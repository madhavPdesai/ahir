-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant R1_base_address : std_logic_vector(0 downto 0) := "0";
  constant R2_base_address : std_logic_vector(0 downto 0) := "0";
  constant R3_base_address : std_logic_vector(0 downto 0) := "0";
  constant frame_base_address : std_logic_vector(0 downto 0) := "0";
  constant key_base_address : std_logic_vector(1 downto 0) := "00";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity a5init is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(1 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    a5reg_call_reqs : out  std_logic_vector(0 downto 0);
    a5reg_call_acks : in   std_logic_vector(0 downto 0);
    a5reg_call_tag  :  out  std_logic_vector(0 downto 0);
    a5reg_return_reqs : out  std_logic_vector(0 downto 0);
    a5reg_return_acks : in   std_logic_vector(0 downto 0);
    a5reg_return_data : in   std_logic_vector(31 downto 0);
    a5reg_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity a5init;
architecture Default of a5init is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal a5init_CP_1104_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_905_gather_scatter_ack_0 : boolean;
  signal binary_957_inst_req_0 : boolean;
  signal binary_992_inst_req_0 : boolean;
  signal binary_986_inst_req_0 : boolean;
  signal simple_obj_ref_899_load_0_ack_1 : boolean;
  signal phi_stmt_912_req_1 : boolean;
  signal binary_986_inst_ack_0 : boolean;
  signal simple_obj_ref_899_load_0_req_1 : boolean;
  signal simple_obj_ref_899_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_899_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_902_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_899_load_0_req_0 : boolean;
  signal simple_obj_ref_895_store_0_req_1 : boolean;
  signal binary_1019_inst_ack_0 : boolean;
  signal binary_1013_inst_req_1 : boolean;
  signal simple_obj_ref_905_gather_scatter_req_0 : boolean;
  signal if_stmt_882_branch_ack_1 : boolean;
  signal simple_obj_ref_892_gather_scatter_req_0 : boolean;
  signal binary_1008_inst_ack_0 : boolean;
  signal simple_obj_ref_899_load_0_ack_0 : boolean;
  signal binary_968_inst_ack_1 : boolean;
  signal simple_obj_ref_902_load_0_ack_0 : boolean;
  signal simple_obj_ref_905_load_0_ack_1 : boolean;
  signal type_cast_934_inst_req_0 : boolean;
  signal if_stmt_882_branch_ack_0 : boolean;
  signal binary_968_inst_req_1 : boolean;
  signal binary_986_inst_req_1 : boolean;
  signal binary_879_inst_req_0 : boolean;
  signal binary_968_inst_ack_0 : boolean;
  signal binary_998_inst_req_1 : boolean;
  signal binary_1008_inst_req_0 : boolean;
  signal binary_968_inst_req_0 : boolean;
  signal binary_1003_inst_ack_0 : boolean;
  signal phi_stmt_651_req_0 : boolean;
  signal binary_952_inst_ack_1 : boolean;
  signal binary_952_inst_req_1 : boolean;
  signal simple_obj_ref_895_store_0_ack_0 : boolean;
  signal simple_obj_ref_895_store_0_req_0 : boolean;
  signal binary_952_inst_ack_0 : boolean;
  signal simple_obj_ref_905_load_0_ack_0 : boolean;
  signal simple_obj_ref_895_store_0_ack_1 : boolean;
  signal binary_1003_inst_ack_1 : boolean;
  signal simple_obj_ref_902_gather_scatter_req_0 : boolean;
  signal binary_952_inst_req_0 : boolean;
  signal binary_879_inst_req_1 : boolean;
  signal simple_obj_ref_905_load_0_req_1 : boolean;
  signal binary_879_inst_ack_0 : boolean;
  signal binary_974_inst_ack_0 : boolean;
  signal binary_998_inst_req_0 : boolean;
  signal binary_749_inst_req_1 : boolean;
  signal binary_727_inst_req_0 : boolean;
  signal binary_727_inst_ack_0 : boolean;
  signal binary_749_inst_ack_1 : boolean;
  signal binary_727_inst_req_1 : boolean;
  signal binary_727_inst_ack_1 : boolean;
  signal binary_703_inst_req_0 : boolean;
  signal binary_879_inst_ack_1 : boolean;
  signal binary_974_inst_ack_1 : boolean;
  signal simple_obj_ref_895_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_902_load_0_ack_1 : boolean;
  signal binary_986_inst_ack_1 : boolean;
  signal simple_obj_ref_895_gather_scatter_ack_0 : boolean;
  signal if_stmt_882_branch_req_0 : boolean;
  signal binary_1013_inst_ack_0 : boolean;
  signal simple_obj_ref_902_load_0_req_0 : boolean;
  signal type_cast_648_inst_ack_0 : boolean;
  signal binary_1003_inst_req_0 : boolean;
  signal simple_obj_ref_905_load_0_req_0 : boolean;
  signal binary_974_inst_req_1 : boolean;
  signal simple_obj_ref_889_store_0_ack_0 : boolean;
  signal binary_962_inst_ack_0 : boolean;
  signal binary_873_inst_ack_1 : boolean;
  signal binary_947_inst_req_0 : boolean;
  signal binary_873_inst_req_1 : boolean;
  signal binary_873_inst_ack_0 : boolean;
  signal simple_obj_ref_889_store_0_req_0 : boolean;
  signal binary_947_inst_ack_1 : boolean;
  signal binary_873_inst_req_0 : boolean;
  signal binary_947_inst_ack_0 : boolean;
  signal binary_980_inst_ack_1 : boolean;
  signal binary_947_inst_req_1 : boolean;
  signal binary_715_inst_ack_1 : boolean;
  signal binary_739_inst_req_0 : boolean;
  signal binary_739_inst_ack_0 : boolean;
  signal binary_739_inst_req_1 : boolean;
  signal simple_obj_ref_908_gather_scatter_ack_0 : boolean;
  signal binary_698_inst_req_0 : boolean;
  signal binary_698_inst_ack_0 : boolean;
  signal binary_754_inst_req_0 : boolean;
  signal simple_obj_ref_902_load_0_req_1 : boolean;
  signal binary_698_inst_req_1 : boolean;
  signal binary_739_inst_ack_1 : boolean;
  signal binary_721_inst_req_0 : boolean;
  signal binary_992_inst_ack_1 : boolean;
  signal binary_721_inst_ack_0 : boolean;
  signal binary_749_inst_req_0 : boolean;
  signal binary_721_inst_req_1 : boolean;
  signal binary_698_inst_ack_1 : boolean;
  signal binary_754_inst_ack_0 : boolean;
  signal binary_721_inst_ack_1 : boolean;
  signal simple_obj_ref_889_gather_scatter_ack_0 : boolean;
  signal binary_749_inst_ack_0 : boolean;
  signal binary_754_inst_req_1 : boolean;
  signal type_cast_654_inst_ack_0 : boolean;
  signal binary_703_inst_ack_0 : boolean;
  signal binary_867_inst_ack_1 : boolean;
  signal simple_obj_ref_892_store_0_ack_1 : boolean;
  signal binary_941_inst_ack_1 : boolean;
  signal binary_703_inst_req_1 : boolean;
  signal binary_703_inst_ack_1 : boolean;
  signal binary_754_inst_ack_1 : boolean;
  signal binary_974_inst_req_0 : boolean;
  signal binary_941_inst_req_1 : boolean;
  signal binary_941_inst_ack_0 : boolean;
  signal binary_733_inst_req_0 : boolean;
  signal binary_867_inst_req_1 : boolean;
  signal binary_733_inst_ack_0 : boolean;
  signal binary_941_inst_req_0 : boolean;
  signal binary_733_inst_req_1 : boolean;
  signal simple_obj_ref_889_gather_scatter_req_0 : boolean;
  signal binary_733_inst_ack_1 : boolean;
  signal binary_744_inst_req_0 : boolean;
  signal binary_709_inst_req_0 : boolean;
  signal binary_709_inst_ack_0 : boolean;
  signal binary_744_inst_ack_0 : boolean;
  signal binary_709_inst_req_1 : boolean;
  signal binary_1003_inst_req_1 : boolean;
  signal binary_709_inst_ack_1 : boolean;
  signal binary_744_inst_req_1 : boolean;
  signal binary_962_inst_req_0 : boolean;
  signal binary_744_inst_ack_1 : boolean;
  signal binary_957_inst_ack_1 : boolean;
  signal binary_715_inst_req_0 : boolean;
  signal binary_715_inst_ack_0 : boolean;
  signal simple_obj_ref_892_store_0_req_1 : boolean;
  signal binary_715_inst_req_1 : boolean;
  signal binary_957_inst_ack_0 : boolean;
  signal binary_957_inst_req_1 : boolean;
  signal binary_992_inst_ack_0 : boolean;
  signal binary_992_inst_req_1 : boolean;
  signal phi_stmt_639_req_0 : boolean;
  signal binary_1042_inst_req_1 : boolean;
  signal type_cast_642_inst_ack_0 : boolean;
  signal binary_1042_inst_ack_1 : boolean;
  signal type_cast_648_inst_req_0 : boolean;
  signal binary_1036_inst_ack_1 : boolean;
  signal binary_980_inst_ack_0 : boolean;
  signal binary_1053_inst_req_0 : boolean;
  signal binary_1053_inst_ack_0 : boolean;
  signal binary_1053_inst_req_1 : boolean;
  signal phi_stmt_919_req_0 : boolean;
  signal type_cast_928_inst_ack_0 : boolean;
  signal type_cast_922_inst_req_0 : boolean;
  signal binary_1042_inst_req_0 : boolean;
  signal binary_1042_inst_ack_0 : boolean;
  signal type_cast_918_inst_ack_0 : boolean;
  signal binary_1019_inst_req_0 : boolean;
  signal binary_980_inst_req_1 : boolean;
  signal binary_1024_inst_req_0 : boolean;
  signal binary_1024_inst_ack_0 : boolean;
  signal binary_998_inst_ack_0 : boolean;
  signal binary_1048_inst_req_1 : boolean;
  signal type_cast_642_inst_req_0 : boolean;
  signal binary_1048_inst_ack_1 : boolean;
  signal binary_1030_inst_req_1 : boolean;
  signal type_cast_928_inst_req_0 : boolean;
  signal binary_1036_inst_ack_0 : boolean;
  signal binary_1036_inst_req_1 : boolean;
  signal binary_980_inst_req_0 : boolean;
  signal binary_998_inst_ack_1 : boolean;
  signal binary_1030_inst_req_0 : boolean;
  signal binary_1030_inst_ack_0 : boolean;
  signal binary_1013_inst_ack_1 : boolean;
  signal binary_1036_inst_req_0 : boolean;
  signal simple_obj_ref_889_store_0_req_1 : boolean;
  signal binary_1024_inst_req_1 : boolean;
  signal binary_1048_inst_req_0 : boolean;
  signal binary_1048_inst_ack_0 : boolean;
  signal simple_obj_ref_889_store_0_ack_1 : boolean;
  signal phi_stmt_925_req_0 : boolean;
  signal type_cast_922_inst_ack_0 : boolean;
  signal binary_1024_inst_ack_1 : boolean;
  signal binary_1030_inst_ack_1 : boolean;
  signal simple_obj_ref_622_load_0_req_0 : boolean;
  signal simple_obj_ref_622_load_0_ack_0 : boolean;
  signal simple_obj_ref_622_load_0_req_1 : boolean;
  signal simple_obj_ref_622_load_0_ack_1 : boolean;
  signal simple_obj_ref_622_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_622_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_625_load_0_req_0 : boolean;
  signal simple_obj_ref_625_load_0_ack_0 : boolean;
  signal simple_obj_ref_625_load_0_req_1 : boolean;
  signal simple_obj_ref_625_load_0_ack_1 : boolean;
  signal simple_obj_ref_625_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_625_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_628_load_0_req_0 : boolean;
  signal simple_obj_ref_628_load_0_ack_0 : boolean;
  signal simple_obj_ref_628_load_0_req_1 : boolean;
  signal simple_obj_ref_628_load_0_ack_1 : boolean;
  signal simple_obj_ref_628_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_628_gather_scatter_ack_0 : boolean;
  signal binary_662_inst_req_0 : boolean;
  signal binary_662_inst_ack_0 : boolean;
  signal binary_662_inst_req_1 : boolean;
  signal binary_662_inst_ack_1 : boolean;
  signal array_obj_ref_666_index_0_resize_req_0 : boolean;
  signal array_obj_ref_666_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_666_index_0_rename_req_0 : boolean;
  signal array_obj_ref_666_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_666_offset_inst_req_0 : boolean;
  signal array_obj_ref_666_offset_inst_ack_0 : boolean;
  signal array_obj_ref_666_root_address_inst_req_0 : boolean;
  signal array_obj_ref_666_root_address_inst_ack_0 : boolean;
  signal addr_of_667_final_reg_req_0 : boolean;
  signal addr_of_667_final_reg_ack_0 : boolean;
  signal ptr_deref_671_base_resize_req_0 : boolean;
  signal ptr_deref_671_base_resize_ack_0 : boolean;
  signal ptr_deref_671_root_address_inst_req_0 : boolean;
  signal ptr_deref_671_root_address_inst_ack_0 : boolean;
  signal ptr_deref_671_addr_0_req_0 : boolean;
  signal ptr_deref_671_addr_0_ack_0 : boolean;
  signal ptr_deref_671_load_0_req_0 : boolean;
  signal ptr_deref_671_load_0_ack_0 : boolean;
  signal ptr_deref_671_load_0_req_1 : boolean;
  signal ptr_deref_671_load_0_ack_1 : boolean;
  signal ptr_deref_671_gather_scatter_req_0 : boolean;
  signal ptr_deref_671_gather_scatter_ack_0 : boolean;
  signal binary_677_inst_req_0 : boolean;
  signal binary_677_inst_ack_0 : boolean;
  signal binary_677_inst_req_1 : boolean;
  signal binary_677_inst_ack_1 : boolean;
  signal binary_682_inst_req_0 : boolean;
  signal binary_682_inst_ack_0 : boolean;
  signal binary_682_inst_req_1 : boolean;
  signal binary_682_inst_ack_1 : boolean;
  signal binary_688_inst_req_0 : boolean;
  signal binary_688_inst_ack_0 : boolean;
  signal binary_688_inst_req_1 : boolean;
  signal binary_688_inst_ack_1 : boolean;
  signal binary_693_inst_req_0 : boolean;
  signal binary_693_inst_ack_0 : boolean;
  signal binary_693_inst_req_1 : boolean;
  signal binary_693_inst_ack_1 : boolean;
  signal binary_867_inst_ack_0 : boolean;
  signal simple_obj_ref_908_gather_scatter_req_0 : boolean;
  signal binary_760_inst_req_0 : boolean;
  signal binary_760_inst_ack_0 : boolean;
  signal simple_obj_ref_908_load_0_ack_1 : boolean;
  signal binary_760_inst_req_1 : boolean;
  signal binary_867_inst_req_0 : boolean;
  signal binary_760_inst_ack_1 : boolean;
  signal binary_1013_inst_req_0 : boolean;
  signal simple_obj_ref_908_load_0_req_1 : boolean;
  signal phi_stmt_645_req_0 : boolean;
  signal binary_765_inst_req_0 : boolean;
  signal binary_765_inst_ack_0 : boolean;
  signal binary_765_inst_req_1 : boolean;
  signal binary_765_inst_ack_1 : boolean;
  signal simple_obj_ref_892_store_0_ack_0 : boolean;
  signal simple_obj_ref_908_load_0_ack_0 : boolean;
  signal simple_obj_ref_908_load_0_req_0 : boolean;
  signal simple_obj_ref_892_store_0_req_0 : boolean;
  signal type_cast_654_inst_req_0 : boolean;
  signal binary_771_inst_req_0 : boolean;
  signal binary_771_inst_ack_0 : boolean;
  signal binary_771_inst_req_1 : boolean;
  signal binary_771_inst_ack_1 : boolean;
  signal binary_1019_inst_ack_1 : boolean;
  signal binary_1008_inst_ack_1 : boolean;
  signal binary_777_inst_req_0 : boolean;
  signal binary_962_inst_ack_1 : boolean;
  signal binary_777_inst_ack_0 : boolean;
  signal binary_777_inst_req_1 : boolean;
  signal binary_777_inst_ack_1 : boolean;
  signal binary_1019_inst_req_1 : boolean;
  signal binary_1008_inst_req_1 : boolean;
  signal simple_obj_ref_892_gather_scatter_ack_0 : boolean;
  signal binary_962_inst_req_1 : boolean;
  signal type_cast_934_inst_ack_0 : boolean;
  signal binary_783_inst_req_0 : boolean;
  signal binary_783_inst_ack_0 : boolean;
  signal binary_783_inst_req_1 : boolean;
  signal binary_783_inst_ack_1 : boolean;
  signal phi_stmt_632_ack_0 : boolean;
  signal binary_789_inst_req_0 : boolean;
  signal binary_789_inst_ack_0 : boolean;
  signal binary_789_inst_req_1 : boolean;
  signal phi_stmt_645_ack_0 : boolean;
  signal binary_789_inst_ack_1 : boolean;
  signal phi_stmt_639_ack_0 : boolean;
  signal binary_794_inst_req_0 : boolean;
  signal binary_794_inst_ack_0 : boolean;
  signal binary_794_inst_req_1 : boolean;
  signal binary_794_inst_ack_1 : boolean;
  signal phi_stmt_931_req_0 : boolean;
  signal phi_stmt_651_ack_0 : boolean;
  signal binary_800_inst_req_0 : boolean;
  signal binary_800_inst_ack_0 : boolean;
  signal binary_800_inst_req_1 : boolean;
  signal binary_800_inst_ack_1 : boolean;
  signal type_cast_918_inst_req_0 : boolean;
  signal phi_stmt_912_ack_0 : boolean;
  signal binary_805_inst_req_0 : boolean;
  signal binary_805_inst_ack_0 : boolean;
  signal binary_805_inst_req_1 : boolean;
  signal binary_805_inst_ack_1 : boolean;
  signal binary_811_inst_req_0 : boolean;
  signal binary_811_inst_ack_0 : boolean;
  signal binary_811_inst_req_1 : boolean;
  signal binary_811_inst_ack_1 : boolean;
  signal phi_stmt_919_ack_0 : boolean;
  signal phi_stmt_925_ack_0 : boolean;
  signal binary_817_inst_req_0 : boolean;
  signal binary_817_inst_ack_0 : boolean;
  signal binary_817_inst_req_1 : boolean;
  signal binary_817_inst_ack_1 : boolean;
  signal phi_stmt_931_ack_0 : boolean;
  signal binary_823_inst_req_0 : boolean;
  signal binary_823_inst_ack_0 : boolean;
  signal binary_823_inst_req_1 : boolean;
  signal binary_823_inst_ack_1 : boolean;
  signal binary_829_inst_req_0 : boolean;
  signal binary_829_inst_ack_0 : boolean;
  signal binary_829_inst_req_1 : boolean;
  signal binary_829_inst_ack_1 : boolean;
  signal binary_835_inst_req_0 : boolean;
  signal binary_835_inst_ack_0 : boolean;
  signal binary_835_inst_req_1 : boolean;
  signal binary_835_inst_ack_1 : boolean;
  signal binary_841_inst_req_0 : boolean;
  signal binary_841_inst_ack_0 : boolean;
  signal binary_841_inst_req_1 : boolean;
  signal binary_841_inst_ack_1 : boolean;
  signal binary_846_inst_req_0 : boolean;
  signal binary_846_inst_ack_0 : boolean;
  signal binary_846_inst_req_1 : boolean;
  signal binary_846_inst_ack_1 : boolean;
  signal binary_851_inst_req_0 : boolean;
  signal binary_851_inst_ack_0 : boolean;
  signal binary_851_inst_req_1 : boolean;
  signal binary_851_inst_ack_1 : boolean;
  signal binary_856_inst_req_0 : boolean;
  signal binary_856_inst_ack_0 : boolean;
  signal binary_856_inst_req_1 : boolean;
  signal binary_856_inst_ack_1 : boolean;
  signal binary_862_inst_req_0 : boolean;
  signal binary_862_inst_ack_0 : boolean;
  signal binary_862_inst_req_1 : boolean;
  signal binary_862_inst_ack_1 : boolean;
  signal binary_1053_inst_ack_1 : boolean;
  signal binary_1059_inst_req_0 : boolean;
  signal binary_1059_inst_ack_0 : boolean;
  signal binary_1059_inst_req_1 : boolean;
  signal binary_1059_inst_ack_1 : boolean;
  signal phi_stmt_912_req_0 : boolean;
  signal binary_1064_inst_req_0 : boolean;
  signal binary_1064_inst_ack_0 : boolean;
  signal binary_1064_inst_req_1 : boolean;
  signal binary_1064_inst_ack_1 : boolean;
  signal binary_1070_inst_req_0 : boolean;
  signal binary_1070_inst_ack_0 : boolean;
  signal binary_1070_inst_req_1 : boolean;
  signal binary_1070_inst_ack_1 : boolean;
  signal binary_1076_inst_req_0 : boolean;
  signal binary_1076_inst_ack_0 : boolean;
  signal binary_1076_inst_req_1 : boolean;
  signal binary_1076_inst_ack_1 : boolean;
  signal phi_stmt_931_req_1 : boolean;
  signal binary_1082_inst_req_0 : boolean;
  signal binary_1082_inst_ack_0 : boolean;
  signal binary_1082_inst_req_1 : boolean;
  signal phi_stmt_632_req_0 : boolean;
  signal binary_1082_inst_ack_1 : boolean;
  signal type_cast_936_inst_ack_0 : boolean;
  signal type_cast_936_inst_req_0 : boolean;
  signal binary_1088_inst_req_0 : boolean;
  signal binary_1088_inst_ack_0 : boolean;
  signal binary_1088_inst_req_1 : boolean;
  signal binary_1088_inst_ack_1 : boolean;
  signal binary_1094_inst_req_0 : boolean;
  signal binary_1094_inst_ack_0 : boolean;
  signal binary_1094_inst_req_1 : boolean;
  signal binary_1094_inst_ack_1 : boolean;
  signal binary_1100_inst_req_0 : boolean;
  signal binary_1100_inst_ack_0 : boolean;
  signal binary_1100_inst_req_1 : boolean;
  signal binary_1100_inst_ack_1 : boolean;
  signal phi_stmt_925_req_1 : boolean;
  signal binary_1105_inst_req_0 : boolean;
  signal binary_1105_inst_ack_0 : boolean;
  signal binary_1105_inst_req_1 : boolean;
  signal binary_1105_inst_ack_1 : boolean;
  signal type_cast_930_inst_ack_0 : boolean;
  signal type_cast_930_inst_req_0 : boolean;
  signal binary_1110_inst_req_0 : boolean;
  signal binary_1110_inst_ack_0 : boolean;
  signal binary_1110_inst_req_1 : boolean;
  signal binary_1110_inst_ack_1 : boolean;
  signal binary_1115_inst_req_0 : boolean;
  signal binary_1115_inst_ack_0 : boolean;
  signal binary_1115_inst_req_1 : boolean;
  signal binary_1115_inst_ack_1 : boolean;
  signal phi_stmt_1158_ack_0 : boolean;
  signal binary_1121_inst_req_0 : boolean;
  signal binary_1121_inst_ack_0 : boolean;
  signal phi_stmt_1158_req_0 : boolean;
  signal binary_1121_inst_req_1 : boolean;
  signal binary_1121_inst_ack_1 : boolean;
  signal phi_stmt_919_req_1 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal binary_1126_inst_req_0 : boolean;
  signal binary_1126_inst_ack_0 : boolean;
  signal binary_1126_inst_req_1 : boolean;
  signal binary_1126_inst_ack_1 : boolean;
  signal binary_1132_inst_req_0 : boolean;
  signal binary_1132_inst_ack_0 : boolean;
  signal phi_stmt_1158_req_1 : boolean;
  signal binary_1132_inst_req_1 : boolean;
  signal binary_1132_inst_ack_1 : boolean;
  signal type_cast_1165_inst_ack_0 : boolean;
  signal type_cast_1165_inst_req_0 : boolean;
  signal binary_1138_inst_req_0 : boolean;
  signal binary_1138_inst_ack_0 : boolean;
  signal binary_1138_inst_req_1 : boolean;
  signal binary_1138_inst_ack_1 : boolean;
  signal if_stmt_1140_branch_req_0 : boolean;
  signal if_stmt_1140_branch_ack_1 : boolean;
  signal if_stmt_1140_branch_ack_0 : boolean;
  signal simple_obj_ref_1147_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1147_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1147_store_0_req_0 : boolean;
  signal simple_obj_ref_1147_store_0_ack_0 : boolean;
  signal simple_obj_ref_1147_store_0_req_1 : boolean;
  signal simple_obj_ref_1147_store_0_ack_1 : boolean;
  signal simple_obj_ref_1150_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1150_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1150_store_0_req_0 : boolean;
  signal simple_obj_ref_1150_store_0_ack_0 : boolean;
  signal simple_obj_ref_1150_store_0_req_1 : boolean;
  signal simple_obj_ref_1150_store_0_ack_1 : boolean;
  signal simple_obj_ref_1153_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1153_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1153_store_0_req_0 : boolean;
  signal simple_obj_ref_1153_store_0_ack_0 : boolean;
  signal simple_obj_ref_1153_store_0_req_1 : boolean;
  signal simple_obj_ref_1153_store_0_ack_1 : boolean;
  signal call_stmt_1168_call_req_0 : boolean;
  signal call_stmt_1168_call_ack_0 : boolean;
  signal call_stmt_1168_call_req_1 : boolean;
  signal call_stmt_1168_call_ack_1 : boolean;
  signal binary_1173_inst_req_0 : boolean;
  signal binary_1173_inst_ack_0 : boolean;
  signal binary_1173_inst_req_1 : boolean;
  signal binary_1173_inst_ack_1 : boolean;
  signal binary_1179_inst_req_0 : boolean;
  signal binary_1179_inst_ack_0 : boolean;
  signal binary_1179_inst_req_1 : boolean;
  signal binary_1179_inst_ack_1 : boolean;
  signal if_stmt_1181_branch_req_0 : boolean;
  signal if_stmt_1181_branch_ack_1 : boolean;
  signal if_stmt_1181_branch_ack_0 : boolean;
  signal type_cast_638_inst_req_0 : boolean;
  signal type_cast_638_inst_ack_0 : boolean;
  signal phi_stmt_632_req_1 : boolean;
  signal type_cast_644_inst_req_0 : boolean;
  signal type_cast_644_inst_ack_0 : boolean;
  signal phi_stmt_639_req_1 : boolean;
  signal type_cast_650_inst_req_0 : boolean;
  signal type_cast_650_inst_ack_0 : boolean;
  signal phi_stmt_645_req_1 : boolean;
  signal type_cast_656_inst_req_0 : boolean;
  signal type_cast_656_inst_ack_0 : boolean;
  signal phi_stmt_651_req_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  a5init_CP_1104: Block -- control-path 
    signal cp_elements: BooleanArray(582 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(10);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(10), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(24);
    cp_elements(2) <= cp_elements(528);
    cp_elements(3) <= cp_elements(215);
    cp_elements(4) <= OrReduce(cp_elements(222) & cp_elements(530));
    cp_elements(5) <= cp_elements(266);
    cp_elements(6) <= cp_elements(574);
    cp_elements(7) <= cp_elements(434);
    cp_elements(8) <= OrReduce(cp_elements(441) & cp_elements(576));
    cp_elements(9) <= cp_elements(463);
    phi_stmt_1158_req_0 <= cp_elements(9);
    cp_elements(10) <= OrReduce(cp_elements(482) & cp_elements(582));
    cp_elements(11) <= cp_elements(0);
    cp_elements(12) <= cp_elements(11);
    simple_obj_ref_622_load_0_req_0 <= cp_elements(12);
    cp_elements(13) <= simple_obj_ref_622_load_0_ack_0;
    simple_obj_ref_622_load_0_req_1 <= cp_elements(13);
    cp_elements(14) <= simple_obj_ref_622_load_0_ack_1;
    simple_obj_ref_622_gather_scatter_req_0 <= cp_elements(14);
    cp_elements(15) <= simple_obj_ref_622_gather_scatter_ack_0;
    cp_elements(16) <= cp_elements(11);
    simple_obj_ref_625_load_0_req_0 <= cp_elements(16);
    cp_elements(17) <= simple_obj_ref_625_load_0_ack_0;
    simple_obj_ref_625_load_0_req_1 <= cp_elements(17);
    cp_elements(18) <= simple_obj_ref_625_load_0_ack_1;
    simple_obj_ref_625_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= simple_obj_ref_625_gather_scatter_ack_0;
    cp_elements(20) <= cp_elements(11);
    simple_obj_ref_628_load_0_req_0 <= cp_elements(20);
    cp_elements(21) <= simple_obj_ref_628_load_0_ack_0;
    simple_obj_ref_628_load_0_req_1 <= cp_elements(21);
    cp_elements(22) <= simple_obj_ref_628_load_0_ack_1;
    simple_obj_ref_628_gather_scatter_req_0 <= cp_elements(22);
    cp_elements(23) <= simple_obj_ref_628_gather_scatter_ack_0;
    cpelement_group_24 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(23) & cp_elements(15));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(24),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(25) <= cp_elements(2);
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(28));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_662_inst_req_0 <= cp_elements(26);
    cp_elements(27) <= cp_elements(25);
    cp_elements(28) <= cp_elements(25);
    cp_elements(29) <= binary_662_inst_ack_0;
    binary_662_inst_req_1 <= cp_elements(29);
    cp_elements(30) <= binary_662_inst_ack_1;
    array_obj_ref_666_index_0_resize_req_0 <= cp_elements(30);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(36));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_667_final_reg_req_0 <= cp_elements(31);
    cp_elements(32) <= cp_elements(25);
    cp_elements(33) <= array_obj_ref_666_index_0_resize_ack_0;
    array_obj_ref_666_index_0_rename_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_666_index_0_rename_ack_0;
    array_obj_ref_666_offset_inst_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_666_offset_inst_ack_0;
    array_obj_ref_666_root_address_inst_req_0 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_666_root_address_inst_ack_0;
    cp_elements(37) <= addr_of_667_final_reg_ack_0;
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(37));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_671_load_0_req_0 <= cp_elements(38);
    cp_elements(39) <= cp_elements(37);
    ptr_deref_671_base_resize_req_0 <= cp_elements(39);
    cp_elements(40) <= ptr_deref_671_base_resize_ack_0;
    ptr_deref_671_root_address_inst_req_0 <= cp_elements(40);
    cp_elements(41) <= ptr_deref_671_root_address_inst_ack_0;
    ptr_deref_671_addr_0_req_0 <= cp_elements(41);
    cp_elements(42) <= ptr_deref_671_addr_0_ack_0;
    cp_elements(43) <= ptr_deref_671_load_0_ack_0;
    ptr_deref_671_load_0_req_1 <= cp_elements(43);
    cp_elements(44) <= ptr_deref_671_load_0_ack_1;
    ptr_deref_671_gather_scatter_req_0 <= cp_elements(44);
    cp_elements(45) <= ptr_deref_671_gather_scatter_ack_0;
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(47) & cp_elements(48));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_677_inst_req_0 <= cp_elements(46);
    cp_elements(47) <= cp_elements(25);
    cp_elements(48) <= cp_elements(25);
    cp_elements(49) <= binary_677_inst_ack_0;
    binary_677_inst_req_1 <= cp_elements(49);
    cp_elements(50) <= binary_677_inst_ack_1;
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(50) & cp_elements(52));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_682_inst_req_0 <= cp_elements(51);
    cp_elements(52) <= cp_elements(25);
    cp_elements(53) <= binary_682_inst_ack_0;
    binary_682_inst_req_1 <= cp_elements(53);
    cp_elements(54) <= binary_682_inst_ack_1;
    cpelement_group_55 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(54) & cp_elements(56));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(55),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_688_inst_req_0 <= cp_elements(55);
    cp_elements(56) <= cp_elements(25);
    cp_elements(57) <= binary_688_inst_ack_0;
    binary_688_inst_req_1 <= cp_elements(57);
    cp_elements(58) <= binary_688_inst_ack_1;
    cpelement_group_59 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(59),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_693_inst_req_0 <= cp_elements(59);
    cp_elements(60) <= cp_elements(25);
    cp_elements(61) <= cp_elements(58);
    cp_elements(62) <= cp_elements(25);
    cp_elements(63) <= binary_693_inst_ack_0;
    binary_693_inst_req_1 <= cp_elements(63);
    cp_elements(64) <= binary_693_inst_ack_1;
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(67) & cp_elements(68));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_698_inst_req_0 <= cp_elements(65);
    cp_elements(66) <= cp_elements(25);
    cp_elements(67) <= cp_elements(25);
    cp_elements(68) <= cp_elements(58);
    cp_elements(69) <= binary_698_inst_ack_0;
    binary_698_inst_req_1 <= cp_elements(69);
    cp_elements(70) <= binary_698_inst_ack_1;
    cpelement_group_71 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(72) & cp_elements(73) & cp_elements(74));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(71),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_703_inst_req_0 <= cp_elements(71);
    cp_elements(72) <= cp_elements(25);
    cp_elements(73) <= cp_elements(25);
    cp_elements(74) <= cp_elements(58);
    cp_elements(75) <= binary_703_inst_ack_0;
    binary_703_inst_req_1 <= cp_elements(75);
    cp_elements(76) <= binary_703_inst_ack_1;
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(79));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_709_inst_req_0 <= cp_elements(77);
    cp_elements(78) <= cp_elements(25);
    cp_elements(79) <= cp_elements(64);
    cp_elements(80) <= binary_709_inst_ack_0;
    binary_709_inst_req_1 <= cp_elements(80);
    cp_elements(81) <= binary_709_inst_ack_1;
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(84));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_715_inst_req_0 <= cp_elements(82);
    cp_elements(83) <= cp_elements(25);
    cp_elements(84) <= cp_elements(64);
    cp_elements(85) <= binary_715_inst_ack_0;
    binary_715_inst_req_1 <= cp_elements(85);
    cp_elements(86) <= binary_715_inst_ack_1;
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(88) & cp_elements(89));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_721_inst_req_0 <= cp_elements(87);
    cp_elements(88) <= cp_elements(25);
    cp_elements(89) <= cp_elements(64);
    cp_elements(90) <= binary_721_inst_ack_0;
    binary_721_inst_req_1 <= cp_elements(90);
    cp_elements(91) <= binary_721_inst_ack_1;
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(94));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_727_inst_req_0 <= cp_elements(92);
    cp_elements(93) <= cp_elements(25);
    cp_elements(94) <= cp_elements(64);
    cp_elements(95) <= binary_727_inst_ack_0;
    binary_727_inst_req_1 <= cp_elements(95);
    cp_elements(96) <= binary_727_inst_ack_1;
    cpelement_group_97 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(98) & cp_elements(99));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(97),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_733_inst_req_0 <= cp_elements(97);
    cp_elements(98) <= cp_elements(25);
    cp_elements(99) <= cp_elements(64);
    cp_elements(100) <= binary_733_inst_ack_0;
    binary_733_inst_req_1 <= cp_elements(100);
    cp_elements(101) <= binary_733_inst_ack_1;
    cpelement_group_102 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(101) & cp_elements(103));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(102),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_739_inst_req_0 <= cp_elements(102);
    cp_elements(103) <= cp_elements(25);
    cp_elements(104) <= binary_739_inst_ack_0;
    binary_739_inst_req_1 <= cp_elements(104);
    cp_elements(105) <= binary_739_inst_ack_1;
    cpelement_group_106 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(86) & cp_elements(107));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(106),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_744_inst_req_0 <= cp_elements(106);
    cp_elements(107) <= cp_elements(25);
    cp_elements(108) <= binary_744_inst_ack_0;
    binary_744_inst_req_1 <= cp_elements(108);
    cp_elements(109) <= binary_744_inst_ack_1;
    cpelement_group_110 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(96) & cp_elements(109) & cp_elements(111));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(110),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_749_inst_req_0 <= cp_elements(110);
    cp_elements(111) <= cp_elements(25);
    cp_elements(112) <= binary_749_inst_ack_0;
    binary_749_inst_req_1 <= cp_elements(112);
    cp_elements(113) <= binary_749_inst_ack_1;
    cpelement_group_114 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(113) & cp_elements(115));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(114),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_754_inst_req_0 <= cp_elements(114);
    cp_elements(115) <= cp_elements(25);
    cp_elements(116) <= binary_754_inst_ack_0;
    binary_754_inst_req_1 <= cp_elements(116);
    cp_elements(117) <= binary_754_inst_ack_1;
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(117) & cp_elements(119));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_760_inst_req_0 <= cp_elements(118);
    cp_elements(119) <= cp_elements(25);
    cp_elements(120) <= binary_760_inst_ack_0;
    binary_760_inst_req_1 <= cp_elements(120);
    cp_elements(121) <= binary_760_inst_ack_1;
    cpelement_group_122 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(105) & cp_elements(121) & cp_elements(123));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(122),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_765_inst_req_0 <= cp_elements(122);
    cp_elements(123) <= cp_elements(25);
    cp_elements(124) <= binary_765_inst_ack_0;
    binary_765_inst_req_1 <= cp_elements(124);
    cp_elements(125) <= binary_765_inst_ack_1;
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(128));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_771_inst_req_0 <= cp_elements(126);
    cp_elements(127) <= cp_elements(25);
    cp_elements(128) <= cp_elements(70);
    cp_elements(129) <= binary_771_inst_ack_0;
    binary_771_inst_req_1 <= cp_elements(129);
    cp_elements(130) <= binary_771_inst_ack_1;
    cpelement_group_131 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(132) & cp_elements(133));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(131),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_777_inst_req_0 <= cp_elements(131);
    cp_elements(132) <= cp_elements(25);
    cp_elements(133) <= cp_elements(70);
    cp_elements(134) <= binary_777_inst_ack_0;
    binary_777_inst_req_1 <= cp_elements(134);
    cp_elements(135) <= binary_777_inst_ack_1;
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(138));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_783_inst_req_0 <= cp_elements(136);
    cp_elements(137) <= cp_elements(25);
    cp_elements(138) <= cp_elements(70);
    cp_elements(139) <= binary_783_inst_ack_0;
    binary_783_inst_req_1 <= cp_elements(139);
    cp_elements(140) <= binary_783_inst_ack_1;
    cpelement_group_141 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(140) & cp_elements(142));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(141),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_789_inst_req_0 <= cp_elements(141);
    cp_elements(142) <= cp_elements(25);
    cp_elements(143) <= binary_789_inst_ack_0;
    binary_789_inst_req_1 <= cp_elements(143);
    cp_elements(144) <= binary_789_inst_ack_1;
    cpelement_group_145 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(130) & cp_elements(135) & cp_elements(146));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(145),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_794_inst_req_0 <= cp_elements(145);
    cp_elements(146) <= cp_elements(25);
    cp_elements(147) <= binary_794_inst_ack_0;
    binary_794_inst_req_1 <= cp_elements(147);
    cp_elements(148) <= binary_794_inst_ack_1;
    cpelement_group_149 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(149),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_800_inst_req_0 <= cp_elements(149);
    cp_elements(150) <= cp_elements(25);
    cp_elements(151) <= binary_800_inst_ack_0;
    binary_800_inst_req_1 <= cp_elements(151);
    cp_elements(152) <= binary_800_inst_ack_1;
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(144) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_805_inst_req_0 <= cp_elements(153);
    cp_elements(154) <= cp_elements(25);
    cp_elements(155) <= binary_805_inst_ack_0;
    binary_805_inst_req_1 <= cp_elements(155);
    cp_elements(156) <= binary_805_inst_ack_1;
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(158) & cp_elements(159));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_811_inst_req_0 <= cp_elements(157);
    cp_elements(158) <= cp_elements(25);
    cp_elements(159) <= cp_elements(76);
    cp_elements(160) <= binary_811_inst_ack_0;
    binary_811_inst_req_1 <= cp_elements(160);
    cp_elements(161) <= binary_811_inst_ack_1;
    cpelement_group_162 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(163) & cp_elements(164));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(162),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_817_inst_req_0 <= cp_elements(162);
    cp_elements(163) <= cp_elements(25);
    cp_elements(164) <= cp_elements(76);
    cp_elements(165) <= binary_817_inst_ack_0;
    binary_817_inst_req_1 <= cp_elements(165);
    cp_elements(166) <= binary_817_inst_ack_1;
    cpelement_group_167 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(168) & cp_elements(169));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(167),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_823_inst_req_0 <= cp_elements(167);
    cp_elements(168) <= cp_elements(25);
    cp_elements(169) <= cp_elements(76);
    cp_elements(170) <= binary_823_inst_ack_0;
    binary_823_inst_req_1 <= cp_elements(170);
    cp_elements(171) <= binary_823_inst_ack_1;
    cpelement_group_172 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(173) & cp_elements(174));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(172),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_829_inst_req_0 <= cp_elements(172);
    cp_elements(173) <= cp_elements(25);
    cp_elements(174) <= cp_elements(76);
    cp_elements(175) <= binary_829_inst_ack_0;
    binary_829_inst_req_1 <= cp_elements(175);
    cp_elements(176) <= binary_829_inst_ack_1;
    cpelement_group_177 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(179));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(177),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_835_inst_req_0 <= cp_elements(177);
    cp_elements(178) <= cp_elements(25);
    cp_elements(179) <= cp_elements(76);
    cp_elements(180) <= binary_835_inst_ack_0;
    binary_835_inst_req_1 <= cp_elements(180);
    cp_elements(181) <= binary_835_inst_ack_1;
    cpelement_group_182 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(183));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(182),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_841_inst_req_0 <= cp_elements(182);
    cp_elements(183) <= cp_elements(25);
    cp_elements(184) <= binary_841_inst_ack_0;
    binary_841_inst_req_1 <= cp_elements(184);
    cp_elements(185) <= binary_841_inst_ack_1;
    cpelement_group_186 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(161) & cp_elements(166) & cp_elements(187));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(186),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_846_inst_req_0 <= cp_elements(186);
    cp_elements(187) <= cp_elements(25);
    cp_elements(188) <= binary_846_inst_ack_0;
    binary_846_inst_req_1 <= cp_elements(188);
    cp_elements(189) <= binary_846_inst_ack_1;
    cpelement_group_190 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(176) & cp_elements(189) & cp_elements(191));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(190),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_851_inst_req_0 <= cp_elements(190);
    cp_elements(191) <= cp_elements(25);
    cp_elements(192) <= binary_851_inst_ack_0;
    binary_851_inst_req_1 <= cp_elements(192);
    cp_elements(193) <= binary_851_inst_ack_1;
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(171) & cp_elements(193) & cp_elements(195));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_856_inst_req_0 <= cp_elements(194);
    cp_elements(195) <= cp_elements(25);
    cp_elements(196) <= binary_856_inst_ack_0;
    binary_856_inst_req_1 <= cp_elements(196);
    cp_elements(197) <= binary_856_inst_ack_1;
    cpelement_group_198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(197) & cp_elements(199));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_862_inst_req_0 <= cp_elements(198);
    cp_elements(199) <= cp_elements(25);
    cp_elements(200) <= binary_862_inst_ack_0;
    binary_862_inst_req_1 <= cp_elements(200);
    cp_elements(201) <= binary_862_inst_ack_1;
    cpelement_group_202 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(185) & cp_elements(201) & cp_elements(203));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(202),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_867_inst_req_0 <= cp_elements(202);
    cp_elements(203) <= cp_elements(25);
    cp_elements(204) <= binary_867_inst_ack_0;
    binary_867_inst_req_1 <= cp_elements(204);
    cp_elements(205) <= binary_867_inst_ack_1;
    cpelement_group_206 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(207) & cp_elements(208));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(206),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_873_inst_req_0 <= cp_elements(206);
    cp_elements(207) <= cp_elements(25);
    cp_elements(208) <= cp_elements(25);
    cp_elements(209) <= binary_873_inst_ack_0;
    binary_873_inst_req_1 <= cp_elements(209);
    cp_elements(210) <= binary_873_inst_ack_1;
    cpelement_group_211 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(210) & cp_elements(212));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_879_inst_req_0 <= cp_elements(211);
    cp_elements(212) <= cp_elements(25);
    cp_elements(213) <= binary_879_inst_ack_0;
    binary_879_inst_req_1 <= cp_elements(213);
    cp_elements(214) <= binary_879_inst_ack_1;
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(205) & cp_elements(214) & cp_elements(125));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= cp_elements(3);
    cp_elements(217) <= false;
    cp_elements(218) <= cp_elements(217);
    cp_elements(219) <= cp_elements(3);
    if_stmt_882_branch_req_0 <= cp_elements(219);
    cp_elements(220) <= cp_elements(219);
    cp_elements(221) <= cp_elements(220);
    cp_elements(222) <= if_stmt_882_branch_ack_1;
    cp_elements(223) <= cp_elements(220);
    cp_elements(224) <= if_stmt_882_branch_ack_0;
    cp_elements(225) <= cp_elements(4);
    cp_elements(226) <= cp_elements(225);
    cpelement_group_227 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(226) & cp_elements(228));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(227),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_889_gather_scatter_req_0 <= cp_elements(227);
    cp_elements(228) <= cp_elements(225);
    cp_elements(229) <= simple_obj_ref_889_gather_scatter_ack_0;
    simple_obj_ref_889_store_0_req_0 <= cp_elements(229);
    cp_elements(230) <= simple_obj_ref_889_store_0_ack_0;
    cp_elements(231) <= cp_elements(230);
    simple_obj_ref_889_store_0_req_1 <= cp_elements(231);
    cp_elements(232) <= simple_obj_ref_889_store_0_ack_1;
    cp_elements(233) <= cp_elements(225);
    cpelement_group_234 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(233) & cp_elements(235));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(234),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_892_gather_scatter_req_0 <= cp_elements(234);
    cp_elements(235) <= cp_elements(225);
    cp_elements(236) <= simple_obj_ref_892_gather_scatter_ack_0;
    simple_obj_ref_892_store_0_req_0 <= cp_elements(236);
    cp_elements(237) <= simple_obj_ref_892_store_0_ack_0;
    cp_elements(238) <= cp_elements(237);
    simple_obj_ref_892_store_0_req_1 <= cp_elements(238);
    cp_elements(239) <= simple_obj_ref_892_store_0_ack_1;
    cp_elements(240) <= cp_elements(225);
    cpelement_group_241 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(240) & cp_elements(242));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(241),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_895_gather_scatter_req_0 <= cp_elements(241);
    cp_elements(242) <= cp_elements(225);
    cp_elements(243) <= simple_obj_ref_895_gather_scatter_ack_0;
    simple_obj_ref_895_store_0_req_0 <= cp_elements(243);
    cp_elements(244) <= simple_obj_ref_895_store_0_ack_0;
    cp_elements(245) <= cp_elements(244);
    simple_obj_ref_895_store_0_req_1 <= cp_elements(245);
    cp_elements(246) <= simple_obj_ref_895_store_0_ack_1;
    cp_elements(247) <= cp_elements(225);
    simple_obj_ref_899_load_0_req_0 <= cp_elements(247);
    cp_elements(248) <= simple_obj_ref_899_load_0_ack_0;
    simple_obj_ref_899_load_0_req_1 <= cp_elements(248);
    cp_elements(249) <= simple_obj_ref_899_load_0_ack_1;
    simple_obj_ref_899_gather_scatter_req_0 <= cp_elements(249);
    cp_elements(250) <= simple_obj_ref_899_gather_scatter_ack_0;
    cpelement_group_251 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(244) & cp_elements(252));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(251),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_902_load_0_req_0 <= cp_elements(251);
    cp_elements(252) <= cp_elements(225);
    cp_elements(253) <= simple_obj_ref_902_load_0_ack_0;
    simple_obj_ref_902_load_0_req_1 <= cp_elements(253);
    cp_elements(254) <= simple_obj_ref_902_load_0_ack_1;
    simple_obj_ref_902_gather_scatter_req_0 <= cp_elements(254);
    cp_elements(255) <= simple_obj_ref_902_gather_scatter_ack_0;
    cpelement_group_256 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(237) & cp_elements(257));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(256),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_905_load_0_req_0 <= cp_elements(256);
    cp_elements(257) <= cp_elements(225);
    cp_elements(258) <= simple_obj_ref_905_load_0_ack_0;
    simple_obj_ref_905_load_0_req_1 <= cp_elements(258);
    cp_elements(259) <= simple_obj_ref_905_load_0_ack_1;
    simple_obj_ref_905_gather_scatter_req_0 <= cp_elements(259);
    cp_elements(260) <= simple_obj_ref_905_gather_scatter_ack_0;
    cpelement_group_261 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(262));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(261),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_908_load_0_req_0 <= cp_elements(261);
    cp_elements(262) <= cp_elements(225);
    cp_elements(263) <= simple_obj_ref_908_load_0_ack_0;
    simple_obj_ref_908_load_0_req_1 <= cp_elements(263);
    cp_elements(264) <= simple_obj_ref_908_load_0_ack_1;
    simple_obj_ref_908_gather_scatter_req_0 <= cp_elements(264);
    cp_elements(265) <= simple_obj_ref_908_gather_scatter_ack_0;
    cpelement_group_266 : Block -- 
      signal predecessors: BooleanArray(6 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(232) & cp_elements(239) & cp_elements(246) & cp_elements(250) & cp_elements(255) & cp_elements(260) & cp_elements(265));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(266),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(267) <= cp_elements(6);
    cpelement_group_268 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(269) & cp_elements(270) & cp_elements(271));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(268),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_941_inst_req_0 <= cp_elements(268);
    cp_elements(269) <= cp_elements(267);
    cp_elements(270) <= cp_elements(267);
    cp_elements(271) <= cp_elements(267);
    cp_elements(272) <= binary_941_inst_ack_0;
    binary_941_inst_req_1 <= cp_elements(272);
    cp_elements(273) <= binary_941_inst_ack_1;
    cpelement_group_274 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(273) & cp_elements(275));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(274),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_947_inst_req_0 <= cp_elements(274);
    cp_elements(275) <= cp_elements(267);
    cp_elements(276) <= binary_947_inst_ack_0;
    binary_947_inst_req_1 <= cp_elements(276);
    cp_elements(277) <= binary_947_inst_ack_1;
    cpelement_group_278 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(279) & cp_elements(280) & cp_elements(281));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(278),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_952_inst_req_0 <= cp_elements(278);
    cp_elements(279) <= cp_elements(267);
    cp_elements(280) <= cp_elements(277);
    cp_elements(281) <= cp_elements(267);
    cp_elements(282) <= binary_952_inst_ack_0;
    binary_952_inst_req_1 <= cp_elements(282);
    cp_elements(283) <= binary_952_inst_ack_1;
    cpelement_group_284 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(285) & cp_elements(286) & cp_elements(287));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(284),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_957_inst_req_0 <= cp_elements(284);
    cp_elements(285) <= cp_elements(267);
    cp_elements(286) <= cp_elements(267);
    cp_elements(287) <= cp_elements(277);
    cp_elements(288) <= binary_957_inst_ack_0;
    binary_957_inst_req_1 <= cp_elements(288);
    cp_elements(289) <= binary_957_inst_ack_1;
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(292) & cp_elements(293));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_962_inst_req_0 <= cp_elements(290);
    cp_elements(291) <= cp_elements(267);
    cp_elements(292) <= cp_elements(267);
    cp_elements(293) <= cp_elements(277);
    cp_elements(294) <= binary_962_inst_ack_0;
    binary_962_inst_req_1 <= cp_elements(294);
    cp_elements(295) <= binary_962_inst_ack_1;
    cpelement_group_296 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(297) & cp_elements(298));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(296),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_968_inst_req_0 <= cp_elements(296);
    cp_elements(297) <= cp_elements(267);
    cp_elements(298) <= cp_elements(283);
    cp_elements(299) <= binary_968_inst_ack_0;
    binary_968_inst_req_1 <= cp_elements(299);
    cp_elements(300) <= binary_968_inst_ack_1;
    cpelement_group_301 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(302) & cp_elements(303));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(301),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_974_inst_req_0 <= cp_elements(301);
    cp_elements(302) <= cp_elements(267);
    cp_elements(303) <= cp_elements(283);
    cp_elements(304) <= binary_974_inst_ack_0;
    binary_974_inst_req_1 <= cp_elements(304);
    cp_elements(305) <= binary_974_inst_ack_1;
    cpelement_group_306 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(307) & cp_elements(308));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(306),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_980_inst_req_0 <= cp_elements(306);
    cp_elements(307) <= cp_elements(267);
    cp_elements(308) <= cp_elements(283);
    cp_elements(309) <= binary_980_inst_ack_0;
    binary_980_inst_req_1 <= cp_elements(309);
    cp_elements(310) <= binary_980_inst_ack_1;
    cpelement_group_311 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(312) & cp_elements(313));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(311),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_986_inst_req_0 <= cp_elements(311);
    cp_elements(312) <= cp_elements(267);
    cp_elements(313) <= cp_elements(283);
    cp_elements(314) <= binary_986_inst_ack_0;
    binary_986_inst_req_1 <= cp_elements(314);
    cp_elements(315) <= binary_986_inst_ack_1;
    cpelement_group_316 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(317) & cp_elements(318));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(316),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_992_inst_req_0 <= cp_elements(316);
    cp_elements(317) <= cp_elements(267);
    cp_elements(318) <= cp_elements(283);
    cp_elements(319) <= binary_992_inst_ack_0;
    binary_992_inst_req_1 <= cp_elements(319);
    cp_elements(320) <= binary_992_inst_ack_1;
    cpelement_group_321 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(320) & cp_elements(322));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(321),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_998_inst_req_0 <= cp_elements(321);
    cp_elements(322) <= cp_elements(267);
    cp_elements(323) <= binary_998_inst_ack_0;
    binary_998_inst_req_1 <= cp_elements(323);
    cp_elements(324) <= binary_998_inst_ack_1;
    cpelement_group_325 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(300) & cp_elements(305) & cp_elements(326));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(325),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1003_inst_req_0 <= cp_elements(325);
    cp_elements(326) <= cp_elements(267);
    cp_elements(327) <= binary_1003_inst_ack_0;
    binary_1003_inst_req_1 <= cp_elements(327);
    cp_elements(328) <= binary_1003_inst_ack_1;
    cpelement_group_329 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(315) & cp_elements(328) & cp_elements(330));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(329),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1008_inst_req_0 <= cp_elements(329);
    cp_elements(330) <= cp_elements(267);
    cp_elements(331) <= binary_1008_inst_ack_0;
    binary_1008_inst_req_1 <= cp_elements(331);
    cp_elements(332) <= binary_1008_inst_ack_1;
    cpelement_group_333 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(310) & cp_elements(332) & cp_elements(334));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(333),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1013_inst_req_0 <= cp_elements(333);
    cp_elements(334) <= cp_elements(267);
    cp_elements(335) <= binary_1013_inst_ack_0;
    binary_1013_inst_req_1 <= cp_elements(335);
    cp_elements(336) <= binary_1013_inst_ack_1;
    cpelement_group_337 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(336) & cp_elements(338));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(337),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1019_inst_req_0 <= cp_elements(337);
    cp_elements(338) <= cp_elements(267);
    cp_elements(339) <= binary_1019_inst_ack_0;
    binary_1019_inst_req_1 <= cp_elements(339);
    cp_elements(340) <= binary_1019_inst_ack_1;
    cpelement_group_341 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(324) & cp_elements(340) & cp_elements(342));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(341),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1024_inst_req_0 <= cp_elements(341);
    cp_elements(342) <= cp_elements(267);
    cp_elements(343) <= binary_1024_inst_ack_0;
    binary_1024_inst_req_1 <= cp_elements(343);
    cp_elements(344) <= binary_1024_inst_ack_1;
    cpelement_group_345 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(346) & cp_elements(347));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(345),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1030_inst_req_0 <= cp_elements(345);
    cp_elements(346) <= cp_elements(267);
    cp_elements(347) <= cp_elements(289);
    cp_elements(348) <= binary_1030_inst_ack_0;
    binary_1030_inst_req_1 <= cp_elements(348);
    cp_elements(349) <= binary_1030_inst_ack_1;
    cpelement_group_350 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(351) & cp_elements(352));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(350),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1036_inst_req_0 <= cp_elements(350);
    cp_elements(351) <= cp_elements(267);
    cp_elements(352) <= cp_elements(289);
    cp_elements(353) <= binary_1036_inst_ack_0;
    binary_1036_inst_req_1 <= cp_elements(353);
    cp_elements(354) <= binary_1036_inst_ack_1;
    cpelement_group_355 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(356) & cp_elements(357));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(355),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1042_inst_req_0 <= cp_elements(355);
    cp_elements(356) <= cp_elements(267);
    cp_elements(357) <= cp_elements(289);
    cp_elements(358) <= binary_1042_inst_ack_0;
    binary_1042_inst_req_1 <= cp_elements(358);
    cp_elements(359) <= binary_1042_inst_ack_1;
    cpelement_group_360 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(359) & cp_elements(361));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(360),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1048_inst_req_0 <= cp_elements(360);
    cp_elements(361) <= cp_elements(267);
    cp_elements(362) <= binary_1048_inst_ack_0;
    binary_1048_inst_req_1 <= cp_elements(362);
    cp_elements(363) <= binary_1048_inst_ack_1;
    cpelement_group_364 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(349) & cp_elements(354) & cp_elements(365));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1053_inst_req_0 <= cp_elements(364);
    cp_elements(365) <= cp_elements(267);
    cp_elements(366) <= binary_1053_inst_ack_0;
    binary_1053_inst_req_1 <= cp_elements(366);
    cp_elements(367) <= binary_1053_inst_ack_1;
    cpelement_group_368 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(367) & cp_elements(369));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(368),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1059_inst_req_0 <= cp_elements(368);
    cp_elements(369) <= cp_elements(267);
    cp_elements(370) <= binary_1059_inst_ack_0;
    binary_1059_inst_req_1 <= cp_elements(370);
    cp_elements(371) <= binary_1059_inst_ack_1;
    cpelement_group_372 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(363) & cp_elements(371) & cp_elements(373));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(372),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1064_inst_req_0 <= cp_elements(372);
    cp_elements(373) <= cp_elements(267);
    cp_elements(374) <= binary_1064_inst_ack_0;
    binary_1064_inst_req_1 <= cp_elements(374);
    cp_elements(375) <= binary_1064_inst_ack_1;
    cpelement_group_376 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(377) & cp_elements(378));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(376),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1070_inst_req_0 <= cp_elements(376);
    cp_elements(377) <= cp_elements(267);
    cp_elements(378) <= cp_elements(295);
    cp_elements(379) <= binary_1070_inst_ack_0;
    binary_1070_inst_req_1 <= cp_elements(379);
    cp_elements(380) <= binary_1070_inst_ack_1;
    cpelement_group_381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(382) & cp_elements(383));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1076_inst_req_0 <= cp_elements(381);
    cp_elements(382) <= cp_elements(267);
    cp_elements(383) <= cp_elements(295);
    cp_elements(384) <= binary_1076_inst_ack_0;
    binary_1076_inst_req_1 <= cp_elements(384);
    cp_elements(385) <= binary_1076_inst_ack_1;
    cpelement_group_386 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(387) & cp_elements(388));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1082_inst_req_0 <= cp_elements(386);
    cp_elements(387) <= cp_elements(267);
    cp_elements(388) <= cp_elements(295);
    cp_elements(389) <= binary_1082_inst_ack_0;
    binary_1082_inst_req_1 <= cp_elements(389);
    cp_elements(390) <= binary_1082_inst_ack_1;
    cpelement_group_391 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(392) & cp_elements(393));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(391),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1088_inst_req_0 <= cp_elements(391);
    cp_elements(392) <= cp_elements(267);
    cp_elements(393) <= cp_elements(295);
    cp_elements(394) <= binary_1088_inst_ack_0;
    binary_1088_inst_req_1 <= cp_elements(394);
    cp_elements(395) <= binary_1088_inst_ack_1;
    cpelement_group_396 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(397) & cp_elements(398));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(396),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1094_inst_req_0 <= cp_elements(396);
    cp_elements(397) <= cp_elements(267);
    cp_elements(398) <= cp_elements(295);
    cp_elements(399) <= binary_1094_inst_ack_0;
    binary_1094_inst_req_1 <= cp_elements(399);
    cp_elements(400) <= binary_1094_inst_ack_1;
    cpelement_group_401 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(400) & cp_elements(402));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(401),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1100_inst_req_0 <= cp_elements(401);
    cp_elements(402) <= cp_elements(267);
    cp_elements(403) <= binary_1100_inst_ack_0;
    binary_1100_inst_req_1 <= cp_elements(403);
    cp_elements(404) <= binary_1100_inst_ack_1;
    cpelement_group_405 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(380) & cp_elements(385) & cp_elements(406));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(405),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1105_inst_req_0 <= cp_elements(405);
    cp_elements(406) <= cp_elements(267);
    cp_elements(407) <= binary_1105_inst_ack_0;
    binary_1105_inst_req_1 <= cp_elements(407);
    cp_elements(408) <= binary_1105_inst_ack_1;
    cpelement_group_409 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(395) & cp_elements(408) & cp_elements(410));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(409),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1110_inst_req_0 <= cp_elements(409);
    cp_elements(410) <= cp_elements(267);
    cp_elements(411) <= binary_1110_inst_ack_0;
    binary_1110_inst_req_1 <= cp_elements(411);
    cp_elements(412) <= binary_1110_inst_ack_1;
    cpelement_group_413 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(390) & cp_elements(412) & cp_elements(414));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(413),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1115_inst_req_0 <= cp_elements(413);
    cp_elements(414) <= cp_elements(267);
    cp_elements(415) <= binary_1115_inst_ack_0;
    binary_1115_inst_req_1 <= cp_elements(415);
    cp_elements(416) <= binary_1115_inst_ack_1;
    cpelement_group_417 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(416) & cp_elements(418));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(417),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1121_inst_req_0 <= cp_elements(417);
    cp_elements(418) <= cp_elements(267);
    cp_elements(419) <= binary_1121_inst_ack_0;
    binary_1121_inst_req_1 <= cp_elements(419);
    cp_elements(420) <= binary_1121_inst_ack_1;
    cpelement_group_421 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(404) & cp_elements(420) & cp_elements(422));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(421),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1126_inst_req_0 <= cp_elements(421);
    cp_elements(422) <= cp_elements(267);
    cp_elements(423) <= binary_1126_inst_ack_0;
    binary_1126_inst_req_1 <= cp_elements(423);
    cp_elements(424) <= binary_1126_inst_ack_1;
    cpelement_group_425 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(426) & cp_elements(427));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(425),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1132_inst_req_0 <= cp_elements(425);
    cp_elements(426) <= cp_elements(267);
    cp_elements(427) <= cp_elements(267);
    cp_elements(428) <= binary_1132_inst_ack_0;
    binary_1132_inst_req_1 <= cp_elements(428);
    cp_elements(429) <= binary_1132_inst_ack_1;
    cpelement_group_430 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(429) & cp_elements(431));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(430),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1138_inst_req_0 <= cp_elements(430);
    cp_elements(431) <= cp_elements(267);
    cp_elements(432) <= binary_1138_inst_ack_0;
    binary_1138_inst_req_1 <= cp_elements(432);
    cp_elements(433) <= binary_1138_inst_ack_1;
    cpelement_group_434 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(344) & cp_elements(375) & cp_elements(424) & cp_elements(433));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(434),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(435) <= cp_elements(7);
    cp_elements(436) <= false;
    cp_elements(437) <= cp_elements(436);
    cp_elements(438) <= cp_elements(7);
    if_stmt_1140_branch_req_0 <= cp_elements(438);
    cp_elements(439) <= cp_elements(438);
    cp_elements(440) <= cp_elements(439);
    cp_elements(441) <= if_stmt_1140_branch_ack_1;
    cp_elements(442) <= cp_elements(439);
    cp_elements(443) <= if_stmt_1140_branch_ack_0;
    cp_elements(444) <= cp_elements(8);
    cp_elements(445) <= cp_elements(444);
    cpelement_group_446 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(445) & cp_elements(447));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(446),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1147_gather_scatter_req_0 <= cp_elements(446);
    cp_elements(447) <= cp_elements(444);
    cp_elements(448) <= simple_obj_ref_1147_gather_scatter_ack_0;
    simple_obj_ref_1147_store_0_req_0 <= cp_elements(448);
    cp_elements(449) <= simple_obj_ref_1147_store_0_ack_0;
    simple_obj_ref_1147_store_0_req_1 <= cp_elements(449);
    cp_elements(450) <= simple_obj_ref_1147_store_0_ack_1;
    cp_elements(451) <= cp_elements(444);
    cpelement_group_452 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(451) & cp_elements(453));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(452),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1150_gather_scatter_req_0 <= cp_elements(452);
    cp_elements(453) <= cp_elements(444);
    cp_elements(454) <= simple_obj_ref_1150_gather_scatter_ack_0;
    simple_obj_ref_1150_store_0_req_0 <= cp_elements(454);
    cp_elements(455) <= simple_obj_ref_1150_store_0_ack_0;
    simple_obj_ref_1150_store_0_req_1 <= cp_elements(455);
    cp_elements(456) <= simple_obj_ref_1150_store_0_ack_1;
    cp_elements(457) <= cp_elements(444);
    cpelement_group_458 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(457) & cp_elements(459));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(458),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1153_gather_scatter_req_0 <= cp_elements(458);
    cp_elements(459) <= cp_elements(444);
    cp_elements(460) <= simple_obj_ref_1153_gather_scatter_ack_0;
    simple_obj_ref_1153_store_0_req_0 <= cp_elements(460);
    cp_elements(461) <= simple_obj_ref_1153_store_0_ack_0;
    simple_obj_ref_1153_store_0_req_1 <= cp_elements(461);
    cp_elements(462) <= simple_obj_ref_1153_store_0_ack_1;
    cpelement_group_463 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(450) & cp_elements(456) & cp_elements(462));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(463),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(464) <= call_stmt_1168_call_ack_0;
    call_stmt_1168_call_req_1 <= cp_elements(464);
    cp_elements(465) <= call_stmt_1168_call_ack_1;
    cp_elements(466) <= cp_elements(465);
    cpelement_group_467 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(468) & cp_elements(469));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(467),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1173_inst_req_0 <= cp_elements(467);
    cp_elements(468) <= cp_elements(466);
    cp_elements(469) <= cp_elements(466);
    cp_elements(470) <= binary_1173_inst_ack_0;
    binary_1173_inst_req_1 <= cp_elements(470);
    cp_elements(471) <= binary_1173_inst_ack_1;
    cpelement_group_472 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(471) & cp_elements(473));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(472),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1179_inst_req_0 <= cp_elements(472);
    cp_elements(473) <= cp_elements(466);
    cp_elements(474) <= binary_1179_inst_ack_0;
    binary_1179_inst_req_1 <= cp_elements(474);
    cp_elements(475) <= binary_1179_inst_ack_1;
    cp_elements(476) <= cp_elements(475);
    cp_elements(477) <= false;
    cp_elements(478) <= cp_elements(477);
    cp_elements(479) <= cp_elements(475);
    if_stmt_1181_branch_req_0 <= cp_elements(479);
    cp_elements(480) <= cp_elements(479);
    cp_elements(481) <= cp_elements(480);
    cp_elements(482) <= if_stmt_1181_branch_ack_1;
    cp_elements(483) <= cp_elements(480);
    cp_elements(484) <= if_stmt_1181_branch_ack_0;
    type_cast_1165_inst_req_0 <= cp_elements(484);
    cp_elements(485) <= cp_elements(224);
    cp_elements(486) <= cp_elements(485);
    type_cast_638_inst_req_0 <= cp_elements(486);
    cp_elements(487) <= type_cast_638_inst_ack_0;
    phi_stmt_632_req_1 <= cp_elements(487);
    cp_elements(488) <= cp_elements(485);
    cp_elements(489) <= cp_elements(488);
    cp_elements(490) <= cp_elements(488);
    type_cast_644_inst_req_0 <= cp_elements(490);
    cp_elements(491) <= type_cast_644_inst_ack_0;
    cpelement_group_492 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(489) & cp_elements(491));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(492),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_639_req_1 <= cp_elements(492);
    cp_elements(493) <= cp_elements(485);
    cp_elements(494) <= cp_elements(493);
    cp_elements(495) <= cp_elements(493);
    type_cast_650_inst_req_0 <= cp_elements(495);
    cp_elements(496) <= type_cast_650_inst_ack_0;
    cpelement_group_497 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(494) & cp_elements(496));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(497),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_645_req_1 <= cp_elements(497);
    cp_elements(498) <= cp_elements(485);
    cp_elements(499) <= cp_elements(498);
    cp_elements(500) <= cp_elements(498);
    type_cast_656_inst_req_0 <= cp_elements(500);
    cp_elements(501) <= type_cast_656_inst_ack_0;
    cpelement_group_502 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(499) & cp_elements(501));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(502),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_651_req_1 <= cp_elements(502);
    cpelement_group_503 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(487) & cp_elements(492) & cp_elements(497) & cp_elements(502));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(503),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(504) <= cp_elements(1);
    cp_elements(505) <= cp_elements(504);
    phi_stmt_632_req_0 <= cp_elements(505);
    cp_elements(506) <= cp_elements(504);
    cp_elements(507) <= cp_elements(506);
    type_cast_642_inst_req_0 <= cp_elements(507);
    cp_elements(508) <= type_cast_642_inst_ack_0;
    cp_elements(509) <= cp_elements(506);
    cpelement_group_510 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(508) & cp_elements(509));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(510),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_639_req_0 <= cp_elements(510);
    cp_elements(511) <= cp_elements(504);
    cp_elements(512) <= cp_elements(511);
    type_cast_648_inst_req_0 <= cp_elements(512);
    cp_elements(513) <= type_cast_648_inst_ack_0;
    cp_elements(514) <= cp_elements(511);
    cpelement_group_515 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(513) & cp_elements(514));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(515),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_645_req_0 <= cp_elements(515);
    cp_elements(516) <= cp_elements(504);
    cp_elements(517) <= cp_elements(516);
    type_cast_654_inst_req_0 <= cp_elements(517);
    cp_elements(518) <= type_cast_654_inst_ack_0;
    cp_elements(519) <= cp_elements(516);
    cpelement_group_520 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(518) & cp_elements(519));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(520),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_651_req_0 <= cp_elements(520);
    cpelement_group_521 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(505) & cp_elements(510) & cp_elements(515) & cp_elements(520));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(521),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(522) <= OrReduce(cp_elements(503) & cp_elements(521));
    cp_elements(523) <= cp_elements(522);
    cp_elements(524) <= phi_stmt_632_ack_0;
    cp_elements(525) <= phi_stmt_639_ack_0;
    cp_elements(526) <= phi_stmt_645_ack_0;
    cp_elements(527) <= phi_stmt_651_ack_0;
    cpelement_group_528 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(524) & cp_elements(525) & cp_elements(526) & cp_elements(527));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(528),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(529) <= false;
    cp_elements(530) <= cp_elements(529);
    cp_elements(531) <= cp_elements(443);
    cp_elements(532) <= cp_elements(531);
    type_cast_918_inst_req_0 <= cp_elements(532);
    cp_elements(533) <= type_cast_918_inst_ack_0;
    phi_stmt_912_req_1 <= cp_elements(533);
    cp_elements(534) <= cp_elements(531);
    cp_elements(535) <= cp_elements(534);
    cp_elements(536) <= cp_elements(534);
    type_cast_924_inst_req_0 <= cp_elements(536);
    cp_elements(537) <= type_cast_924_inst_ack_0;
    cpelement_group_538 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(535) & cp_elements(537));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(538),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_919_req_1 <= cp_elements(538);
    cp_elements(539) <= cp_elements(531);
    cp_elements(540) <= cp_elements(539);
    cp_elements(541) <= cp_elements(539);
    type_cast_930_inst_req_0 <= cp_elements(541);
    cp_elements(542) <= type_cast_930_inst_ack_0;
    cpelement_group_543 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(540) & cp_elements(542));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(543),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_925_req_1 <= cp_elements(543);
    cp_elements(544) <= cp_elements(531);
    cp_elements(545) <= cp_elements(544);
    cp_elements(546) <= cp_elements(544);
    type_cast_936_inst_req_0 <= cp_elements(546);
    cp_elements(547) <= type_cast_936_inst_ack_0;
    cpelement_group_548 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(545) & cp_elements(547));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(548),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_931_req_1 <= cp_elements(548);
    cpelement_group_549 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(533) & cp_elements(538) & cp_elements(543) & cp_elements(548));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(549),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(550) <= cp_elements(5);
    cp_elements(551) <= cp_elements(550);
    phi_stmt_912_req_0 <= cp_elements(551);
    cp_elements(552) <= cp_elements(550);
    cp_elements(553) <= cp_elements(552);
    type_cast_922_inst_req_0 <= cp_elements(553);
    cp_elements(554) <= type_cast_922_inst_ack_0;
    cp_elements(555) <= cp_elements(552);
    cpelement_group_556 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(554) & cp_elements(555));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(556),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_919_req_0 <= cp_elements(556);
    cp_elements(557) <= cp_elements(550);
    cp_elements(558) <= cp_elements(557);
    type_cast_928_inst_req_0 <= cp_elements(558);
    cp_elements(559) <= type_cast_928_inst_ack_0;
    cp_elements(560) <= cp_elements(557);
    cpelement_group_561 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(559) & cp_elements(560));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(561),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_925_req_0 <= cp_elements(561);
    cp_elements(562) <= cp_elements(550);
    cp_elements(563) <= cp_elements(562);
    type_cast_934_inst_req_0 <= cp_elements(563);
    cp_elements(564) <= type_cast_934_inst_ack_0;
    cp_elements(565) <= cp_elements(562);
    cpelement_group_566 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(564) & cp_elements(565));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(566),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_931_req_0 <= cp_elements(566);
    cpelement_group_567 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(551) & cp_elements(556) & cp_elements(561) & cp_elements(566));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(567),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(568) <= OrReduce(cp_elements(549) & cp_elements(567));
    cp_elements(569) <= cp_elements(568);
    cp_elements(570) <= phi_stmt_912_ack_0;
    cp_elements(571) <= phi_stmt_919_ack_0;
    cp_elements(572) <= phi_stmt_925_ack_0;
    cp_elements(573) <= phi_stmt_931_ack_0;
    cpelement_group_574 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(570) & cp_elements(571) & cp_elements(572) & cp_elements(573));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(574),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(575) <= false;
    cp_elements(576) <= cp_elements(575);
    cp_elements(577) <= type_cast_1165_inst_ack_0;
    phi_stmt_1158_req_1 <= cp_elements(577);
    cp_elements(578) <= OrReduce(cp_elements(9) & cp_elements(577));
    cp_elements(579) <= cp_elements(578);
    cp_elements(580) <= phi_stmt_1158_ack_0;
    call_stmt_1168_call_req_0 <= cp_elements(580);
    cp_elements(581) <= false;
    cp_elements(582) <= cp_elements(581);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R1x_xpromoted9_623 : std_logic_vector(31 downto 0);
    signal R1x_xpromoted_903 : std_logic_vector(31 downto 0);
    signal R2x_xpromoted10_626 : std_logic_vector(31 downto 0);
    signal R2x_xpromoted_906 : std_logic_vector(31 downto 0);
    signal R3x_xpromoted11_629 : std_logic_vector(31 downto 0);
    signal R3x_xpromoted_909 : std_logic_vector(31 downto 0);
    signal array_obj_ref_666_final_offset : std_logic_vector(1 downto 0);
    signal array_obj_ref_666_offset_scale_factor_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_666_resized_base_address : std_logic_vector(1 downto 0);
    signal array_obj_ref_666_root_address : std_logic_vector(1 downto 0);
    signal exitcond17_1139 : std_logic_vector(0 downto 0);
    signal exitcond23_881 : std_logic_vector(0 downto 0);
    signal exitcond_1180 : std_logic_vector(0 downto 0);
    signal iNsTr_10_694 : std_logic_vector(31 downto 0);
    signal iNsTr_11_699 : std_logic_vector(31 downto 0);
    signal iNsTr_12_704 : std_logic_vector(31 downto 0);
    signal iNsTr_13_710 : std_logic_vector(31 downto 0);
    signal iNsTr_14_716 : std_logic_vector(31 downto 0);
    signal iNsTr_15_722 : std_logic_vector(31 downto 0);
    signal iNsTr_16_728 : std_logic_vector(31 downto 0);
    signal iNsTr_17_734 : std_logic_vector(31 downto 0);
    signal iNsTr_18_740 : std_logic_vector(31 downto 0);
    signal iNsTr_19_745 : std_logic_vector(31 downto 0);
    signal iNsTr_1_639 : std_logic_vector(31 downto 0);
    signal iNsTr_20_750 : std_logic_vector(31 downto 0);
    signal iNsTr_21_755 : std_logic_vector(31 downto 0);
    signal iNsTr_22_761 : std_logic_vector(31 downto 0);
    signal iNsTr_23_766 : std_logic_vector(31 downto 0);
    signal iNsTr_24_772 : std_logic_vector(31 downto 0);
    signal iNsTr_25_778 : std_logic_vector(31 downto 0);
    signal iNsTr_26_784 : std_logic_vector(31 downto 0);
    signal iNsTr_27_790 : std_logic_vector(31 downto 0);
    signal iNsTr_28_795 : std_logic_vector(31 downto 0);
    signal iNsTr_29_801 : std_logic_vector(31 downto 0);
    signal iNsTr_2_645 : std_logic_vector(31 downto 0);
    signal iNsTr_30_806 : std_logic_vector(31 downto 0);
    signal iNsTr_31_812 : std_logic_vector(31 downto 0);
    signal iNsTr_32_818 : std_logic_vector(31 downto 0);
    signal iNsTr_33_824 : std_logic_vector(31 downto 0);
    signal iNsTr_34_830 : std_logic_vector(31 downto 0);
    signal iNsTr_35_836 : std_logic_vector(31 downto 0);
    signal iNsTr_36_842 : std_logic_vector(31 downto 0);
    signal iNsTr_37_847 : std_logic_vector(31 downto 0);
    signal iNsTr_38_852 : std_logic_vector(31 downto 0);
    signal iNsTr_39_857 : std_logic_vector(31 downto 0);
    signal iNsTr_3_651 : std_logic_vector(31 downto 0);
    signal iNsTr_40_863 : std_logic_vector(31 downto 0);
    signal iNsTr_41_868 : std_logic_vector(31 downto 0);
    signal iNsTr_46_900 : std_logic_vector(31 downto 0);
    signal iNsTr_48_919 : std_logic_vector(31 downto 0);
    signal iNsTr_49_925 : std_logic_vector(31 downto 0);
    signal iNsTr_4_663 : std_logic_vector(31 downto 0);
    signal iNsTr_50_931 : std_logic_vector(31 downto 0);
    signal iNsTr_51_942 : std_logic_vector(31 downto 0);
    signal iNsTr_52_948 : std_logic_vector(31 downto 0);
    signal iNsTr_53_953 : std_logic_vector(31 downto 0);
    signal iNsTr_54_958 : std_logic_vector(31 downto 0);
    signal iNsTr_55_963 : std_logic_vector(31 downto 0);
    signal iNsTr_56_969 : std_logic_vector(31 downto 0);
    signal iNsTr_57_975 : std_logic_vector(31 downto 0);
    signal iNsTr_58_981 : std_logic_vector(31 downto 0);
    signal iNsTr_59_987 : std_logic_vector(31 downto 0);
    signal iNsTr_5_668 : std_logic_vector(31 downto 0);
    signal iNsTr_60_993 : std_logic_vector(31 downto 0);
    signal iNsTr_61_999 : std_logic_vector(31 downto 0);
    signal iNsTr_62_1004 : std_logic_vector(31 downto 0);
    signal iNsTr_63_1009 : std_logic_vector(31 downto 0);
    signal iNsTr_64_1014 : std_logic_vector(31 downto 0);
    signal iNsTr_65_1020 : std_logic_vector(31 downto 0);
    signal iNsTr_66_1025 : std_logic_vector(31 downto 0);
    signal iNsTr_67_1031 : std_logic_vector(31 downto 0);
    signal iNsTr_68_1037 : std_logic_vector(31 downto 0);
    signal iNsTr_69_1043 : std_logic_vector(31 downto 0);
    signal iNsTr_6_672 : std_logic_vector(31 downto 0);
    signal iNsTr_70_1049 : std_logic_vector(31 downto 0);
    signal iNsTr_71_1054 : std_logic_vector(31 downto 0);
    signal iNsTr_72_1060 : std_logic_vector(31 downto 0);
    signal iNsTr_73_1065 : std_logic_vector(31 downto 0);
    signal iNsTr_74_1071 : std_logic_vector(31 downto 0);
    signal iNsTr_75_1077 : std_logic_vector(31 downto 0);
    signal iNsTr_76_1083 : std_logic_vector(31 downto 0);
    signal iNsTr_77_1089 : std_logic_vector(31 downto 0);
    signal iNsTr_78_1095 : std_logic_vector(31 downto 0);
    signal iNsTr_79_1101 : std_logic_vector(31 downto 0);
    signal iNsTr_7_678 : std_logic_vector(31 downto 0);
    signal iNsTr_80_1106 : std_logic_vector(31 downto 0);
    signal iNsTr_81_1111 : std_logic_vector(31 downto 0);
    signal iNsTr_82_1116 : std_logic_vector(31 downto 0);
    signal iNsTr_83_1122 : std_logic_vector(31 downto 0);
    signal iNsTr_84_1127 : std_logic_vector(31 downto 0);
    signal iNsTr_8_683 : std_logic_vector(31 downto 0);
    signal iNsTr_90_1168 : std_logic_vector(31 downto 0);
    signal iNsTr_91_1174 : std_logic_vector(7 downto 0);
    signal iNsTr_9_689 : std_logic_vector(31 downto 0);
    signal indvar21_632 : std_logic_vector(31 downto 0);
    signal indvar_912 : std_logic_vector(31 downto 0);
    signal indvarx_xnext22_874 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1133 : std_logic_vector(31 downto 0);
    signal ix_x21_1158 : std_logic_vector(7 downto 0);
    signal ptr_deref_671_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_671_resized_base_address : std_logic_vector(1 downto 0);
    signal ptr_deref_671_root_address : std_logic_vector(1 downto 0);
    signal ptr_deref_671_word_address_0 : std_logic_vector(1 downto 0);
    signal ptr_deref_671_word_offset_0 : std_logic_vector(1 downto 0);
    signal simple_obj_ref_1147_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1147_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1150_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1150_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1153_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1153_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_622_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_622_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_625_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_625_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_628_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_628_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_665_resized : std_logic_vector(1 downto 0);
    signal simple_obj_ref_665_scaled : std_logic_vector(1 downto 0);
    signal simple_obj_ref_889_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_889_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_892_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_892_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_895_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_895_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_899_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_899_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_902_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_902_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_905_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_905_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_908_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_908_word_address_0 : std_logic_vector(0 downto 0);
    signal type_cast_1018_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1029_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1035_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1041_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1058_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1069_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1081_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1087_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1093_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1099_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1120_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1131_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1137_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1165_wire : std_logic_vector(7 downto 0);
    signal type_cast_1172_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_638_wire : std_logic_vector(31 downto 0);
    signal type_cast_642_wire : std_logic_vector(31 downto 0);
    signal type_cast_644_wire : std_logic_vector(31 downto 0);
    signal type_cast_648_wire : std_logic_vector(31 downto 0);
    signal type_cast_650_wire : std_logic_vector(31 downto 0);
    signal type_cast_654_wire : std_logic_vector(31 downto 0);
    signal type_cast_656_wire : std_logic_vector(31 downto 0);
    signal type_cast_661_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_687_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_708_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_726_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_759_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_770_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_776_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_782_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_799_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_810_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_822_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_834_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_840_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_861_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_918_wire : std_logic_vector(31 downto 0);
    signal type_cast_922_wire : std_logic_vector(31 downto 0);
    signal type_cast_924_wire : std_logic_vector(31 downto 0);
    signal type_cast_928_wire : std_logic_vector(31 downto 0);
    signal type_cast_930_wire : std_logic_vector(31 downto 0);
    signal type_cast_934_wire : std_logic_vector(31 downto 0);
    signal type_cast_936_wire : std_logic_vector(31 downto 0);
    signal type_cast_946_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_967_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_973_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_979_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_985_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_991_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_666_offset_scale_factor_0 <= "01";
    array_obj_ref_666_resized_base_address <= "00";
    ptr_deref_671_word_offset_0 <= "00";
    simple_obj_ref_1147_word_address_0 <= "0";
    simple_obj_ref_1150_word_address_0 <= "0";
    simple_obj_ref_1153_word_address_0 <= "0";
    simple_obj_ref_622_word_address_0 <= "0";
    simple_obj_ref_625_word_address_0 <= "0";
    simple_obj_ref_628_word_address_0 <= "0";
    simple_obj_ref_889_word_address_0 <= "0";
    simple_obj_ref_892_word_address_0 <= "0";
    simple_obj_ref_895_word_address_0 <= "0";
    simple_obj_ref_899_word_address_0 <= "0";
    simple_obj_ref_902_word_address_0 <= "0";
    simple_obj_ref_905_word_address_0 <= "0";
    simple_obj_ref_908_word_address_0 <= "0";
    type_cast_1018_wire_constant <= "00000000000000000000000000000001";
    type_cast_1029_wire_constant <= "00000000000000000000000000010101";
    type_cast_1035_wire_constant <= "00000000000000000000000000010100";
    type_cast_1041_wire_constant <= "00000000000000000000000000000001";
    type_cast_1047_wire_constant <= "00000000001111111111111111111110";
    type_cast_1058_wire_constant <= "00000000000000000000000000000001";
    type_cast_1069_wire_constant <= "00000000000000000000000000010110";
    type_cast_1075_wire_constant <= "00000000000000000000000000010101";
    type_cast_1081_wire_constant <= "00000000000000000000000000010100";
    type_cast_1087_wire_constant <= "00000000000000000000000000000111";
    type_cast_1093_wire_constant <= "00000000000000000000000000000001";
    type_cast_1099_wire_constant <= "00000000011111111111111111111110";
    type_cast_1120_wire_constant <= "00000000000000000000000000000001";
    type_cast_1131_wire_constant <= "00000000000000000000000000000001";
    type_cast_1137_wire_constant <= "00000000000000000000000000010110";
    type_cast_1163_wire_constant <= "00000000";
    type_cast_1172_wire_constant <= "00000001";
    type_cast_1178_wire_constant <= "01100100";
    type_cast_636_wire_constant <= "00000000000000000000000000000000";
    type_cast_661_wire_constant <= "00000000000000000000000000000101";
    type_cast_676_wire_constant <= "00000000000000000000000000011111";
    type_cast_687_wire_constant <= "00000000000000000000000000000001";
    type_cast_708_wire_constant <= "00000000000000000000000000010010";
    type_cast_714_wire_constant <= "00000000000000000000000000010001";
    type_cast_720_wire_constant <= "00000000000000000000000000010000";
    type_cast_726_wire_constant <= "00000000000000000000000000001101";
    type_cast_732_wire_constant <= "00000000000000000000000000000001";
    type_cast_738_wire_constant <= "00000000000001111111111111111110";
    type_cast_759_wire_constant <= "00000000000000000000000000000001";
    type_cast_770_wire_constant <= "00000000000000000000000000010101";
    type_cast_776_wire_constant <= "00000000000000000000000000010100";
    type_cast_782_wire_constant <= "00000000000000000000000000000001";
    type_cast_788_wire_constant <= "00000000001111111111111111111110";
    type_cast_799_wire_constant <= "00000000000000000000000000000001";
    type_cast_810_wire_constant <= "00000000000000000000000000010110";
    type_cast_816_wire_constant <= "00000000000000000000000000010101";
    type_cast_822_wire_constant <= "00000000000000000000000000010100";
    type_cast_828_wire_constant <= "00000000000000000000000000000111";
    type_cast_834_wire_constant <= "00000000000000000000000000000001";
    type_cast_840_wire_constant <= "00000000011111111111111111111110";
    type_cast_861_wire_constant <= "00000000000000000000000000000001";
    type_cast_872_wire_constant <= "00000000000000000000000000000001";
    type_cast_878_wire_constant <= "00000000000000000000000001000000";
    type_cast_916_wire_constant <= "00000000000000000000000000000000";
    type_cast_946_wire_constant <= "00000000000000000000000000000001";
    type_cast_967_wire_constant <= "00000000000000000000000000010010";
    type_cast_973_wire_constant <= "00000000000000000000000000010001";
    type_cast_979_wire_constant <= "00000000000000000000000000010000";
    type_cast_985_wire_constant <= "00000000000000000000000000001101";
    type_cast_991_wire_constant <= "00000000000000000000000000000001";
    type_cast_997_wire_constant <= "00000000000001111111111111111110";
    phi_stmt_1158: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1163_wire_constant & type_cast_1165_wire;
      req <= phi_stmt_1158_req_0 & phi_stmt_1158_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1158_ack_0,
          idata => idata,
          odata => ix_x21_1158,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1158
    phi_stmt_632: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_636_wire_constant & type_cast_638_wire;
      req <= phi_stmt_632_req_0 & phi_stmt_632_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_632_ack_0,
          idata => idata,
          odata => indvar21_632,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_632
    phi_stmt_639: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_642_wire & type_cast_644_wire;
      req <= phi_stmt_639_req_0 & phi_stmt_639_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_639_ack_0,
          idata => idata,
          odata => iNsTr_1_639,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_639
    phi_stmt_645: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_648_wire & type_cast_650_wire;
      req <= phi_stmt_645_req_0 & phi_stmt_645_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_645_ack_0,
          idata => idata,
          odata => iNsTr_2_645,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_645
    phi_stmt_651: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_654_wire & type_cast_656_wire;
      req <= phi_stmt_651_req_0 & phi_stmt_651_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_651_ack_0,
          idata => idata,
          odata => iNsTr_3_651,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_651
    phi_stmt_912: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_916_wire_constant & type_cast_918_wire;
      req <= phi_stmt_912_req_0 & phi_stmt_912_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_912_ack_0,
          idata => idata,
          odata => indvar_912,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_912
    phi_stmt_919: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_922_wire & type_cast_924_wire;
      req <= phi_stmt_919_req_0 & phi_stmt_919_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_919_ack_0,
          idata => idata,
          odata => iNsTr_48_919,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_919
    phi_stmt_925: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_928_wire & type_cast_930_wire;
      req <= phi_stmt_925_req_0 & phi_stmt_925_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_925_ack_0,
          idata => idata,
          odata => iNsTr_49_925,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_925
    phi_stmt_931: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_934_wire & type_cast_936_wire;
      req <= phi_stmt_931_req_0 & phi_stmt_931_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_931_ack_0,
          idata => idata,
          odata => iNsTr_50_931,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_931
    addr_of_667_final_reg: RegisterBase --
      generic map(in_data_width => 2,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_666_root_address, dout => iNsTr_5_668, req => addr_of_667_final_reg_req_0, ack => addr_of_667_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_666_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 2, flow_through => true ) 
      port map( din => iNsTr_4_663, dout => simple_obj_ref_665_resized, req => array_obj_ref_666_index_0_resize_req_0, ack => array_obj_ref_666_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_666_offset_inst: RegisterBase --
      generic map(in_data_width => 2,out_data_width => 2, flow_through => true ) 
      port map( din => simple_obj_ref_665_scaled, dout => array_obj_ref_666_final_offset, req => array_obj_ref_666_offset_inst_req_0, ack => array_obj_ref_666_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_671_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 2, flow_through => true ) 
      port map( din => iNsTr_5_668, dout => ptr_deref_671_resized_base_address, req => ptr_deref_671_base_resize_req_0, ack => ptr_deref_671_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1165_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => iNsTr_91_1174, dout => type_cast_1165_wire, req => type_cast_1165_inst_req_0, ack => type_cast_1165_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_638_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnext22_874, dout => type_cast_638_wire, req => type_cast_638_inst_req_0, ack => type_cast_638_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_642_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => R3x_xpromoted11_629, dout => type_cast_642_wire, req => type_cast_642_inst_req_0, ack => type_cast_642_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_644_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_41_868, dout => type_cast_644_wire, req => type_cast_644_inst_req_0, ack => type_cast_644_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_648_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => R2x_xpromoted10_626, dout => type_cast_648_wire, req => type_cast_648_inst_req_0, ack => type_cast_648_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_650_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_30_806, dout => type_cast_650_wire, req => type_cast_650_inst_req_0, ack => type_cast_650_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_654_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => R1x_xpromoted9_623, dout => type_cast_654_wire, req => type_cast_654_inst_req_0, ack => type_cast_654_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_656_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_23_766, dout => type_cast_656_wire, req => type_cast_656_inst_req_0, ack => type_cast_656_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_918_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnext_1133, dout => type_cast_918_wire, req => type_cast_918_inst_req_0, ack => type_cast_918_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_922_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => R3x_xpromoted_909, dout => type_cast_922_wire, req => type_cast_922_inst_req_0, ack => type_cast_922_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_924_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_84_1127, dout => type_cast_924_wire, req => type_cast_924_inst_req_0, ack => type_cast_924_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_928_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => R2x_xpromoted_906, dout => type_cast_928_wire, req => type_cast_928_inst_req_0, ack => type_cast_928_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_930_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_73_1065, dout => type_cast_930_wire, req => type_cast_930_inst_req_0, ack => type_cast_930_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_934_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => R1x_xpromoted_903, dout => type_cast_934_wire, req => type_cast_934_inst_req_0, ack => type_cast_934_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_936_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_66_1025, dout => type_cast_936_wire, req => type_cast_936_inst_req_0, ack => type_cast_936_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_666_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      array_obj_ref_666_index_0_rename_ack_0 <= array_obj_ref_666_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_665_resized;
      simple_obj_ref_665_scaled <= aggregated_sig(1 downto 0);
      --
    end Block;
    array_obj_ref_666_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      array_obj_ref_666_root_address_inst_ack_0 <= array_obj_ref_666_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_666_final_offset;
      array_obj_ref_666_root_address <= aggregated_sig(1 downto 0);
      --
    end Block;
    ptr_deref_671_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      ptr_deref_671_addr_0_ack_0 <= ptr_deref_671_addr_0_req_0;
      aggregated_sig <= ptr_deref_671_root_address;
      ptr_deref_671_word_address_0 <= aggregated_sig(1 downto 0);
      --
    end Block;
    ptr_deref_671_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_671_gather_scatter_ack_0 <= ptr_deref_671_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_671_data_0;
      iNsTr_6_672 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_671_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      ptr_deref_671_root_address_inst_ack_0 <= ptr_deref_671_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_671_resized_base_address;
      ptr_deref_671_root_address <= aggregated_sig(1 downto 0);
      --
    end Block;
    simple_obj_ref_1147_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1147_gather_scatter_ack_0 <= simple_obj_ref_1147_gather_scatter_req_0;
      aggregated_sig <= iNsTr_84_1127;
      simple_obj_ref_1147_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1150_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1150_gather_scatter_ack_0 <= simple_obj_ref_1150_gather_scatter_req_0;
      aggregated_sig <= iNsTr_73_1065;
      simple_obj_ref_1150_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1153_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1153_gather_scatter_ack_0 <= simple_obj_ref_1153_gather_scatter_req_0;
      aggregated_sig <= iNsTr_66_1025;
      simple_obj_ref_1153_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_622_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_622_gather_scatter_ack_0 <= simple_obj_ref_622_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_622_data_0;
      R1x_xpromoted9_623 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_625_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_625_gather_scatter_ack_0 <= simple_obj_ref_625_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_625_data_0;
      R2x_xpromoted10_626 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_628_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_628_gather_scatter_ack_0 <= simple_obj_ref_628_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_628_data_0;
      R3x_xpromoted11_629 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_889_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_889_gather_scatter_ack_0 <= simple_obj_ref_889_gather_scatter_req_0;
      aggregated_sig <= iNsTr_41_868;
      simple_obj_ref_889_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_892_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_892_gather_scatter_ack_0 <= simple_obj_ref_892_gather_scatter_req_0;
      aggregated_sig <= iNsTr_30_806;
      simple_obj_ref_892_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_895_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_895_gather_scatter_ack_0 <= simple_obj_ref_895_gather_scatter_req_0;
      aggregated_sig <= iNsTr_23_766;
      simple_obj_ref_895_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_899_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_899_gather_scatter_ack_0 <= simple_obj_ref_899_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_899_data_0;
      iNsTr_46_900 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_902_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_902_gather_scatter_ack_0 <= simple_obj_ref_902_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_902_data_0;
      R1x_xpromoted_903 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_905_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_905_gather_scatter_ack_0 <= simple_obj_ref_905_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_905_data_0;
      R2x_xpromoted_906 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_908_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_908_gather_scatter_ack_0 <= simple_obj_ref_908_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_908_data_0;
      R3x_xpromoted_909 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_1140_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond17_1139;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1140_branch_req_0,
          ack0 => if_stmt_1140_branch_ack_0,
          ack1 => if_stmt_1140_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1181_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1180;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1181_branch_req_0,
          ack0 => if_stmt_1181_branch_ack_0,
          ack1 => if_stmt_1181_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_882_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond23_881;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_882_branch_req_0,
          ack0 => if_stmt_882_branch_ack_0,
          ack1 => if_stmt_882_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_1003_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_57_975 & iNsTr_56_969;
      iNsTr_62_1004 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1003_inst_req_0,
          ackL => binary_1003_inst_ack_0,
          reqR => binary_1003_inst_req_1,
          ackR => binary_1003_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_1008_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_62_1004 & iNsTr_59_987;
      iNsTr_63_1009 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1008_inst_req_0,
          ackL => binary_1008_inst_ack_0,
          reqR => binary_1008_inst_req_1,
          ackR => binary_1008_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1013_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_63_1009 & iNsTr_58_981;
      iNsTr_64_1014 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1013_inst_req_0,
          ackL => binary_1013_inst_ack_0,
          reqR => binary_1013_inst_req_1,
          ackR => binary_1013_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1019_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_64_1014;
      iNsTr_65_1020 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1019_inst_req_0,
          ackL => binary_1019_inst_ack_0,
          reqR => binary_1019_inst_req_1,
          ackR => binary_1019_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_1024_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_65_1020 & iNsTr_61_999;
      iNsTr_66_1025 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1024_inst_req_0,
          ackL => binary_1024_inst_ack_0,
          reqR => binary_1024_inst_req_1,
          ackR => binary_1024_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_1030_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_54_958;
      iNsTr_67_1031 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1030_inst_req_0,
          ackL => binary_1030_inst_ack_0,
          reqR => binary_1030_inst_req_1,
          ackR => binary_1030_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_1036_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_54_958;
      iNsTr_68_1037 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1036_inst_req_0,
          ackL => binary_1036_inst_ack_0,
          reqR => binary_1036_inst_req_1,
          ackR => binary_1036_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_1042_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_54_958;
      iNsTr_69_1043 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1042_inst_req_0,
          ackL => binary_1042_inst_ack_0,
          reqR => binary_1042_inst_req_1,
          ackR => binary_1042_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_1048_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_69_1043;
      iNsTr_70_1049 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000001111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1048_inst_req_0,
          ackL => binary_1048_inst_ack_0,
          reqR => binary_1048_inst_req_1,
          ackR => binary_1048_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_1053_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_67_1031 & iNsTr_68_1037;
      iNsTr_71_1054 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1053_inst_req_0,
          ackL => binary_1053_inst_ack_0,
          reqR => binary_1053_inst_req_1,
          ackR => binary_1053_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_1059_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_71_1054;
      iNsTr_72_1060 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1059_inst_req_0,
          ackL => binary_1059_inst_ack_0,
          reqR => binary_1059_inst_req_1,
          ackR => binary_1059_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_1064_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_72_1060 & iNsTr_70_1049;
      iNsTr_73_1065 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1064_inst_req_0,
          ackL => binary_1064_inst_ack_0,
          reqR => binary_1064_inst_req_1,
          ackR => binary_1064_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_1070_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_55_963;
      iNsTr_74_1071 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1070_inst_req_0,
          ackL => binary_1070_inst_ack_0,
          reqR => binary_1070_inst_req_1,
          ackR => binary_1070_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_1076_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_55_963;
      iNsTr_75_1077 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1076_inst_req_0,
          ackL => binary_1076_inst_ack_0,
          reqR => binary_1076_inst_req_1,
          ackR => binary_1076_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_1082_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_55_963;
      iNsTr_76_1083 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1082_inst_req_0,
          ackL => binary_1082_inst_ack_0,
          reqR => binary_1082_inst_req_1,
          ackR => binary_1082_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1088_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_55_963;
      iNsTr_77_1089 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1088_inst_req_0,
          ackL => binary_1088_inst_ack_0,
          reqR => binary_1088_inst_req_1,
          ackR => binary_1088_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1094_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_55_963;
      iNsTr_78_1095 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1094_inst_req_0,
          ackL => binary_1094_inst_ack_0,
          reqR => binary_1094_inst_req_1,
          ackR => binary_1094_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1100_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_78_1095;
      iNsTr_79_1101 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1100_inst_req_0,
          ackL => binary_1100_inst_ack_0,
          reqR => binary_1100_inst_req_1,
          ackR => binary_1100_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1105_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_75_1077 & iNsTr_74_1071;
      iNsTr_80_1106 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1105_inst_req_0,
          ackL => binary_1105_inst_ack_0,
          reqR => binary_1105_inst_req_1,
          ackR => binary_1105_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1110_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_80_1106 & iNsTr_77_1089;
      iNsTr_81_1111 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1110_inst_req_0,
          ackL => binary_1110_inst_ack_0,
          reqR => binary_1110_inst_req_1,
          ackR => binary_1110_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1115_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_81_1111 & iNsTr_76_1083;
      iNsTr_82_1116 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1115_inst_req_0,
          ackL => binary_1115_inst_ack_0,
          reqR => binary_1115_inst_req_1,
          ackR => binary_1115_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1121_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_82_1116;
      iNsTr_83_1122 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1121_inst_req_0,
          ackL => binary_1121_inst_ack_0,
          reqR => binary_1121_inst_req_1,
          ackR => binary_1121_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1126_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_83_1122 & iNsTr_79_1101;
      iNsTr_84_1127 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1126_inst_req_0,
          ackL => binary_1126_inst_ack_0,
          reqR => binary_1126_inst_req_1,
          ackR => binary_1126_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1132_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_912;
      indvarx_xnext_1133 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1132_inst_req_0,
          ackL => binary_1132_inst_ack_0,
          reqR => binary_1132_inst_req_1,
          ackR => binary_1132_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1138_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext_1133;
      exitcond17_1139 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1138_inst_req_0,
          ackL => binary_1138_inst_ack_0,
          reqR => binary_1138_inst_req_1,
          ackR => binary_1138_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1173_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ix_x21_1158;
      iNsTr_91_1174 <= data_out(7 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1173_inst_req_0,
          ackL => binary_1173_inst_ack_0,
          reqR => binary_1173_inst_req_1,
          ackR => binary_1173_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1179_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_91_1174;
      exitcond_1180 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01100100",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1179_inst_req_0,
          ackL => binary_1179_inst_ack_0,
          reqR => binary_1179_inst_req_1,
          ackR => binary_1179_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_662_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar21_632;
      iNsTr_4_663 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_662_inst_req_0,
          ackL => binary_662_inst_ack_0,
          reqR => binary_662_inst_req_1,
          ackR => binary_662_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_677_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar21_632;
      iNsTr_7_678 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000011111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_677_inst_req_0,
          ackL => binary_677_inst_ack_0,
          reqR => binary_677_inst_req_1,
          ackR => binary_677_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_682_inst binary_941_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_6_672 & iNsTr_7_678 & iNsTr_46_900 & indvar_912;
      iNsTr_8_683 <= data_out(63 downto 32);
      iNsTr_51_942 <= data_out(31 downto 0);
      reqL(1) <= binary_682_inst_req_0;
      reqL(0) <= binary_941_inst_req_0;
      binary_682_inst_ack_0 <= ackL(1);
      binary_941_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_682_inst_req_1;
      reqR(0) <= binary_941_inst_req_1;
      binary_682_inst_ack_1 <= ackR(1);
      binary_941_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_688_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_8_683;
      iNsTr_9_689 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_688_inst_req_0,
          ackL => binary_688_inst_ack_0,
          reqR => binary_688_inst_req_1,
          ackR => binary_688_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_693_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_689 & iNsTr_3_651;
      iNsTr_10_694 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_693_inst_req_0,
          ackL => binary_693_inst_ack_0,
          reqR => binary_693_inst_req_1,
          ackR => binary_693_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_698_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_645 & iNsTr_9_689;
      iNsTr_11_699 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_698_inst_req_0,
          ackL => binary_698_inst_ack_0,
          reqR => binary_698_inst_req_1,
          ackR => binary_698_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_703_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_1_639 & iNsTr_9_689;
      iNsTr_12_704 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_703_inst_req_0,
          ackL => binary_703_inst_ack_0,
          reqR => binary_703_inst_req_1,
          ackR => binary_703_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_709_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_694;
      iNsTr_13_710 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_709_inst_req_0,
          ackL => binary_709_inst_ack_0,
          reqR => binary_709_inst_req_1,
          ackR => binary_709_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_715_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_694;
      iNsTr_14_716 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_715_inst_req_0,
          ackL => binary_715_inst_ack_0,
          reqR => binary_715_inst_req_1,
          ackR => binary_715_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_721_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_694;
      iNsTr_15_722 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_721_inst_req_0,
          ackL => binary_721_inst_ack_0,
          reqR => binary_721_inst_req_1,
          ackR => binary_721_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_727_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_694;
      iNsTr_16_728 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_727_inst_req_0,
          ackL => binary_727_inst_ack_0,
          reqR => binary_727_inst_req_1,
          ackR => binary_727_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_733_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_694;
      iNsTr_17_734 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_733_inst_req_0,
          ackL => binary_733_inst_ack_0,
          reqR => binary_733_inst_req_1,
          ackR => binary_733_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_739_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_17_734;
      iNsTr_18_740 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000001111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_739_inst_req_0,
          ackL => binary_739_inst_ack_0,
          reqR => binary_739_inst_req_1,
          ackR => binary_739_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_744_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_14_716 & iNsTr_13_710;
      iNsTr_19_745 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_744_inst_req_0,
          ackL => binary_744_inst_ack_0,
          reqR => binary_744_inst_req_1,
          ackR => binary_744_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_749_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_19_745 & iNsTr_16_728;
      iNsTr_20_750 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_749_inst_req_0,
          ackL => binary_749_inst_ack_0,
          reqR => binary_749_inst_req_1,
          ackR => binary_749_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_754_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_20_750 & iNsTr_15_722;
      iNsTr_21_755 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_754_inst_req_0,
          ackL => binary_754_inst_ack_0,
          reqR => binary_754_inst_req_1,
          ackR => binary_754_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_760_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_21_755;
      iNsTr_22_761 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_760_inst_req_0,
          ackL => binary_760_inst_ack_0,
          reqR => binary_760_inst_req_1,
          ackR => binary_760_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_765_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_22_761 & iNsTr_18_740;
      iNsTr_23_766 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_765_inst_req_0,
          ackL => binary_765_inst_ack_0,
          reqR => binary_765_inst_req_1,
          ackR => binary_765_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_771_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_11_699;
      iNsTr_24_772 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_771_inst_req_0,
          ackL => binary_771_inst_ack_0,
          reqR => binary_771_inst_req_1,
          ackR => binary_771_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_777_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_11_699;
      iNsTr_25_778 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_777_inst_req_0,
          ackL => binary_777_inst_ack_0,
          reqR => binary_777_inst_req_1,
          ackR => binary_777_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_783_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_11_699;
      iNsTr_26_784 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_783_inst_req_0,
          ackL => binary_783_inst_ack_0,
          reqR => binary_783_inst_req_1,
          ackR => binary_783_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_789_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_26_784;
      iNsTr_27_790 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000001111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_789_inst_req_0,
          ackL => binary_789_inst_ack_0,
          reqR => binary_789_inst_req_1,
          ackR => binary_789_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_794_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_24_772 & iNsTr_25_778;
      iNsTr_28_795 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_794_inst_req_0,
          ackL => binary_794_inst_ack_0,
          reqR => binary_794_inst_req_1,
          ackR => binary_794_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_800_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_28_795;
      iNsTr_29_801 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_800_inst_req_0,
          ackL => binary_800_inst_ack_0,
          reqR => binary_800_inst_req_1,
          ackR => binary_800_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_805_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_29_801 & iNsTr_27_790;
      iNsTr_30_806 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_805_inst_req_0,
          ackL => binary_805_inst_ack_0,
          reqR => binary_805_inst_req_1,
          ackR => binary_805_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_811_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_704;
      iNsTr_31_812 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_811_inst_req_0,
          ackL => binary_811_inst_ack_0,
          reqR => binary_811_inst_req_1,
          ackR => binary_811_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_817_inst 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_704;
      iNsTr_32_818 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_817_inst_req_0,
          ackL => binary_817_inst_ack_0,
          reqR => binary_817_inst_req_1,
          ackR => binary_817_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : binary_823_inst 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_704;
      iNsTr_33_824 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_823_inst_req_0,
          ackL => binary_823_inst_ack_0,
          reqR => binary_823_inst_req_1,
          ackR => binary_823_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : binary_829_inst 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_704;
      iNsTr_34_830 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_829_inst_req_0,
          ackL => binary_829_inst_ack_0,
          reqR => binary_829_inst_req_1,
          ackR => binary_829_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : binary_835_inst 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_704;
      iNsTr_35_836 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_835_inst_req_0,
          ackL => binary_835_inst_ack_0,
          reqR => binary_835_inst_req_1,
          ackR => binary_835_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : binary_841_inst 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_35_836;
      iNsTr_36_842 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_841_inst_req_0,
          ackL => binary_841_inst_ack_0,
          reqR => binary_841_inst_req_1,
          ackR => binary_841_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : binary_846_inst 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_32_818 & iNsTr_31_812;
      iNsTr_37_847 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_846_inst_req_0,
          ackL => binary_846_inst_ack_0,
          reqR => binary_846_inst_req_1,
          ackR => binary_846_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : binary_851_inst 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_37_847 & iNsTr_34_830;
      iNsTr_38_852 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_851_inst_req_0,
          ackL => binary_851_inst_ack_0,
          reqR => binary_851_inst_req_1,
          ackR => binary_851_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : binary_856_inst 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_38_852 & iNsTr_33_824;
      iNsTr_39_857 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_856_inst_req_0,
          ackL => binary_856_inst_ack_0,
          reqR => binary_856_inst_req_1,
          ackR => binary_856_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : binary_862_inst 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_39_857;
      iNsTr_40_863 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_862_inst_req_0,
          ackL => binary_862_inst_ack_0,
          reqR => binary_862_inst_req_1,
          ackR => binary_862_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : binary_867_inst 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_40_863 & iNsTr_36_842;
      iNsTr_41_868 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_867_inst_req_0,
          ackL => binary_867_inst_ack_0,
          reqR => binary_867_inst_req_1,
          ackR => binary_867_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : binary_873_inst 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar21_632;
      indvarx_xnext22_874 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_873_inst_req_0,
          ackL => binary_873_inst_ack_0,
          reqR => binary_873_inst_req_1,
          ackR => binary_873_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : binary_879_inst 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext22_874;
      exitcond23_881 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_879_inst_req_0,
          ackL => binary_879_inst_ack_0,
          reqR => binary_879_inst_req_1,
          ackR => binary_879_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : binary_947_inst 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_51_942;
      iNsTr_52_948 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_947_inst_req_0,
          ackL => binary_947_inst_ack_0,
          reqR => binary_947_inst_req_1,
          ackR => binary_947_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : binary_952_inst 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_52_948 & iNsTr_50_931;
      iNsTr_53_953 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_952_inst_req_0,
          ackL => binary_952_inst_ack_0,
          reqR => binary_952_inst_req_1,
          ackR => binary_952_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : binary_957_inst 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_49_925 & iNsTr_52_948;
      iNsTr_54_958 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_957_inst_req_0,
          ackL => binary_957_inst_ack_0,
          reqR => binary_957_inst_req_1,
          ackR => binary_957_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : binary_962_inst 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_48_919 & iNsTr_52_948;
      iNsTr_55_963 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_962_inst_req_0,
          ackL => binary_962_inst_ack_0,
          reqR => binary_962_inst_req_1,
          ackR => binary_962_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : binary_968_inst 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_53_953;
      iNsTr_56_969 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_968_inst_req_0,
          ackL => binary_968_inst_ack_0,
          reqR => binary_968_inst_req_1,
          ackR => binary_968_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : binary_974_inst 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_53_953;
      iNsTr_57_975 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_974_inst_req_0,
          ackL => binary_974_inst_ack_0,
          reqR => binary_974_inst_req_1,
          ackR => binary_974_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : binary_980_inst 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_53_953;
      iNsTr_58_981 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_980_inst_req_0,
          ackL => binary_980_inst_ack_0,
          reqR => binary_980_inst_req_1,
          ackR => binary_980_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : binary_986_inst 
    SplitOperatorGroup72: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_53_953;
      iNsTr_59_987 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_986_inst_req_0,
          ackL => binary_986_inst_ack_0,
          reqR => binary_986_inst_req_1,
          ackR => binary_986_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : binary_992_inst 
    SplitOperatorGroup73: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_53_953;
      iNsTr_60_993 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_992_inst_req_0,
          ackL => binary_992_inst_ack_0,
          reqR => binary_992_inst_req_1,
          ackR => binary_992_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : binary_998_inst 
    SplitOperatorGroup74: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_60_993;
      iNsTr_61_999 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000001111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_998_inst_req_0,
          ackL => binary_998_inst_ack_0,
          reqR => binary_998_inst_req_1,
          ackR => binary_998_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared load operator group (0) : ptr_deref_671_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_671_load_0_req_0;
      ptr_deref_671_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_671_load_0_req_1;
      ptr_deref_671_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_671_word_address_0;
      ptr_deref_671_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 2,  num_reqs => 1,  tag_length => 1, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(1 downto 0),
          mtag => memory_space_3_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : simple_obj_ref_622_load_0 simple_obj_ref_902_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= simple_obj_ref_622_load_0_req_0;
      reqL(0) <= simple_obj_ref_902_load_0_req_0;
      simple_obj_ref_622_load_0_ack_0 <= ackL(1);
      simple_obj_ref_902_load_0_ack_0 <= ackL(0);
      reqR(1) <= simple_obj_ref_622_load_0_req_1;
      reqR(0) <= simple_obj_ref_902_load_0_req_1;
      simple_obj_ref_622_load_0_ack_1 <= ackR(1);
      simple_obj_ref_902_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_622_word_address_0 & simple_obj_ref_902_word_address_0;
      simple_obj_ref_622_data_0 <= data_out(63 downto 32);
      simple_obj_ref_902_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : simple_obj_ref_625_load_0 simple_obj_ref_905_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= simple_obj_ref_625_load_0_req_0;
      reqL(0) <= simple_obj_ref_905_load_0_req_0;
      simple_obj_ref_625_load_0_ack_0 <= ackL(1);
      simple_obj_ref_905_load_0_ack_0 <= ackL(0);
      reqR(1) <= simple_obj_ref_625_load_0_req_1;
      reqR(0) <= simple_obj_ref_905_load_0_req_1;
      simple_obj_ref_625_load_0_ack_1 <= ackR(1);
      simple_obj_ref_905_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_625_word_address_0 & simple_obj_ref_905_word_address_0;
      simple_obj_ref_625_data_0 <= data_out(63 downto 32);
      simple_obj_ref_905_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : simple_obj_ref_628_load_0 simple_obj_ref_908_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= simple_obj_ref_628_load_0_req_0;
      reqL(0) <= simple_obj_ref_908_load_0_req_0;
      simple_obj_ref_628_load_0_ack_0 <= ackL(1);
      simple_obj_ref_908_load_0_ack_0 <= ackL(0);
      reqR(1) <= simple_obj_ref_628_load_0_req_1;
      reqR(0) <= simple_obj_ref_908_load_0_req_1;
      simple_obj_ref_628_load_0_ack_1 <= ackR(1);
      simple_obj_ref_908_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_628_word_address_0 & simple_obj_ref_908_word_address_0;
      simple_obj_ref_628_data_0 <= data_out(63 downto 32);
      simple_obj_ref_908_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : simple_obj_ref_899_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_899_load_0_req_0;
      simple_obj_ref_899_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_899_load_0_req_1;
      simple_obj_ref_899_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_899_word_address_0;
      simple_obj_ref_899_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared store operator group (0) : simple_obj_ref_889_store_0 simple_obj_ref_1147_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= simple_obj_ref_889_store_0_req_0;
      reqL(0) <= simple_obj_ref_1147_store_0_req_0;
      simple_obj_ref_889_store_0_ack_0 <= ackL(1);
      simple_obj_ref_1147_store_0_ack_0 <= ackL(0);
      reqR(1) <= simple_obj_ref_889_store_0_req_1;
      reqR(0) <= simple_obj_ref_1147_store_0_req_1;
      simple_obj_ref_889_store_0_ack_1 <= ackR(1);
      simple_obj_ref_1147_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_889_word_address_0 & simple_obj_ref_1147_word_address_0;
      data_in <= simple_obj_ref_889_data_0 & simple_obj_ref_1147_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : simple_obj_ref_892_store_0 simple_obj_ref_1150_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= simple_obj_ref_892_store_0_req_0;
      reqL(0) <= simple_obj_ref_1150_store_0_req_0;
      simple_obj_ref_892_store_0_ack_0 <= ackL(1);
      simple_obj_ref_1150_store_0_ack_0 <= ackL(0);
      reqR(1) <= simple_obj_ref_892_store_0_req_1;
      reqR(0) <= simple_obj_ref_1150_store_0_req_1;
      simple_obj_ref_892_store_0_ack_1 <= ackR(1);
      simple_obj_ref_1150_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_892_word_address_0 & simple_obj_ref_1150_word_address_0;
      data_in <= simple_obj_ref_892_data_0 & simple_obj_ref_1150_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : simple_obj_ref_895_store_0 simple_obj_ref_1153_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= simple_obj_ref_895_store_0_req_0;
      reqL(0) <= simple_obj_ref_1153_store_0_req_0;
      simple_obj_ref_895_store_0_ack_0 <= ackL(1);
      simple_obj_ref_1153_store_0_ack_0 <= ackL(0);
      reqR(1) <= simple_obj_ref_895_store_0_req_1;
      reqR(0) <= simple_obj_ref_1153_store_0_req_1;
      simple_obj_ref_895_store_0_ack_1 <= ackR(1);
      simple_obj_ref_1153_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_895_word_address_0 & simple_obj_ref_1153_word_address_0;
      data_in <= simple_obj_ref_895_data_0 & simple_obj_ref_1153_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared call operator group (0) : call_stmt_1168_call 
    CallGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1168_call_req_0;
      call_stmt_1168_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1168_call_req_1;
      call_stmt_1168_call_ack_1 <= ackR(0);
      iNsTr_90_1168 <= data_out(31 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => a5reg_call_reqs(0),
          ackR => a5reg_call_acks(0),
          tagR => a5reg_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 32, owidth => 32, twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => a5reg_return_acks(0), -- cross-over
          ackL => a5reg_return_reqs(0), -- cross-over
          dataL => a5reg_return_data(31 downto 0),
          tagL => a5reg_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity a5reg is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(31 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity a5reg;
architecture Default of a5reg is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(31 downto 0);
  signal a5reg_CP_0_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_15_load_0_req_0 : boolean;
  signal simple_obj_ref_15_load_0_ack_0 : boolean;
  signal simple_obj_ref_15_load_0_req_1 : boolean;
  signal simple_obj_ref_15_load_0_ack_1 : boolean;
  signal simple_obj_ref_15_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_15_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_12_load_0_req_0 : boolean;
  signal simple_obj_ref_12_load_0_ack_0 : boolean;
  signal simple_obj_ref_12_load_0_req_1 : boolean;
  signal simple_obj_ref_12_load_0_ack_1 : boolean;
  signal simple_obj_ref_12_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_12_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_18_load_0_req_0 : boolean;
  signal simple_obj_ref_18_load_0_ack_0 : boolean;
  signal simple_obj_ref_18_load_0_req_1 : boolean;
  signal simple_obj_ref_18_load_0_ack_1 : boolean;
  signal simple_obj_ref_18_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_18_gather_scatter_ack_0 : boolean;
  signal binary_24_inst_req_0 : boolean;
  signal binary_24_inst_ack_0 : boolean;
  signal binary_24_inst_req_1 : boolean;
  signal binary_24_inst_ack_1 : boolean;
  signal binary_30_inst_req_0 : boolean;
  signal binary_30_inst_ack_0 : boolean;
  signal binary_30_inst_req_1 : boolean;
  signal binary_30_inst_ack_1 : boolean;
  signal binary_36_inst_req_0 : boolean;
  signal binary_36_inst_ack_0 : boolean;
  signal binary_36_inst_req_1 : boolean;
  signal binary_36_inst_ack_1 : boolean;
  signal binary_42_inst_req_0 : boolean;
  signal binary_42_inst_ack_0 : boolean;
  signal binary_42_inst_req_1 : boolean;
  signal binary_42_inst_ack_1 : boolean;
  signal binary_48_inst_req_0 : boolean;
  signal binary_48_inst_ack_0 : boolean;
  signal binary_48_inst_req_1 : boolean;
  signal binary_48_inst_ack_1 : boolean;
  signal binary_54_inst_req_0 : boolean;
  signal binary_54_inst_ack_0 : boolean;
  signal binary_54_inst_req_1 : boolean;
  signal binary_54_inst_ack_1 : boolean;
  signal binary_125_inst_req_1 : boolean;
  signal binary_125_inst_ack_1 : boolean;
  signal binary_60_inst_req_0 : boolean;
  signal binary_60_inst_ack_0 : boolean;
  signal binary_60_inst_req_1 : boolean;
  signal simple_obj_ref_424_store_0_ack_1 : boolean;
  signal binary_60_inst_ack_1 : boolean;
  signal binary_66_inst_req_0 : boolean;
  signal binary_66_inst_ack_0 : boolean;
  signal binary_66_inst_req_1 : boolean;
  signal simple_obj_ref_424_store_0_req_1 : boolean;
  signal binary_66_inst_ack_1 : boolean;
  signal binary_72_inst_req_0 : boolean;
  signal binary_72_inst_ack_0 : boolean;
  signal binary_72_inst_req_1 : boolean;
  signal binary_72_inst_ack_1 : boolean;
  signal binary_78_inst_req_0 : boolean;
  signal binary_78_inst_ack_0 : boolean;
  signal binary_78_inst_req_1 : boolean;
  signal binary_78_inst_ack_1 : boolean;
  signal binary_84_inst_req_0 : boolean;
  signal binary_84_inst_ack_0 : boolean;
  signal binary_84_inst_req_1 : boolean;
  signal binary_84_inst_ack_1 : boolean;
  signal binary_89_inst_req_0 : boolean;
  signal binary_89_inst_ack_0 : boolean;
  signal binary_89_inst_req_1 : boolean;
  signal binary_89_inst_ack_1 : boolean;
  signal binary_95_inst_req_0 : boolean;
  signal binary_95_inst_ack_0 : boolean;
  signal binary_95_inst_req_1 : boolean;
  signal binary_95_inst_ack_1 : boolean;
  signal binary_100_inst_req_0 : boolean;
  signal binary_100_inst_ack_0 : boolean;
  signal binary_100_inst_req_1 : boolean;
  signal binary_100_inst_ack_1 : boolean;
  signal binary_105_inst_req_0 : boolean;
  signal binary_105_inst_ack_0 : boolean;
  signal binary_105_inst_req_1 : boolean;
  signal simple_obj_ref_424_store_0_ack_0 : boolean;
  signal binary_105_inst_ack_1 : boolean;
  signal binary_110_inst_req_0 : boolean;
  signal binary_110_inst_ack_0 : boolean;
  signal binary_110_inst_req_1 : boolean;
  signal simple_obj_ref_424_store_0_req_0 : boolean;
  signal binary_110_inst_ack_1 : boolean;
  signal binary_115_inst_req_0 : boolean;
  signal binary_115_inst_ack_0 : boolean;
  signal binary_115_inst_req_1 : boolean;
  signal binary_115_inst_ack_1 : boolean;
  signal binary_120_inst_req_0 : boolean;
  signal binary_120_inst_ack_0 : boolean;
  signal binary_120_inst_req_1 : boolean;
  signal binary_120_inst_ack_1 : boolean;
  signal binary_125_inst_req_0 : boolean;
  signal binary_125_inst_ack_0 : boolean;
  signal binary_275_inst_req_0 : boolean;
  signal binary_275_inst_ack_0 : boolean;
  signal binary_275_inst_req_1 : boolean;
  signal binary_275_inst_ack_1 : boolean;
  signal binary_281_inst_req_0 : boolean;
  signal binary_281_inst_ack_0 : boolean;
  signal binary_281_inst_req_1 : boolean;
  signal binary_281_inst_ack_1 : boolean;
  signal binary_130_inst_req_0 : boolean;
  signal binary_130_inst_ack_0 : boolean;
  signal binary_130_inst_req_1 : boolean;
  signal binary_130_inst_ack_1 : boolean;
  signal binary_135_inst_req_0 : boolean;
  signal binary_135_inst_ack_0 : boolean;
  signal binary_135_inst_req_1 : boolean;
  signal simple_obj_ref_424_gather_scatter_ack_0 : boolean;
  signal binary_135_inst_ack_1 : boolean;
  signal binary_140_inst_req_0 : boolean;
  signal binary_140_inst_ack_0 : boolean;
  signal binary_140_inst_req_1 : boolean;
  signal simple_obj_ref_424_gather_scatter_req_0 : boolean;
  signal binary_140_inst_ack_1 : boolean;
  signal binary_145_inst_req_0 : boolean;
  signal binary_145_inst_ack_0 : boolean;
  signal binary_145_inst_req_1 : boolean;
  signal binary_145_inst_ack_1 : boolean;
  signal binary_150_inst_req_0 : boolean;
  signal binary_150_inst_ack_0 : boolean;
  signal binary_150_inst_req_1 : boolean;
  signal binary_150_inst_ack_1 : boolean;
  signal binary_155_inst_req_0 : boolean;
  signal binary_155_inst_ack_0 : boolean;
  signal binary_155_inst_req_1 : boolean;
  signal binary_155_inst_ack_1 : boolean;
  signal binary_161_inst_req_0 : boolean;
  signal binary_161_inst_ack_0 : boolean;
  signal binary_161_inst_req_1 : boolean;
  signal binary_161_inst_ack_1 : boolean;
  signal binary_167_inst_req_0 : boolean;
  signal binary_167_inst_ack_0 : boolean;
  signal binary_167_inst_req_1 : boolean;
  signal binary_167_inst_ack_1 : boolean;
  signal binary_173_inst_req_0 : boolean;
  signal binary_173_inst_ack_0 : boolean;
  signal binary_173_inst_req_1 : boolean;
  signal binary_173_inst_ack_1 : boolean;
  signal binary_179_inst_req_0 : boolean;
  signal binary_179_inst_ack_0 : boolean;
  signal binary_179_inst_req_1 : boolean;
  signal binary_179_inst_ack_1 : boolean;
  signal binary_184_inst_req_0 : boolean;
  signal binary_184_inst_ack_0 : boolean;
  signal binary_184_inst_req_1 : boolean;
  signal binary_184_inst_ack_1 : boolean;
  signal binary_189_inst_req_0 : boolean;
  signal binary_189_inst_ack_0 : boolean;
  signal binary_189_inst_req_1 : boolean;
  signal binary_189_inst_ack_1 : boolean;
  signal binary_194_inst_req_0 : boolean;
  signal binary_194_inst_ack_0 : boolean;
  signal binary_194_inst_req_1 : boolean;
  signal binary_194_inst_ack_1 : boolean;
  signal binary_200_inst_req_0 : boolean;
  signal binary_200_inst_ack_0 : boolean;
  signal binary_200_inst_req_1 : boolean;
  signal binary_200_inst_ack_1 : boolean;
  signal binary_206_inst_req_0 : boolean;
  signal binary_206_inst_ack_0 : boolean;
  signal binary_206_inst_req_1 : boolean;
  signal binary_206_inst_ack_1 : boolean;
  signal binary_212_inst_req_0 : boolean;
  signal binary_212_inst_ack_0 : boolean;
  signal binary_212_inst_req_1 : boolean;
  signal binary_212_inst_ack_1 : boolean;
  signal binary_217_inst_req_0 : boolean;
  signal binary_217_inst_ack_0 : boolean;
  signal binary_217_inst_req_1 : boolean;
  signal binary_217_inst_ack_1 : boolean;
  signal binary_223_inst_req_0 : boolean;
  signal binary_223_inst_ack_0 : boolean;
  signal binary_223_inst_req_1 : boolean;
  signal binary_223_inst_ack_1 : boolean;
  signal binary_229_inst_req_0 : boolean;
  signal binary_229_inst_ack_0 : boolean;
  signal binary_229_inst_req_1 : boolean;
  signal binary_229_inst_ack_1 : boolean;
  signal binary_234_inst_req_0 : boolean;
  signal binary_234_inst_ack_0 : boolean;
  signal binary_234_inst_req_1 : boolean;
  signal binary_234_inst_ack_1 : boolean;
  signal binary_240_inst_req_0 : boolean;
  signal binary_240_inst_ack_0 : boolean;
  signal binary_240_inst_req_1 : boolean;
  signal binary_240_inst_ack_1 : boolean;
  signal binary_246_inst_req_0 : boolean;
  signal binary_246_inst_ack_0 : boolean;
  signal binary_246_inst_req_1 : boolean;
  signal binary_246_inst_ack_1 : boolean;
  signal binary_252_inst_req_0 : boolean;
  signal binary_252_inst_ack_0 : boolean;
  signal binary_252_inst_req_1 : boolean;
  signal binary_252_inst_ack_1 : boolean;
  signal binary_257_inst_req_0 : boolean;
  signal binary_257_inst_ack_0 : boolean;
  signal binary_257_inst_req_1 : boolean;
  signal binary_257_inst_ack_1 : boolean;
  signal binary_263_inst_req_0 : boolean;
  signal binary_263_inst_ack_0 : boolean;
  signal binary_263_inst_req_1 : boolean;
  signal binary_263_inst_ack_1 : boolean;
  signal binary_269_inst_req_0 : boolean;
  signal binary_269_inst_ack_0 : boolean;
  signal binary_269_inst_req_1 : boolean;
  signal binary_269_inst_ack_1 : boolean;
  signal binary_286_inst_req_0 : boolean;
  signal binary_286_inst_ack_0 : boolean;
  signal binary_286_inst_req_1 : boolean;
  signal binary_286_inst_ack_1 : boolean;
  signal binary_291_inst_req_0 : boolean;
  signal binary_291_inst_ack_0 : boolean;
  signal binary_291_inst_req_1 : boolean;
  signal binary_291_inst_ack_1 : boolean;
  signal binary_296_inst_req_0 : boolean;
  signal binary_296_inst_ack_0 : boolean;
  signal binary_296_inst_req_1 : boolean;
  signal binary_296_inst_ack_1 : boolean;
  signal binary_302_inst_req_0 : boolean;
  signal binary_302_inst_ack_0 : boolean;
  signal binary_302_inst_req_1 : boolean;
  signal binary_302_inst_ack_1 : boolean;
  signal binary_308_inst_req_0 : boolean;
  signal binary_308_inst_ack_0 : boolean;
  signal binary_308_inst_req_1 : boolean;
  signal binary_308_inst_ack_1 : boolean;
  signal binary_314_inst_req_0 : boolean;
  signal binary_314_inst_ack_0 : boolean;
  signal binary_314_inst_req_1 : boolean;
  signal binary_314_inst_ack_1 : boolean;
  signal binary_319_inst_req_0 : boolean;
  signal binary_319_inst_ack_0 : boolean;
  signal binary_319_inst_req_1 : boolean;
  signal binary_319_inst_ack_1 : boolean;
  signal binary_324_inst_req_0 : boolean;
  signal binary_324_inst_ack_0 : boolean;
  signal binary_324_inst_req_1 : boolean;
  signal binary_324_inst_ack_1 : boolean;
  signal binary_330_inst_req_0 : boolean;
  signal binary_330_inst_ack_0 : boolean;
  signal binary_330_inst_req_1 : boolean;
  signal binary_330_inst_ack_1 : boolean;
  signal binary_335_inst_req_0 : boolean;
  signal binary_335_inst_ack_0 : boolean;
  signal binary_335_inst_req_1 : boolean;
  signal binary_335_inst_ack_1 : boolean;
  signal binary_340_inst_req_0 : boolean;
  signal binary_340_inst_ack_0 : boolean;
  signal binary_340_inst_req_1 : boolean;
  signal binary_340_inst_ack_1 : boolean;
  signal binary_345_inst_req_0 : boolean;
  signal binary_345_inst_ack_0 : boolean;
  signal binary_345_inst_req_1 : boolean;
  signal binary_345_inst_ack_1 : boolean;
  signal binary_351_inst_req_0 : boolean;
  signal binary_351_inst_ack_0 : boolean;
  signal binary_351_inst_req_1 : boolean;
  signal binary_351_inst_ack_1 : boolean;
  signal binary_356_inst_req_0 : boolean;
  signal binary_356_inst_ack_0 : boolean;
  signal binary_356_inst_req_1 : boolean;
  signal binary_356_inst_ack_1 : boolean;
  signal binary_361_inst_req_0 : boolean;
  signal binary_361_inst_ack_0 : boolean;
  signal binary_361_inst_req_1 : boolean;
  signal binary_361_inst_ack_1 : boolean;
  signal binary_366_inst_req_0 : boolean;
  signal binary_366_inst_ack_0 : boolean;
  signal binary_366_inst_req_1 : boolean;
  signal binary_366_inst_ack_1 : boolean;
  signal binary_372_inst_req_0 : boolean;
  signal binary_372_inst_ack_0 : boolean;
  signal binary_372_inst_req_1 : boolean;
  signal binary_372_inst_ack_1 : boolean;
  signal binary_377_inst_req_0 : boolean;
  signal binary_377_inst_ack_0 : boolean;
  signal binary_377_inst_req_1 : boolean;
  signal binary_377_inst_ack_1 : boolean;
  signal binary_382_inst_req_0 : boolean;
  signal binary_382_inst_ack_0 : boolean;
  signal binary_382_inst_req_1 : boolean;
  signal binary_382_inst_ack_1 : boolean;
  signal binary_388_inst_req_0 : boolean;
  signal binary_388_inst_ack_0 : boolean;
  signal binary_388_inst_req_1 : boolean;
  signal binary_388_inst_ack_1 : boolean;
  signal binary_394_inst_req_0 : boolean;
  signal binary_394_inst_ack_0 : boolean;
  signal binary_394_inst_req_1 : boolean;
  signal binary_394_inst_ack_1 : boolean;
  signal binary_400_inst_req_0 : boolean;
  signal binary_400_inst_ack_0 : boolean;
  signal binary_400_inst_req_1 : boolean;
  signal binary_400_inst_ack_1 : boolean;
  signal binary_405_inst_req_0 : boolean;
  signal binary_405_inst_ack_0 : boolean;
  signal binary_405_inst_req_1 : boolean;
  signal binary_405_inst_ack_1 : boolean;
  signal binary_410_inst_req_0 : boolean;
  signal binary_410_inst_ack_0 : boolean;
  signal binary_410_inst_req_1 : boolean;
  signal binary_410_inst_ack_1 : boolean;
  signal binary_416_inst_req_0 : boolean;
  signal binary_416_inst_ack_0 : boolean;
  signal binary_416_inst_req_1 : boolean;
  signal binary_416_inst_ack_1 : boolean;
  signal simple_obj_ref_418_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_418_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_418_store_0_req_0 : boolean;
  signal simple_obj_ref_418_store_0_ack_0 : boolean;
  signal simple_obj_ref_418_store_0_req_1 : boolean;
  signal simple_obj_ref_418_store_0_ack_1 : boolean;
  signal simple_obj_ref_421_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_421_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_421_store_0_req_0 : boolean;
  signal simple_obj_ref_421_store_0_ack_0 : boolean;
  signal simple_obj_ref_421_store_0_req_1 : boolean;
  signal simple_obj_ref_421_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  ret_val_x_x <= ret_val_x_x_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  a5reg_CP_0: Block -- control-path 
    signal cp_elements: BooleanArray(376 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(376);
    cp_elements(2) <= cp_elements(0);
    cp_elements(3) <= cp_elements(2);
    simple_obj_ref_12_load_0_req_0 <= cp_elements(3);
    cp_elements(4) <= simple_obj_ref_12_load_0_ack_0;
    cp_elements(5) <= cp_elements(4);
    simple_obj_ref_12_load_0_req_1 <= cp_elements(5);
    cp_elements(6) <= simple_obj_ref_12_load_0_ack_1;
    simple_obj_ref_12_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= simple_obj_ref_12_gather_scatter_ack_0;
    cp_elements(8) <= cp_elements(2);
    simple_obj_ref_15_load_0_req_0 <= cp_elements(8);
    cp_elements(9) <= simple_obj_ref_15_load_0_ack_0;
    cp_elements(10) <= cp_elements(9);
    simple_obj_ref_15_load_0_req_1 <= cp_elements(10);
    cp_elements(11) <= simple_obj_ref_15_load_0_ack_1;
    simple_obj_ref_15_gather_scatter_req_0 <= cp_elements(11);
    cp_elements(12) <= simple_obj_ref_15_gather_scatter_ack_0;
    cp_elements(13) <= cp_elements(2);
    simple_obj_ref_18_load_0_req_0 <= cp_elements(13);
    cp_elements(14) <= simple_obj_ref_18_load_0_ack_0;
    cp_elements(15) <= cp_elements(14);
    simple_obj_ref_18_load_0_req_1 <= cp_elements(15);
    cp_elements(16) <= simple_obj_ref_18_load_0_ack_1;
    simple_obj_ref_18_gather_scatter_req_0 <= cp_elements(16);
    cp_elements(17) <= simple_obj_ref_18_gather_scatter_ack_0;
    cpelement_group_18 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(20));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(18),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_24_inst_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(2);
    cp_elements(20) <= cp_elements(7);
    cp_elements(21) <= binary_24_inst_ack_0;
    binary_24_inst_req_1 <= cp_elements(21);
    cp_elements(22) <= binary_24_inst_ack_1;
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(24) & cp_elements(25));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_30_inst_req_0 <= cp_elements(23);
    cp_elements(24) <= cp_elements(2);
    cp_elements(25) <= cp_elements(12);
    cp_elements(26) <= binary_30_inst_ack_0;
    binary_30_inst_req_1 <= cp_elements(26);
    cp_elements(27) <= binary_30_inst_ack_1;
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(29) & cp_elements(30));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_36_inst_req_0 <= cp_elements(28);
    cp_elements(29) <= cp_elements(2);
    cp_elements(30) <= cp_elements(17);
    cp_elements(31) <= binary_36_inst_ack_0;
    binary_36_inst_req_1 <= cp_elements(31);
    cp_elements(32) <= binary_36_inst_ack_1;
    cpelement_group_33 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(34));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(33),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_42_inst_req_0 <= cp_elements(33);
    cp_elements(34) <= cp_elements(2);
    cp_elements(35) <= binary_42_inst_ack_0;
    binary_42_inst_req_1 <= cp_elements(35);
    cp_elements(36) <= binary_42_inst_ack_1;
    cpelement_group_37 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(38) & cp_elements(39));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(37),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_48_inst_req_0 <= cp_elements(37);
    cp_elements(38) <= cp_elements(2);
    cp_elements(39) <= cp_elements(36);
    cp_elements(40) <= binary_48_inst_ack_0;
    binary_48_inst_req_1 <= cp_elements(40);
    cp_elements(41) <= binary_48_inst_ack_1;
    cpelement_group_42 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(43));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(42),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_54_inst_req_0 <= cp_elements(42);
    cp_elements(43) <= cp_elements(2);
    cp_elements(44) <= binary_54_inst_ack_0;
    binary_54_inst_req_1 <= cp_elements(44);
    cp_elements(45) <= binary_54_inst_ack_1;
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(47) & cp_elements(48));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_60_inst_req_0 <= cp_elements(46);
    cp_elements(47) <= cp_elements(2);
    cp_elements(48) <= cp_elements(45);
    cp_elements(49) <= binary_60_inst_ack_0;
    binary_60_inst_req_1 <= cp_elements(49);
    cp_elements(50) <= binary_60_inst_ack_1;
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(52));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_66_inst_req_0 <= cp_elements(51);
    cp_elements(52) <= cp_elements(2);
    cp_elements(53) <= binary_66_inst_ack_0;
    binary_66_inst_req_1 <= cp_elements(53);
    cp_elements(54) <= binary_66_inst_ack_1;
    cpelement_group_55 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(57));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(55),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_72_inst_req_0 <= cp_elements(55);
    cp_elements(56) <= cp_elements(2);
    cp_elements(57) <= cp_elements(54);
    cp_elements(58) <= binary_72_inst_ack_0;
    binary_72_inst_req_1 <= cp_elements(58);
    cp_elements(59) <= binary_72_inst_ack_1;
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_78_inst_req_0 <= cp_elements(60);
    cp_elements(61) <= cp_elements(2);
    cp_elements(62) <= cp_elements(45);
    cp_elements(63) <= binary_78_inst_ack_0;
    binary_78_inst_req_1 <= cp_elements(63);
    cp_elements(64) <= binary_78_inst_ack_1;
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(67));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_84_inst_req_0 <= cp_elements(65);
    cp_elements(66) <= cp_elements(2);
    cp_elements(67) <= cp_elements(54);
    cp_elements(68) <= binary_84_inst_ack_0;
    binary_84_inst_req_1 <= cp_elements(68);
    cp_elements(69) <= binary_84_inst_ack_1;
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(72) & cp_elements(73));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_89_inst_req_0 <= cp_elements(70);
    cp_elements(71) <= cp_elements(2);
    cp_elements(72) <= cp_elements(69);
    cp_elements(73) <= cp_elements(64);
    cp_elements(74) <= binary_89_inst_ack_0;
    binary_89_inst_req_1 <= cp_elements(74);
    cp_elements(75) <= binary_89_inst_ack_1;
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(77) & cp_elements(78));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_95_inst_req_0 <= cp_elements(76);
    cp_elements(77) <= cp_elements(2);
    cp_elements(78) <= cp_elements(36);
    cp_elements(79) <= binary_95_inst_ack_0;
    binary_95_inst_req_1 <= cp_elements(79);
    cp_elements(80) <= binary_95_inst_ack_1;
    cpelement_group_81 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(83) & cp_elements(84));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(81),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_100_inst_req_0 <= cp_elements(81);
    cp_elements(82) <= cp_elements(2);
    cp_elements(83) <= cp_elements(80);
    cp_elements(84) <= cp_elements(59);
    cp_elements(85) <= binary_100_inst_ack_0;
    binary_100_inst_req_1 <= cp_elements(85);
    cp_elements(86) <= binary_100_inst_ack_1;
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(88) & cp_elements(89) & cp_elements(90));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_105_inst_req_0 <= cp_elements(87);
    cp_elements(88) <= cp_elements(2);
    cp_elements(89) <= cp_elements(50);
    cp_elements(90) <= cp_elements(41);
    cp_elements(91) <= binary_105_inst_ack_0;
    binary_105_inst_req_1 <= cp_elements(91);
    cp_elements(92) <= binary_105_inst_ack_1;
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(86) & cp_elements(94) & cp_elements(95));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_110_inst_req_0 <= cp_elements(93);
    cp_elements(94) <= cp_elements(2);
    cp_elements(95) <= cp_elements(92);
    cp_elements(96) <= binary_110_inst_ack_0;
    binary_110_inst_req_1 <= cp_elements(96);
    cp_elements(97) <= binary_110_inst_ack_1;
    cpelement_group_98 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(97) & cp_elements(99) & cp_elements(100));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(98),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_115_inst_req_0 <= cp_elements(98);
    cp_elements(99) <= cp_elements(2);
    cp_elements(100) <= cp_elements(75);
    cp_elements(101) <= binary_115_inst_ack_0;
    binary_115_inst_req_1 <= cp_elements(101);
    cp_elements(102) <= binary_115_inst_ack_1;
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(104) & cp_elements(105) & cp_elements(106));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_120_inst_req_0 <= cp_elements(103);
    cp_elements(104) <= cp_elements(2);
    cp_elements(105) <= cp_elements(80);
    cp_elements(106) <= cp_elements(50);
    cp_elements(107) <= binary_120_inst_ack_0;
    binary_120_inst_req_1 <= cp_elements(107);
    cp_elements(108) <= binary_120_inst_ack_1;
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(111) & cp_elements(112));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_125_inst_req_0 <= cp_elements(109);
    cp_elements(110) <= cp_elements(2);
    cp_elements(111) <= cp_elements(59);
    cp_elements(112) <= cp_elements(41);
    cp_elements(113) <= binary_125_inst_ack_0;
    binary_125_inst_req_1 <= cp_elements(113);
    cp_elements(114) <= binary_125_inst_ack_1;
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(108) & cp_elements(114) & cp_elements(116));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_130_inst_req_0 <= cp_elements(115);
    cp_elements(116) <= cp_elements(2);
    cp_elements(117) <= binary_130_inst_ack_0;
    binary_130_inst_req_1 <= cp_elements(117);
    cp_elements(118) <= binary_130_inst_ack_1;
    cpelement_group_119 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(120) & cp_elements(121));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_135_inst_req_0 <= cp_elements(119);
    cp_elements(120) <= cp_elements(2);
    cp_elements(121) <= cp_elements(75);
    cp_elements(122) <= binary_135_inst_ack_0;
    binary_135_inst_req_1 <= cp_elements(122);
    cp_elements(123) <= binary_135_inst_ack_1;
    cpelement_group_124 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(126) & cp_elements(127));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(124),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_140_inst_req_0 <= cp_elements(124);
    cp_elements(125) <= cp_elements(2);
    cp_elements(126) <= cp_elements(69);
    cp_elements(127) <= cp_elements(80);
    cp_elements(128) <= binary_140_inst_ack_0;
    binary_140_inst_req_1 <= cp_elements(128);
    cp_elements(129) <= binary_140_inst_ack_1;
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(131) & cp_elements(132) & cp_elements(133));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_145_inst_req_0 <= cp_elements(130);
    cp_elements(131) <= cp_elements(2);
    cp_elements(132) <= cp_elements(64);
    cp_elements(133) <= cp_elements(59);
    cp_elements(134) <= binary_145_inst_ack_0;
    binary_145_inst_req_1 <= cp_elements(134);
    cp_elements(135) <= binary_145_inst_ack_1;
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(135) & cp_elements(137) & cp_elements(138));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_150_inst_req_0 <= cp_elements(136);
    cp_elements(137) <= cp_elements(2);
    cp_elements(138) <= cp_elements(92);
    cp_elements(139) <= binary_150_inst_ack_0;
    binary_150_inst_req_1 <= cp_elements(139);
    cp_elements(140) <= binary_150_inst_ack_1;
    cpelement_group_141 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(129) & cp_elements(140) & cp_elements(142));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(141),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_155_inst_req_0 <= cp_elements(141);
    cp_elements(142) <= cp_elements(2);
    cp_elements(143) <= binary_155_inst_ack_0;
    binary_155_inst_req_1 <= cp_elements(143);
    cp_elements(144) <= binary_155_inst_ack_1;
    cpelement_group_145 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(146) & cp_elements(147));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(145),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_161_inst_req_0 <= cp_elements(145);
    cp_elements(146) <= cp_elements(2);
    cp_elements(147) <= cp_elements(7);
    cp_elements(148) <= binary_161_inst_ack_0;
    binary_161_inst_req_1 <= cp_elements(148);
    cp_elements(149) <= binary_161_inst_ack_1;
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(151) & cp_elements(152));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_167_inst_req_0 <= cp_elements(150);
    cp_elements(151) <= cp_elements(2);
    cp_elements(152) <= cp_elements(7);
    cp_elements(153) <= binary_167_inst_ack_0;
    binary_167_inst_req_1 <= cp_elements(153);
    cp_elements(154) <= binary_167_inst_ack_1;
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(157));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_173_inst_req_0 <= cp_elements(155);
    cp_elements(156) <= cp_elements(2);
    cp_elements(157) <= cp_elements(7);
    cp_elements(158) <= binary_173_inst_ack_0;
    binary_173_inst_req_1 <= cp_elements(158);
    cp_elements(159) <= binary_173_inst_ack_1;
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(161) & cp_elements(162));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_179_inst_req_0 <= cp_elements(160);
    cp_elements(161) <= cp_elements(2);
    cp_elements(162) <= cp_elements(7);
    cp_elements(163) <= binary_179_inst_ack_0;
    binary_179_inst_req_1 <= cp_elements(163);
    cp_elements(164) <= binary_179_inst_ack_1;
    cpelement_group_165 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(159) & cp_elements(164) & cp_elements(166));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(165),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_184_inst_req_0 <= cp_elements(165);
    cp_elements(166) <= cp_elements(2);
    cp_elements(167) <= binary_184_inst_ack_0;
    binary_184_inst_req_1 <= cp_elements(167);
    cp_elements(168) <= binary_184_inst_ack_1;
    cpelement_group_169 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(154) & cp_elements(168) & cp_elements(170));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(169),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_189_inst_req_0 <= cp_elements(169);
    cp_elements(170) <= cp_elements(2);
    cp_elements(171) <= binary_189_inst_ack_0;
    binary_189_inst_req_1 <= cp_elements(171);
    cp_elements(172) <= binary_189_inst_ack_1;
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_194_inst_req_0 <= cp_elements(173);
    cp_elements(174) <= cp_elements(2);
    cp_elements(175) <= binary_194_inst_ack_0;
    binary_194_inst_req_1 <= cp_elements(175);
    cp_elements(176) <= binary_194_inst_ack_1;
    cpelement_group_177 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(176) & cp_elements(178));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(177),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_200_inst_req_0 <= cp_elements(177);
    cp_elements(178) <= cp_elements(2);
    cp_elements(179) <= binary_200_inst_ack_0;
    binary_200_inst_req_1 <= cp_elements(179);
    cp_elements(180) <= binary_200_inst_ack_1;
    cpelement_group_181 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(182) & cp_elements(183));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(181),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_206_inst_req_0 <= cp_elements(181);
    cp_elements(182) <= cp_elements(2);
    cp_elements(183) <= cp_elements(7);
    cp_elements(184) <= binary_206_inst_ack_0;
    binary_206_inst_req_1 <= cp_elements(184);
    cp_elements(185) <= binary_206_inst_ack_1;
    cpelement_group_186 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(185) & cp_elements(187));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(186),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_212_inst_req_0 <= cp_elements(186);
    cp_elements(187) <= cp_elements(2);
    cp_elements(188) <= binary_212_inst_ack_0;
    binary_212_inst_req_1 <= cp_elements(188);
    cp_elements(189) <= binary_212_inst_ack_1;
    cpelement_group_190 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(180) & cp_elements(189) & cp_elements(191));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(190),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_217_inst_req_0 <= cp_elements(190);
    cp_elements(191) <= cp_elements(2);
    cp_elements(192) <= binary_217_inst_ack_0;
    binary_217_inst_req_1 <= cp_elements(192);
    cp_elements(193) <= binary_217_inst_ack_1;
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(195) & cp_elements(196));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_223_inst_req_0 <= cp_elements(194);
    cp_elements(195) <= cp_elements(2);
    cp_elements(196) <= cp_elements(12);
    cp_elements(197) <= binary_223_inst_ack_0;
    binary_223_inst_req_1 <= cp_elements(197);
    cp_elements(198) <= binary_223_inst_ack_1;
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(200) & cp_elements(201));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_229_inst_req_0 <= cp_elements(199);
    cp_elements(200) <= cp_elements(2);
    cp_elements(201) <= cp_elements(12);
    cp_elements(202) <= binary_229_inst_ack_0;
    binary_229_inst_req_1 <= cp_elements(202);
    cp_elements(203) <= binary_229_inst_ack_1;
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(198) & cp_elements(203) & cp_elements(205));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_234_inst_req_0 <= cp_elements(204);
    cp_elements(205) <= cp_elements(2);
    cp_elements(206) <= binary_234_inst_ack_0;
    binary_234_inst_req_1 <= cp_elements(206);
    cp_elements(207) <= binary_234_inst_ack_1;
    cpelement_group_208 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(207) & cp_elements(209));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(208),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_240_inst_req_0 <= cp_elements(208);
    cp_elements(209) <= cp_elements(2);
    cp_elements(210) <= binary_240_inst_ack_0;
    binary_240_inst_req_1 <= cp_elements(210);
    cp_elements(211) <= binary_240_inst_ack_1;
    cpelement_group_212 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(213) & cp_elements(214));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_246_inst_req_0 <= cp_elements(212);
    cp_elements(213) <= cp_elements(2);
    cp_elements(214) <= cp_elements(12);
    cp_elements(215) <= binary_246_inst_ack_0;
    binary_246_inst_req_1 <= cp_elements(215);
    cp_elements(216) <= binary_246_inst_ack_1;
    cpelement_group_217 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(216) & cp_elements(218));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(217),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_252_inst_req_0 <= cp_elements(217);
    cp_elements(218) <= cp_elements(2);
    cp_elements(219) <= binary_252_inst_ack_0;
    binary_252_inst_req_1 <= cp_elements(219);
    cp_elements(220) <= binary_252_inst_ack_1;
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(220) & cp_elements(222));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_257_inst_req_0 <= cp_elements(221);
    cp_elements(222) <= cp_elements(2);
    cp_elements(223) <= binary_257_inst_ack_0;
    binary_257_inst_req_1 <= cp_elements(223);
    cp_elements(224) <= binary_257_inst_ack_1;
    cpelement_group_225 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(226) & cp_elements(227));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(225),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_263_inst_req_0 <= cp_elements(225);
    cp_elements(226) <= cp_elements(2);
    cp_elements(227) <= cp_elements(17);
    cp_elements(228) <= binary_263_inst_ack_0;
    binary_263_inst_req_1 <= cp_elements(228);
    cp_elements(229) <= binary_263_inst_ack_1;
    cpelement_group_230 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(231) & cp_elements(232));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(230),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_269_inst_req_0 <= cp_elements(230);
    cp_elements(231) <= cp_elements(2);
    cp_elements(232) <= cp_elements(17);
    cp_elements(233) <= binary_269_inst_ack_0;
    binary_269_inst_req_1 <= cp_elements(233);
    cp_elements(234) <= binary_269_inst_ack_1;
    cpelement_group_235 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(236) & cp_elements(237));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(235),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_275_inst_req_0 <= cp_elements(235);
    cp_elements(236) <= cp_elements(2);
    cp_elements(237) <= cp_elements(17);
    cp_elements(238) <= binary_275_inst_ack_0;
    binary_275_inst_req_1 <= cp_elements(238);
    cp_elements(239) <= binary_275_inst_ack_1;
    cpelement_group_240 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(241) & cp_elements(242));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(240),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_281_inst_req_0 <= cp_elements(240);
    cp_elements(241) <= cp_elements(2);
    cp_elements(242) <= cp_elements(17);
    cp_elements(243) <= binary_281_inst_ack_0;
    binary_281_inst_req_1 <= cp_elements(243);
    cp_elements(244) <= binary_281_inst_ack_1;
    cpelement_group_245 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(239) & cp_elements(244) & cp_elements(246));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(245),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_286_inst_req_0 <= cp_elements(245);
    cp_elements(246) <= cp_elements(2);
    cp_elements(247) <= binary_286_inst_ack_0;
    binary_286_inst_req_1 <= cp_elements(247);
    cp_elements(248) <= binary_286_inst_ack_1;
    cpelement_group_249 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(234) & cp_elements(248) & cp_elements(250));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(249),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_291_inst_req_0 <= cp_elements(249);
    cp_elements(250) <= cp_elements(2);
    cp_elements(251) <= binary_291_inst_ack_0;
    binary_291_inst_req_1 <= cp_elements(251);
    cp_elements(252) <= binary_291_inst_ack_1;
    cpelement_group_253 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(229) & cp_elements(252) & cp_elements(254));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(253),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_296_inst_req_0 <= cp_elements(253);
    cp_elements(254) <= cp_elements(2);
    cp_elements(255) <= binary_296_inst_ack_0;
    binary_296_inst_req_1 <= cp_elements(255);
    cp_elements(256) <= binary_296_inst_ack_1;
    cpelement_group_257 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(256) & cp_elements(258));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(257),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_302_inst_req_0 <= cp_elements(257);
    cp_elements(258) <= cp_elements(2);
    cp_elements(259) <= binary_302_inst_ack_0;
    binary_302_inst_req_1 <= cp_elements(259);
    cp_elements(260) <= binary_302_inst_ack_1;
    cpelement_group_261 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(263));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(261),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_308_inst_req_0 <= cp_elements(261);
    cp_elements(262) <= cp_elements(2);
    cp_elements(263) <= cp_elements(17);
    cp_elements(264) <= binary_308_inst_ack_0;
    binary_308_inst_req_1 <= cp_elements(264);
    cp_elements(265) <= binary_308_inst_ack_1;
    cpelement_group_266 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(265) & cp_elements(267));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(266),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_314_inst_req_0 <= cp_elements(266);
    cp_elements(267) <= cp_elements(2);
    cp_elements(268) <= binary_314_inst_ack_0;
    binary_314_inst_req_1 <= cp_elements(268);
    cp_elements(269) <= binary_314_inst_ack_1;
    cpelement_group_270 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(260) & cp_elements(269) & cp_elements(271));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(270),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_319_inst_req_0 <= cp_elements(270);
    cp_elements(271) <= cp_elements(2);
    cp_elements(272) <= binary_319_inst_ack_0;
    binary_319_inst_req_1 <= cp_elements(272);
    cp_elements(273) <= binary_319_inst_ack_1;
    cpelement_group_274 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(193) & cp_elements(275) & cp_elements(276));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(274),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_324_inst_req_0 <= cp_elements(274);
    cp_elements(275) <= cp_elements(2);
    cp_elements(276) <= cp_elements(144);
    cp_elements(277) <= binary_324_inst_ack_0;
    binary_324_inst_req_1 <= cp_elements(277);
    cp_elements(278) <= binary_324_inst_ack_1;
    cpelement_group_279 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(280) & cp_elements(281));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(279),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_330_inst_req_0 <= cp_elements(279);
    cp_elements(280) <= cp_elements(2);
    cp_elements(281) <= cp_elements(144);
    cp_elements(282) <= binary_330_inst_ack_0;
    binary_330_inst_req_1 <= cp_elements(282);
    cp_elements(283) <= binary_330_inst_ack_1;
    cpelement_group_284 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(286));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(284),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_335_inst_req_0 <= cp_elements(284);
    cp_elements(285) <= cp_elements(2);
    cp_elements(286) <= cp_elements(7);
    cp_elements(287) <= binary_335_inst_ack_0;
    binary_335_inst_req_1 <= cp_elements(287);
    cp_elements(288) <= binary_335_inst_ack_1;
    cpelement_group_289 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(278) & cp_elements(288) & cp_elements(290));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(289),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_340_inst_req_0 <= cp_elements(289);
    cp_elements(290) <= cp_elements(2);
    cp_elements(291) <= binary_340_inst_ack_0;
    binary_340_inst_req_1 <= cp_elements(291);
    cp_elements(292) <= binary_340_inst_ack_1;
    cpelement_group_293 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(224) & cp_elements(294) & cp_elements(295));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(293),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_345_inst_req_0 <= cp_elements(293);
    cp_elements(294) <= cp_elements(2);
    cp_elements(295) <= cp_elements(102);
    cp_elements(296) <= binary_345_inst_ack_0;
    binary_345_inst_req_1 <= cp_elements(296);
    cp_elements(297) <= binary_345_inst_ack_1;
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_351_inst_req_0 <= cp_elements(298);
    cp_elements(299) <= cp_elements(2);
    cp_elements(300) <= cp_elements(102);
    cp_elements(301) <= binary_351_inst_ack_0;
    binary_351_inst_req_1 <= cp_elements(301);
    cp_elements(302) <= binary_351_inst_ack_1;
    cpelement_group_303 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(302) & cp_elements(304) & cp_elements(305));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(303),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_356_inst_req_0 <= cp_elements(303);
    cp_elements(304) <= cp_elements(2);
    cp_elements(305) <= cp_elements(12);
    cp_elements(306) <= binary_356_inst_ack_0;
    binary_356_inst_req_1 <= cp_elements(306);
    cp_elements(307) <= binary_356_inst_ack_1;
    cpelement_group_308 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(297) & cp_elements(307) & cp_elements(309));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_361_inst_req_0 <= cp_elements(308);
    cp_elements(309) <= cp_elements(2);
    cp_elements(310) <= binary_361_inst_ack_0;
    binary_361_inst_req_1 <= cp_elements(310);
    cp_elements(311) <= binary_361_inst_ack_1;
    cpelement_group_312 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(273) & cp_elements(313) & cp_elements(314));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(312),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_366_inst_req_0 <= cp_elements(312);
    cp_elements(313) <= cp_elements(2);
    cp_elements(314) <= cp_elements(123);
    cp_elements(315) <= binary_366_inst_ack_0;
    binary_366_inst_req_1 <= cp_elements(315);
    cp_elements(316) <= binary_366_inst_ack_1;
    cpelement_group_317 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(318) & cp_elements(319));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(317),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_372_inst_req_0 <= cp_elements(317);
    cp_elements(318) <= cp_elements(2);
    cp_elements(319) <= cp_elements(123);
    cp_elements(320) <= binary_372_inst_ack_0;
    binary_372_inst_req_1 <= cp_elements(320);
    cp_elements(321) <= binary_372_inst_ack_1;
    cpelement_group_322 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(321) & cp_elements(323) & cp_elements(324));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(322),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_377_inst_req_0 <= cp_elements(322);
    cp_elements(323) <= cp_elements(2);
    cp_elements(324) <= cp_elements(17);
    cp_elements(325) <= binary_377_inst_ack_0;
    binary_377_inst_req_1 <= cp_elements(325);
    cp_elements(326) <= binary_377_inst_ack_1;
    cpelement_group_327 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(316) & cp_elements(326) & cp_elements(328));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(327),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_382_inst_req_0 <= cp_elements(327);
    cp_elements(328) <= cp_elements(2);
    cp_elements(329) <= binary_382_inst_ack_0;
    binary_382_inst_req_1 <= cp_elements(329);
    cp_elements(330) <= binary_382_inst_ack_1;
    cpelement_group_331 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(332) & cp_elements(333));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(331),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_388_inst_req_0 <= cp_elements(331);
    cp_elements(332) <= cp_elements(2);
    cp_elements(333) <= cp_elements(292);
    cp_elements(334) <= binary_388_inst_ack_0;
    binary_388_inst_req_1 <= cp_elements(334);
    cp_elements(335) <= binary_388_inst_ack_1;
    cpelement_group_336 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(337) & cp_elements(338));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(336),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_394_inst_req_0 <= cp_elements(336);
    cp_elements(337) <= cp_elements(2);
    cp_elements(338) <= cp_elements(311);
    cp_elements(339) <= binary_394_inst_ack_0;
    binary_394_inst_req_1 <= cp_elements(339);
    cp_elements(340) <= binary_394_inst_ack_1;
    cpelement_group_341 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(342) & cp_elements(343));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(341),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_400_inst_req_0 <= cp_elements(341);
    cp_elements(342) <= cp_elements(2);
    cp_elements(343) <= cp_elements(330);
    cp_elements(344) <= binary_400_inst_ack_0;
    binary_400_inst_req_1 <= cp_elements(344);
    cp_elements(345) <= binary_400_inst_ack_1;
    cpelement_group_346 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(335) & cp_elements(340) & cp_elements(347));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(346),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_405_inst_req_0 <= cp_elements(346);
    cp_elements(347) <= cp_elements(2);
    cp_elements(348) <= binary_405_inst_ack_0;
    binary_405_inst_req_1 <= cp_elements(348);
    cp_elements(349) <= binary_405_inst_ack_1;
    cpelement_group_350 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(345) & cp_elements(349) & cp_elements(351));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(350),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_410_inst_req_0 <= cp_elements(350);
    cp_elements(351) <= cp_elements(2);
    cp_elements(352) <= binary_410_inst_ack_0;
    binary_410_inst_req_1 <= cp_elements(352);
    cp_elements(353) <= binary_410_inst_ack_1;
    cpelement_group_354 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(353) & cp_elements(355));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(354),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_416_inst_req_0 <= cp_elements(354);
    cp_elements(355) <= cp_elements(2);
    cp_elements(356) <= binary_416_inst_ack_0;
    binary_416_inst_req_1 <= cp_elements(356);
    cp_elements(357) <= binary_416_inst_ack_1;
    cp_elements(358) <= cp_elements(292);
    cpelement_group_359 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(4) & cp_elements(358) & cp_elements(360));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(359),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_418_gather_scatter_req_0 <= cp_elements(359);
    cp_elements(360) <= cp_elements(2);
    cp_elements(361) <= simple_obj_ref_418_gather_scatter_ack_0;
    simple_obj_ref_418_store_0_req_0 <= cp_elements(361);
    cp_elements(362) <= simple_obj_ref_418_store_0_ack_0;
    simple_obj_ref_418_store_0_req_1 <= cp_elements(362);
    cp_elements(363) <= simple_obj_ref_418_store_0_ack_1;
    cp_elements(364) <= cp_elements(311);
    cpelement_group_365 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(9) & cp_elements(364) & cp_elements(366));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(365),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_421_gather_scatter_req_0 <= cp_elements(365);
    cp_elements(366) <= cp_elements(2);
    cp_elements(367) <= simple_obj_ref_421_gather_scatter_ack_0;
    simple_obj_ref_421_store_0_req_0 <= cp_elements(367);
    cp_elements(368) <= simple_obj_ref_421_store_0_ack_0;
    simple_obj_ref_421_store_0_req_1 <= cp_elements(368);
    cp_elements(369) <= simple_obj_ref_421_store_0_ack_1;
    cp_elements(370) <= cp_elements(330);
    cpelement_group_371 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(370) & cp_elements(372));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_424_gather_scatter_req_0 <= cp_elements(371);
    cp_elements(372) <= cp_elements(2);
    cp_elements(373) <= simple_obj_ref_424_gather_scatter_ack_0;
    simple_obj_ref_424_store_0_req_0 <= cp_elements(373);
    cp_elements(374) <= simple_obj_ref_424_store_0_ack_0;
    simple_obj_ref_424_store_0_req_1 <= cp_elements(374);
    cp_elements(375) <= simple_obj_ref_424_store_0_ack_1;
    cpelement_group_376 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(357) & cp_elements(363) & cp_elements(369) & cp_elements(375));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(376),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal iNsTr_0_13 : std_logic_vector(31 downto 0);
    signal iNsTr_10_67 : std_logic_vector(31 downto 0);
    signal iNsTr_11_73 : std_logic_vector(31 downto 0);
    signal iNsTr_12_79 : std_logic_vector(31 downto 0);
    signal iNsTr_13_85 : std_logic_vector(31 downto 0);
    signal iNsTr_14_90 : std_logic_vector(31 downto 0);
    signal iNsTr_15_96 : std_logic_vector(31 downto 0);
    signal iNsTr_16_101 : std_logic_vector(31 downto 0);
    signal iNsTr_17_106 : std_logic_vector(31 downto 0);
    signal iNsTr_18_111 : std_logic_vector(31 downto 0);
    signal iNsTr_19_116 : std_logic_vector(31 downto 0);
    signal iNsTr_1_16 : std_logic_vector(31 downto 0);
    signal iNsTr_20_121 : std_logic_vector(31 downto 0);
    signal iNsTr_21_126 : std_logic_vector(31 downto 0);
    signal iNsTr_22_131 : std_logic_vector(31 downto 0);
    signal iNsTr_23_136 : std_logic_vector(31 downto 0);
    signal iNsTr_24_141 : std_logic_vector(31 downto 0);
    signal iNsTr_25_146 : std_logic_vector(31 downto 0);
    signal iNsTr_26_151 : std_logic_vector(31 downto 0);
    signal iNsTr_27_156 : std_logic_vector(31 downto 0);
    signal iNsTr_28_162 : std_logic_vector(31 downto 0);
    signal iNsTr_29_168 : std_logic_vector(31 downto 0);
    signal iNsTr_2_19 : std_logic_vector(31 downto 0);
    signal iNsTr_30_174 : std_logic_vector(31 downto 0);
    signal iNsTr_31_180 : std_logic_vector(31 downto 0);
    signal iNsTr_32_185 : std_logic_vector(31 downto 0);
    signal iNsTr_33_190 : std_logic_vector(31 downto 0);
    signal iNsTr_34_195 : std_logic_vector(31 downto 0);
    signal iNsTr_35_201 : std_logic_vector(31 downto 0);
    signal iNsTr_36_207 : std_logic_vector(31 downto 0);
    signal iNsTr_37_213 : std_logic_vector(31 downto 0);
    signal iNsTr_38_218 : std_logic_vector(31 downto 0);
    signal iNsTr_39_224 : std_logic_vector(31 downto 0);
    signal iNsTr_3_25 : std_logic_vector(31 downto 0);
    signal iNsTr_40_230 : std_logic_vector(31 downto 0);
    signal iNsTr_41_235 : std_logic_vector(31 downto 0);
    signal iNsTr_42_241 : std_logic_vector(31 downto 0);
    signal iNsTr_43_247 : std_logic_vector(31 downto 0);
    signal iNsTr_44_253 : std_logic_vector(31 downto 0);
    signal iNsTr_45_258 : std_logic_vector(31 downto 0);
    signal iNsTr_46_264 : std_logic_vector(31 downto 0);
    signal iNsTr_47_270 : std_logic_vector(31 downto 0);
    signal iNsTr_48_276 : std_logic_vector(31 downto 0);
    signal iNsTr_49_282 : std_logic_vector(31 downto 0);
    signal iNsTr_4_31 : std_logic_vector(31 downto 0);
    signal iNsTr_50_287 : std_logic_vector(31 downto 0);
    signal iNsTr_51_292 : std_logic_vector(31 downto 0);
    signal iNsTr_52_297 : std_logic_vector(31 downto 0);
    signal iNsTr_53_303 : std_logic_vector(31 downto 0);
    signal iNsTr_54_309 : std_logic_vector(31 downto 0);
    signal iNsTr_55_315 : std_logic_vector(31 downto 0);
    signal iNsTr_56_320 : std_logic_vector(31 downto 0);
    signal iNsTr_57_325 : std_logic_vector(31 downto 0);
    signal iNsTr_58_331 : std_logic_vector(31 downto 0);
    signal iNsTr_59_336 : std_logic_vector(31 downto 0);
    signal iNsTr_5_37 : std_logic_vector(31 downto 0);
    signal iNsTr_60_341 : std_logic_vector(31 downto 0);
    signal iNsTr_61_346 : std_logic_vector(31 downto 0);
    signal iNsTr_62_352 : std_logic_vector(31 downto 0);
    signal iNsTr_63_357 : std_logic_vector(31 downto 0);
    signal iNsTr_64_362 : std_logic_vector(31 downto 0);
    signal iNsTr_65_367 : std_logic_vector(31 downto 0);
    signal iNsTr_66_373 : std_logic_vector(31 downto 0);
    signal iNsTr_67_378 : std_logic_vector(31 downto 0);
    signal iNsTr_68_383 : std_logic_vector(31 downto 0);
    signal iNsTr_69_389 : std_logic_vector(31 downto 0);
    signal iNsTr_6_43 : std_logic_vector(31 downto 0);
    signal iNsTr_70_395 : std_logic_vector(31 downto 0);
    signal iNsTr_71_401 : std_logic_vector(31 downto 0);
    signal iNsTr_72_406 : std_logic_vector(31 downto 0);
    signal iNsTr_73_411 : std_logic_vector(31 downto 0);
    signal iNsTr_7_49 : std_logic_vector(31 downto 0);
    signal iNsTr_8_55 : std_logic_vector(31 downto 0);
    signal iNsTr_9_61 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_12_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_12_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_15_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_15_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_18_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_18_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_418_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_418_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_421_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_421_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_424_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_424_word_address_0 : std_logic_vector(0 downto 0);
    signal type_cast_160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_166_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_172_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_178_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_205_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_211_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_222_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_228_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_23_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_262_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_274_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_280_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_29_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_301_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_307_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_313_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_329_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_35_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_371_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_387_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_393_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_399_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_415_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_41_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_46_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_53_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_58_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_65_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_77_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_83_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    simple_obj_ref_12_word_address_0 <= "0";
    simple_obj_ref_15_word_address_0 <= "0";
    simple_obj_ref_18_word_address_0 <= "0";
    simple_obj_ref_418_word_address_0 <= "0";
    simple_obj_ref_421_word_address_0 <= "0";
    simple_obj_ref_424_word_address_0 <= "0";
    type_cast_160_wire_constant <= "00000000000000000000000000010010";
    type_cast_166_wire_constant <= "00000000000000000000000000010001";
    type_cast_172_wire_constant <= "00000000000000000000000000010000";
    type_cast_178_wire_constant <= "00000000000000000000000000001101";
    type_cast_199_wire_constant <= "00000000000000000000000000000001";
    type_cast_205_wire_constant <= "00000000000000000000000000000001";
    type_cast_211_wire_constant <= "00000000000001111111111111111110";
    type_cast_222_wire_constant <= "00000000000000000000000000010101";
    type_cast_228_wire_constant <= "00000000000000000000000000010100";
    type_cast_239_wire_constant <= "00000000000000000000000000000001";
    type_cast_23_wire_constant <= "00000000000000000000000000001000";
    type_cast_245_wire_constant <= "00000000000000000000000000000001";
    type_cast_251_wire_constant <= "00000000001111111111111111111110";
    type_cast_262_wire_constant <= "00000000000000000000000000010110";
    type_cast_268_wire_constant <= "00000000000000000000000000010101";
    type_cast_274_wire_constant <= "00000000000000000000000000010100";
    type_cast_280_wire_constant <= "00000000000000000000000000000111";
    type_cast_29_wire_constant <= "00000000000000000000000000001010";
    type_cast_301_wire_constant <= "00000000000000000000000000000001";
    type_cast_307_wire_constant <= "00000000000000000000000000000001";
    type_cast_313_wire_constant <= "00000000011111111111111111111110";
    type_cast_329_wire_constant <= "11111111111111111111111111111111";
    type_cast_350_wire_constant <= "11111111111111111111111111111111";
    type_cast_35_wire_constant <= "00000000000000000000000000001010";
    type_cast_371_wire_constant <= "11111111111111111111111111111111";
    type_cast_387_wire_constant <= "00000000000000000000000000010010";
    type_cast_393_wire_constant <= "00000000000000000000000000010101";
    type_cast_399_wire_constant <= "00000000000000000000000000010110";
    type_cast_415_wire_constant <= "00000000000000000000000000000001";
    type_cast_41_wire_constant <= "00000000000000000000000000000001";
    type_cast_46_wire_constant <= "00000000000000000000000000000000";
    type_cast_53_wire_constant <= "00000000000000000000000000000001";
    type_cast_58_wire_constant <= "00000000000000000000000000000000";
    type_cast_65_wire_constant <= "00000000000000000000000000000001";
    type_cast_70_wire_constant <= "00000000000000000000000000000000";
    type_cast_77_wire_constant <= "11111111111111111111111111111111";
    type_cast_83_wire_constant <= "11111111111111111111111111111111";
    type_cast_94_wire_constant <= "11111111111111111111111111111111";
    simple_obj_ref_12_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_12_gather_scatter_ack_0 <= simple_obj_ref_12_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_12_data_0;
      iNsTr_0_13 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_15_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_15_gather_scatter_ack_0 <= simple_obj_ref_15_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_15_data_0;
      iNsTr_1_16 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_18_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_18_gather_scatter_ack_0 <= simple_obj_ref_18_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_18_data_0;
      iNsTr_2_19 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_418_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_418_gather_scatter_ack_0 <= simple_obj_ref_418_gather_scatter_req_0;
      aggregated_sig <= iNsTr_60_341;
      simple_obj_ref_418_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_421_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_421_gather_scatter_ack_0 <= simple_obj_ref_421_gather_scatter_req_0;
      aggregated_sig <= iNsTr_64_362;
      simple_obj_ref_421_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_424_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_424_gather_scatter_ack_0 <= simple_obj_ref_424_gather_scatter_req_0;
      aggregated_sig <= iNsTr_68_383;
      simple_obj_ref_424_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    -- shared split operator group (0) : binary_100_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_15_96 & iNsTr_11_73;
      iNsTr_16_101 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_100_inst_req_0,
          ackL => binary_100_inst_ack_0,
          reqR => binary_100_inst_req_1,
          ackR => binary_100_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_105_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_61 & iNsTr_7_49;
      iNsTr_17_106 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_105_inst_req_0,
          ackL => binary_105_inst_ack_0,
          reqR => binary_105_inst_req_1,
          ackR => binary_105_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_110_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_16_101 & iNsTr_17_106;
      iNsTr_18_111 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_110_inst_req_0,
          ackL => binary_110_inst_ack_0,
          reqR => binary_110_inst_req_1,
          ackR => binary_110_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_115_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_18_111 & iNsTr_14_90;
      iNsTr_19_116 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_115_inst_req_0,
          ackL => binary_115_inst_ack_0,
          reqR => binary_115_inst_req_1,
          ackR => binary_115_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_120_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_15_96 & iNsTr_9_61;
      iNsTr_20_121 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_120_inst_req_0,
          ackL => binary_120_inst_ack_0,
          reqR => binary_120_inst_req_1,
          ackR => binary_120_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_125_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_11_73 & iNsTr_7_49;
      iNsTr_21_126 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_125_inst_req_0,
          ackL => binary_125_inst_ack_0,
          reqR => binary_125_inst_req_1,
          ackR => binary_125_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_130_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_21_126 & iNsTr_20_121;
      iNsTr_22_131 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_130_inst_req_0,
          ackL => binary_130_inst_ack_0,
          reqR => binary_130_inst_req_1,
          ackR => binary_130_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_135_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_22_131 & iNsTr_14_90;
      iNsTr_23_136 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_135_inst_req_0,
          ackL => binary_135_inst_ack_0,
          reqR => binary_135_inst_req_1,
          ackR => binary_135_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_140_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_13_85 & iNsTr_15_96;
      iNsTr_24_141 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_140_inst_req_0,
          ackL => binary_140_inst_ack_0,
          reqR => binary_140_inst_req_1,
          ackR => binary_140_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_145_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_79 & iNsTr_11_73;
      iNsTr_25_146 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_145_inst_req_0,
          ackL => binary_145_inst_ack_0,
          reqR => binary_145_inst_req_1,
          ackR => binary_145_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_150_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_25_146 & iNsTr_17_106;
      iNsTr_26_151 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_150_inst_req_0,
          ackL => binary_150_inst_ack_0,
          reqR => binary_150_inst_req_1,
          ackR => binary_150_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_155_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_26_151 & iNsTr_24_141;
      iNsTr_27_156 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_155_inst_req_0,
          ackL => binary_155_inst_ack_0,
          reqR => binary_155_inst_req_1,
          ackR => binary_155_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_161_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13;
      iNsTr_28_162 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_161_inst_req_0,
          ackL => binary_161_inst_ack_0,
          reqR => binary_161_inst_req_1,
          ackR => binary_161_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_167_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13;
      iNsTr_29_168 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_167_inst_req_0,
          ackL => binary_167_inst_ack_0,
          reqR => binary_167_inst_req_1,
          ackR => binary_167_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_173_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13;
      iNsTr_30_174 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_173_inst_req_0,
          ackL => binary_173_inst_ack_0,
          reqR => binary_173_inst_req_1,
          ackR => binary_173_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_179_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13;
      iNsTr_31_180 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_179_inst_req_0,
          ackL => binary_179_inst_ack_0,
          reqR => binary_179_inst_req_1,
          ackR => binary_179_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_184_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_31_180 & iNsTr_30_174;
      iNsTr_32_185 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_184_inst_req_0,
          ackL => binary_184_inst_ack_0,
          reqR => binary_184_inst_req_1,
          ackR => binary_184_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_189_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_32_185 & iNsTr_29_168;
      iNsTr_33_190 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_189_inst_req_0,
          ackL => binary_189_inst_ack_0,
          reqR => binary_189_inst_req_1,
          ackR => binary_189_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_194_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_33_190 & iNsTr_28_162;
      iNsTr_34_195 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_194_inst_req_0,
          ackL => binary_194_inst_ack_0,
          reqR => binary_194_inst_req_1,
          ackR => binary_194_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_200_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_34_195;
      iNsTr_35_201 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_200_inst_req_0,
          ackL => binary_200_inst_ack_0,
          reqR => binary_200_inst_req_1,
          ackR => binary_200_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_206_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13;
      iNsTr_36_207 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_206_inst_req_0,
          ackL => binary_206_inst_ack_0,
          reqR => binary_206_inst_req_1,
          ackR => binary_206_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_212_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_36_207;
      iNsTr_37_213 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000001111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_212_inst_req_0,
          ackL => binary_212_inst_ack_0,
          reqR => binary_212_inst_req_1,
          ackR => binary_212_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_217_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_35_201 & iNsTr_37_213;
      iNsTr_38_218 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_217_inst_req_0,
          ackL => binary_217_inst_ack_0,
          reqR => binary_217_inst_req_1,
          ackR => binary_217_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_223_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_1_16;
      iNsTr_39_224 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_223_inst_req_0,
          ackL => binary_223_inst_ack_0,
          reqR => binary_223_inst_req_1,
          ackR => binary_223_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_229_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_1_16;
      iNsTr_40_230 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_229_inst_req_0,
          ackL => binary_229_inst_ack_0,
          reqR => binary_229_inst_req_1,
          ackR => binary_229_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_234_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_39_224 & iNsTr_40_230;
      iNsTr_41_235 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_234_inst_req_0,
          ackL => binary_234_inst_ack_0,
          reqR => binary_234_inst_req_1,
          ackR => binary_234_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_240_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_41_235;
      iNsTr_42_241 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_240_inst_req_0,
          ackL => binary_240_inst_ack_0,
          reqR => binary_240_inst_req_1,
          ackR => binary_240_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_246_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_1_16;
      iNsTr_43_247 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_246_inst_req_0,
          ackL => binary_246_inst_ack_0,
          reqR => binary_246_inst_req_1,
          ackR => binary_246_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_24_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13;
      iNsTr_3_25 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_24_inst_req_0,
          ackL => binary_24_inst_ack_0,
          reqR => binary_24_inst_req_1,
          ackR => binary_24_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_252_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_43_247;
      iNsTr_44_253 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000001111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_252_inst_req_0,
          ackL => binary_252_inst_ack_0,
          reqR => binary_252_inst_req_1,
          ackR => binary_252_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_257_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_42_241 & iNsTr_44_253;
      iNsTr_45_258 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_257_inst_req_0,
          ackL => binary_257_inst_ack_0,
          reqR => binary_257_inst_req_1,
          ackR => binary_257_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_263_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19;
      iNsTr_46_264 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_263_inst_req_0,
          ackL => binary_263_inst_ack_0,
          reqR => binary_263_inst_req_1,
          ackR => binary_263_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_269_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19;
      iNsTr_47_270 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_269_inst_req_0,
          ackL => binary_269_inst_ack_0,
          reqR => binary_269_inst_req_1,
          ackR => binary_269_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_275_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19;
      iNsTr_48_276 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_275_inst_req_0,
          ackL => binary_275_inst_ack_0,
          reqR => binary_275_inst_req_1,
          ackR => binary_275_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_281_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19;
      iNsTr_49_282 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_281_inst_req_0,
          ackL => binary_281_inst_ack_0,
          reqR => binary_281_inst_req_1,
          ackR => binary_281_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_286_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_49_282 & iNsTr_48_276;
      iNsTr_50_287 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_286_inst_req_0,
          ackL => binary_286_inst_ack_0,
          reqR => binary_286_inst_req_1,
          ackR => binary_286_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_291_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_50_287 & iNsTr_47_270;
      iNsTr_51_292 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_291_inst_req_0,
          ackL => binary_291_inst_ack_0,
          reqR => binary_291_inst_req_1,
          ackR => binary_291_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_296_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_51_292 & iNsTr_46_264;
      iNsTr_52_297 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_296_inst_req_0,
          ackL => binary_296_inst_ack_0,
          reqR => binary_296_inst_req_1,
          ackR => binary_296_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_302_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_52_297;
      iNsTr_53_303 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_302_inst_req_0,
          ackL => binary_302_inst_ack_0,
          reqR => binary_302_inst_req_1,
          ackR => binary_302_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_308_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19;
      iNsTr_54_309 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_308_inst_req_0,
          ackL => binary_308_inst_ack_0,
          reqR => binary_308_inst_req_1,
          ackR => binary_308_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_30_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_1_16;
      iNsTr_4_31 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_30_inst_req_0,
          ackL => binary_30_inst_ack_0,
          reqR => binary_30_inst_req_1,
          ackR => binary_30_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_314_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_54_309;
      iNsTr_55_315 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_314_inst_req_0,
          ackL => binary_314_inst_ack_0,
          reqR => binary_314_inst_req_1,
          ackR => binary_314_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_319_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_53_303 & iNsTr_55_315;
      iNsTr_56_320 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_319_inst_req_0,
          ackL => binary_319_inst_ack_0,
          reqR => binary_319_inst_req_1,
          ackR => binary_319_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_324_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_27_156 & iNsTr_38_218;
      iNsTr_57_325 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_324_inst_req_0,
          ackL => binary_324_inst_ack_0,
          reqR => binary_324_inst_req_1,
          ackR => binary_324_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_330_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_27_156;
      iNsTr_58_331 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_330_inst_req_0,
          ackL => binary_330_inst_ack_0,
          reqR => binary_330_inst_req_1,
          ackR => binary_330_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_335_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_0_13 & iNsTr_58_331;
      iNsTr_59_336 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_335_inst_req_0,
          ackL => binary_335_inst_ack_0,
          reqR => binary_335_inst_req_1,
          ackR => binary_335_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_340_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_57_325 & iNsTr_59_336;
      iNsTr_60_341 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_340_inst_req_0,
          ackL => binary_340_inst_ack_0,
          reqR => binary_340_inst_req_1,
          ackR => binary_340_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_345_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_19_116 & iNsTr_45_258;
      iNsTr_61_346 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_345_inst_req_0,
          ackL => binary_345_inst_ack_0,
          reqR => binary_345_inst_req_1,
          ackR => binary_345_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_351_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_19_116;
      iNsTr_62_352 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_351_inst_req_0,
          ackL => binary_351_inst_ack_0,
          reqR => binary_351_inst_req_1,
          ackR => binary_351_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_356_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_1_16 & iNsTr_62_352;
      iNsTr_63_357 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_356_inst_req_0,
          ackL => binary_356_inst_ack_0,
          reqR => binary_356_inst_req_1,
          ackR => binary_356_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_361_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_61_346 & iNsTr_63_357;
      iNsTr_64_362 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_361_inst_req_0,
          ackL => binary_361_inst_ack_0,
          reqR => binary_361_inst_req_1,
          ackR => binary_361_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_366_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_56_320 & iNsTr_23_136;
      iNsTr_65_367 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_366_inst_req_0,
          ackL => binary_366_inst_ack_0,
          reqR => binary_366_inst_req_1,
          ackR => binary_366_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_36_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19;
      iNsTr_5_37 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_36_inst_req_0,
          ackL => binary_36_inst_ack_0,
          reqR => binary_36_inst_req_1,
          ackR => binary_36_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_372_inst 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_23_136;
      iNsTr_66_373 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_372_inst_req_0,
          ackL => binary_372_inst_ack_0,
          reqR => binary_372_inst_req_1,
          ackR => binary_372_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : binary_377_inst 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_19 & iNsTr_66_373;
      iNsTr_67_378 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_377_inst_req_0,
          ackL => binary_377_inst_ack_0,
          reqR => binary_377_inst_req_1,
          ackR => binary_377_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : binary_382_inst 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_65_367 & iNsTr_67_378;
      iNsTr_68_383 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_382_inst_req_0,
          ackL => binary_382_inst_ack_0,
          reqR => binary_382_inst_req_1,
          ackR => binary_382_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : binary_388_inst 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_60_341;
      iNsTr_69_389 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_388_inst_req_0,
          ackL => binary_388_inst_ack_0,
          reqR => binary_388_inst_req_1,
          ackR => binary_388_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : binary_394_inst 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_64_362;
      iNsTr_70_395 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_394_inst_req_0,
          ackL => binary_394_inst_ack_0,
          reqR => binary_394_inst_req_1,
          ackR => binary_394_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : binary_400_inst 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_68_383;
      iNsTr_71_401 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_400_inst_req_0,
          ackL => binary_400_inst_ack_0,
          reqR => binary_400_inst_req_1,
          ackR => binary_400_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : binary_405_inst 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_69_389 & iNsTr_70_395;
      iNsTr_72_406 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_405_inst_req_0,
          ackL => binary_405_inst_ack_0,
          reqR => binary_405_inst_req_1,
          ackR => binary_405_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : binary_410_inst 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_72_406 & iNsTr_71_401;
      iNsTr_73_411 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_410_inst_req_0,
          ackL => binary_410_inst_ack_0,
          reqR => binary_410_inst_req_1,
          ackR => binary_410_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : binary_416_inst 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_73_411;
      ret_val_x_x_buffer <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_416_inst_req_0,
          ackL => binary_416_inst_ack_0,
          reqR => binary_416_inst_req_1,
          ackR => binary_416_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : binary_42_inst 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_3_25;
      iNsTr_6_43 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_42_inst_req_0,
          ackL => binary_42_inst_ack_0,
          reqR => binary_42_inst_req_1,
          ackR => binary_42_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : binary_48_inst 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_46_wire_constant & iNsTr_6_43;
      iNsTr_7_49 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_48_inst_req_0,
          ackL => binary_48_inst_ack_0,
          reqR => binary_48_inst_req_1,
          ackR => binary_48_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : binary_54_inst 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_31;
      iNsTr_8_55 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_54_inst_req_0,
          ackL => binary_54_inst_ack_0,
          reqR => binary_54_inst_req_1,
          ackR => binary_54_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : binary_60_inst 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_58_wire_constant & iNsTr_8_55;
      iNsTr_9_61 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_60_inst_req_0,
          ackL => binary_60_inst_ack_0,
          reqR => binary_60_inst_req_1,
          ackR => binary_60_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : binary_66_inst 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_5_37;
      iNsTr_10_67 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_66_inst_req_0,
          ackL => binary_66_inst_ack_0,
          reqR => binary_66_inst_req_1,
          ackR => binary_66_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : binary_72_inst 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_70_wire_constant & iNsTr_10_67;
      iNsTr_11_73 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_72_inst_req_0,
          ackL => binary_72_inst_ack_0,
          reqR => binary_72_inst_req_1,
          ackR => binary_72_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : binary_78_inst 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_8_55;
      iNsTr_12_79 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_78_inst_req_0,
          ackL => binary_78_inst_ack_0,
          reqR => binary_78_inst_req_1,
          ackR => binary_78_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : binary_84_inst 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_67;
      iNsTr_13_85 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_84_inst_req_0,
          ackL => binary_84_inst_ack_0,
          reqR => binary_84_inst_req_1,
          ackR => binary_84_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : binary_89_inst 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_13_85 & iNsTr_12_79;
      iNsTr_14_90 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_89_inst_req_0,
          ackL => binary_89_inst_ack_0,
          reqR => binary_89_inst_req_1,
          ackR => binary_89_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : binary_95_inst 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_6_43;
      iNsTr_15_96 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_95_inst_req_0,
          ackL => binary_95_inst_ack_0,
          reqR => binary_95_inst_req_1,
          ackR => binary_95_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared load operator group (0) : simple_obj_ref_12_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_12_load_0_req_0;
      simple_obj_ref_12_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_12_load_0_req_1;
      simple_obj_ref_12_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_12_word_address_0;
      simple_obj_ref_12_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : simple_obj_ref_15_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_15_load_0_req_0;
      simple_obj_ref_15_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_15_load_0_req_1;
      simple_obj_ref_15_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_15_word_address_0;
      simple_obj_ref_15_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : simple_obj_ref_18_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_18_load_0_req_0;
      simple_obj_ref_18_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_18_load_0_req_1;
      simple_obj_ref_18_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_18_word_address_0;
      simple_obj_ref_18_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : simple_obj_ref_418_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_418_store_0_req_0;
      simple_obj_ref_418_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_418_store_0_req_1;
      simple_obj_ref_418_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_418_word_address_0;
      data_in <= simple_obj_ref_418_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : simple_obj_ref_421_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_421_store_0_req_0;
      simple_obj_ref_421_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_421_store_0_req_1;
      simple_obj_ref_421_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_421_word_address_0;
      data_in <= simple_obj_ref_421_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : simple_obj_ref_424_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_424_store_0_req_0;
      simple_obj_ref_424_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_424_store_0_req_1;
      simple_obj_ref_424_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_424_word_address_0;
      data_in <= simple_obj_ref_424_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity main_inner is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(31 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(1 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(1 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(1 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(1 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    outpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    outpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    outpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    a5reg_call_reqs : out  std_logic_vector(0 downto 0);
    a5reg_call_acks : in   std_logic_vector(0 downto 0);
    a5reg_call_tag  :  out  std_logic_vector(0 downto 0);
    a5reg_return_reqs : out  std_logic_vector(0 downto 0);
    a5reg_return_acks : in   std_logic_vector(0 downto 0);
    a5reg_return_data : in   std_logic_vector(31 downto 0);
    a5reg_return_tag :  in   std_logic_vector(0 downto 0);
    a5init_call_reqs : out  std_logic_vector(0 downto 0);
    a5init_call_acks : in   std_logic_vector(0 downto 0);
    a5init_call_tag  :  out  std_logic_vector(0 downto 0);
    a5init_return_reqs : out  std_logic_vector(0 downto 0);
    a5init_return_acks : in   std_logic_vector(0 downto 0);
    a5init_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity main_inner;
architecture Default of main_inner is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(31 downto 0);
  signal main_inner_CP_3580_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_1241_load_0_ack_0 : boolean;
  signal ptr_deref_1229_addr_0_ack_0 : boolean;
  signal call_stmt_1233_call_ack_1 : boolean;
  signal ptr_deref_1218_store_0_ack_0 : boolean;
  signal simple_obj_ref_1207_store_0_ack_1 : boolean;
  signal binary_1280_inst_req_1 : boolean;
  signal simple_obj_ref_1207_store_0_req_0 : boolean;
  signal call_stmt_1270_call_ack_1 : boolean;
  signal simple_obj_ref_1241_gather_scatter_req_0 : boolean;
  signal call_stmt_1233_call_req_1 : boolean;
  signal simple_obj_ref_1199_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1229_addr_0_req_0 : boolean;
  signal binary_1285_inst_req_0 : boolean;
  signal call_stmt_1233_call_ack_0 : boolean;
  signal simple_obj_ref_1199_gather_scatter_req_0 : boolean;
  signal ptr_deref_1229_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1241_load_0_ack_1 : boolean;
  signal simple_obj_ref_1241_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1229_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1241_load_0_req_1 : boolean;
  signal simple_obj_ref_1237_inst_req_0 : boolean;
  signal simple_obj_ref_1195_store_0_ack_0 : boolean;
  signal simple_obj_ref_1241_load_0_req_0 : boolean;
  signal binary_1285_inst_ack_1 : boolean;
  signal binary_1275_inst_ack_1 : boolean;
  signal simple_obj_ref_1235_load_0_ack_0 : boolean;
  signal simple_obj_ref_1207_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1195_store_0_ack_1 : boolean;
  signal ptr_deref_1229_root_address_inst_ack_0 : boolean;
  signal binary_1291_inst_req_0 : boolean;
  signal ptr_deref_1229_root_address_inst_req_0 : boolean;
  signal ptr_deref_1218_store_0_req_0 : boolean;
  signal binary_1280_inst_ack_0 : boolean;
  signal simple_obj_ref_1243_inst_req_0 : boolean;
  signal simple_obj_ref_1195_store_0_req_1 : boolean;
  signal call_stmt_1270_call_ack_0 : boolean;
  signal binary_1291_inst_ack_0 : boolean;
  signal simple_obj_ref_1249_inst_req_0 : boolean;
  signal simple_obj_ref_1249_inst_ack_0 : boolean;
  signal ptr_deref_1229_base_resize_req_0 : boolean;
  signal binary_1280_inst_req_0 : boolean;
  signal binary_1291_inst_ack_1 : boolean;
  signal simple_obj_ref_1207_store_0_req_1 : boolean;
  signal binary_1280_inst_ack_1 : boolean;
  signal binary_1275_inst_req_1 : boolean;
  signal simple_obj_ref_1235_load_0_req_0 : boolean;
  signal simple_obj_ref_1247_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1243_inst_ack_0 : boolean;
  signal binary_1275_inst_req_0 : boolean;
  signal ptr_deref_1229_base_resize_ack_0 : boolean;
  signal phi_stmt_1261_req_1 : boolean;
  signal simple_obj_ref_1207_gather_scatter_req_0 : boolean;
  signal call_stmt_1270_call_req_1 : boolean;
  signal simple_obj_ref_1247_load_0_ack_0 : boolean;
  signal binary_1285_inst_req_1 : boolean;
  signal simple_obj_ref_1237_inst_ack_0 : boolean;
  signal simple_obj_ref_1199_store_0_req_1 : boolean;
  signal simple_obj_ref_1247_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1247_load_0_ack_1 : boolean;
  signal simple_obj_ref_1247_load_0_req_1 : boolean;
  signal type_cast_1267_inst_req_0 : boolean;
  signal type_cast_1267_inst_ack_0 : boolean;
  signal simple_obj_ref_1203_store_0_ack_1 : boolean;
  signal simple_obj_ref_1306_inst_req_0 : boolean;
  signal simple_obj_ref_1306_inst_ack_0 : boolean;
  signal simple_obj_ref_1203_store_0_req_1 : boolean;
  signal phi_stmt_1254_req_1 : boolean;
  signal type_cast_1260_inst_ack_0 : boolean;
  signal simple_obj_ref_1203_store_0_ack_0 : boolean;
  signal simple_obj_ref_1203_store_0_req_0 : boolean;
  signal type_cast_1260_inst_req_0 : boolean;
  signal simple_obj_ref_1203_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1203_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1247_load_0_req_0 : boolean;
  signal ptr_deref_1218_store_0_ack_1 : boolean;
  signal simple_obj_ref_1199_store_0_ack_1 : boolean;
  signal call_stmt_1270_call_req_0 : boolean;
  signal simple_obj_ref_1199_store_0_req_0 : boolean;
  signal ptr_deref_1229_store_0_req_0 : boolean;
  signal ptr_deref_1229_store_0_ack_0 : boolean;
  signal ptr_deref_1218_base_resize_req_0 : boolean;
  signal ptr_deref_1218_base_resize_ack_0 : boolean;
  signal ptr_deref_1218_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_1199_store_0_ack_0 : boolean;
  signal ptr_deref_1218_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1218_addr_0_req_0 : boolean;
  signal ptr_deref_1218_addr_0_ack_0 : boolean;
  signal ptr_deref_1218_gather_scatter_req_0 : boolean;
  signal ptr_deref_1218_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1195_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1235_load_0_req_1 : boolean;
  signal simple_obj_ref_1235_load_0_ack_1 : boolean;
  signal simple_obj_ref_1195_gather_scatter_ack_0 : boolean;
  signal binary_1285_inst_ack_0 : boolean;
  signal ptr_deref_1229_store_0_req_1 : boolean;
  signal ptr_deref_1229_store_0_ack_1 : boolean;
  signal simple_obj_ref_1207_store_0_ack_0 : boolean;
  signal call_stmt_1233_call_req_0 : boolean;
  signal simple_obj_ref_1235_gather_scatter_req_0 : boolean;
  signal phi_stmt_1261_req_0 : boolean;
  signal binary_1291_inst_req_1 : boolean;
  signal phi_stmt_1254_req_0 : boolean;
  signal binary_1275_inst_ack_0 : boolean;
  signal if_stmt_1299_branch_ack_0 : boolean;
  signal if_stmt_1299_branch_ack_1 : boolean;
  signal if_stmt_1299_branch_req_0 : boolean;
  signal binary_1297_inst_ack_1 : boolean;
  signal binary_1297_inst_ack_0 : boolean;
  signal binary_1297_inst_req_1 : boolean;
  signal binary_1297_inst_req_0 : boolean;
  signal phi_stmt_1254_ack_0 : boolean;
  signal phi_stmt_1261_ack_0 : boolean;
  signal ptr_deref_1218_store_0_req_1 : boolean;
  signal simple_obj_ref_1235_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1195_store_0_req_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  ret_val_x_x <= ret_val_x_x_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  main_inner_CP_3580: Block -- control-path 
    signal cp_elements: BooleanArray(120 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(103);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(103), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(51);
    call_stmt_1233_call_req_0 <= cp_elements(1);
    cp_elements(2) <= cp_elements(118);
    call_stmt_1270_call_req_0 <= cp_elements(2);
    cp_elements(3) <= cp_elements(93);
    cp_elements(4) <= OrReduce(cp_elements(100) & cp_elements(120));
    simple_obj_ref_1306_inst_req_0 <= cp_elements(4);
    cp_elements(5) <= cp_elements(0);
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1195_gather_scatter_req_0 <= cp_elements(7);
    cp_elements(8) <= cp_elements(5);
    cp_elements(9) <= simple_obj_ref_1195_gather_scatter_ack_0;
    simple_obj_ref_1195_store_0_req_0 <= cp_elements(9);
    cp_elements(10) <= simple_obj_ref_1195_store_0_ack_0;
    simple_obj_ref_1195_store_0_req_1 <= cp_elements(10);
    cp_elements(11) <= simple_obj_ref_1195_store_0_ack_1;
    cp_elements(12) <= cp_elements(5);
    cpelement_group_13 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(14));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(13),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1199_gather_scatter_req_0 <= cp_elements(13);
    cp_elements(14) <= cp_elements(5);
    cp_elements(15) <= simple_obj_ref_1199_gather_scatter_ack_0;
    simple_obj_ref_1199_store_0_req_0 <= cp_elements(15);
    cp_elements(16) <= simple_obj_ref_1199_store_0_ack_0;
    simple_obj_ref_1199_store_0_req_1 <= cp_elements(16);
    cp_elements(17) <= simple_obj_ref_1199_store_0_ack_1;
    cp_elements(18) <= cp_elements(5);
    cpelement_group_19 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(18) & cp_elements(20));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(19),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1203_gather_scatter_req_0 <= cp_elements(19);
    cp_elements(20) <= cp_elements(5);
    cp_elements(21) <= simple_obj_ref_1203_gather_scatter_ack_0;
    simple_obj_ref_1203_store_0_req_0 <= cp_elements(21);
    cp_elements(22) <= simple_obj_ref_1203_store_0_ack_0;
    simple_obj_ref_1203_store_0_req_1 <= cp_elements(22);
    cp_elements(23) <= simple_obj_ref_1203_store_0_ack_1;
    cp_elements(24) <= cp_elements(5);
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(24) & cp_elements(26));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    simple_obj_ref_1207_gather_scatter_req_0 <= cp_elements(25);
    cp_elements(26) <= cp_elements(5);
    cp_elements(27) <= simple_obj_ref_1207_gather_scatter_ack_0;
    simple_obj_ref_1207_store_0_req_0 <= cp_elements(27);
    cp_elements(28) <= simple_obj_ref_1207_store_0_ack_0;
    simple_obj_ref_1207_store_0_req_1 <= cp_elements(28);
    cp_elements(29) <= simple_obj_ref_1207_store_0_ack_1;
    cp_elements(30) <= cp_elements(5);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(32) & cp_elements(36));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1218_gather_scatter_req_0 <= cp_elements(31);
    cp_elements(32) <= cp_elements(5);
    cp_elements(33) <= cp_elements(32);
    ptr_deref_1218_base_resize_req_0 <= cp_elements(33);
    cp_elements(34) <= ptr_deref_1218_base_resize_ack_0;
    ptr_deref_1218_root_address_inst_req_0 <= cp_elements(34);
    cp_elements(35) <= ptr_deref_1218_root_address_inst_ack_0;
    ptr_deref_1218_addr_0_req_0 <= cp_elements(35);
    cp_elements(36) <= ptr_deref_1218_addr_0_ack_0;
    cp_elements(37) <= ptr_deref_1218_gather_scatter_ack_0;
    ptr_deref_1218_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= ptr_deref_1218_store_0_ack_0;
    cp_elements(39) <= cp_elements(38);
    ptr_deref_1218_store_0_req_1 <= cp_elements(39);
    cp_elements(40) <= ptr_deref_1218_store_0_ack_1;
    cp_elements(41) <= cp_elements(5);
    cpelement_group_42 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(38) & cp_elements(41) & cp_elements(43) & cp_elements(47));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(42),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1229_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= cp_elements(5);
    cp_elements(44) <= cp_elements(43);
    ptr_deref_1229_base_resize_req_0 <= cp_elements(44);
    cp_elements(45) <= ptr_deref_1229_base_resize_ack_0;
    ptr_deref_1229_root_address_inst_req_0 <= cp_elements(45);
    cp_elements(46) <= ptr_deref_1229_root_address_inst_ack_0;
    ptr_deref_1229_addr_0_req_0 <= cp_elements(46);
    cp_elements(47) <= ptr_deref_1229_addr_0_ack_0;
    cp_elements(48) <= ptr_deref_1229_gather_scatter_ack_0;
    ptr_deref_1229_store_0_req_0 <= cp_elements(48);
    cp_elements(49) <= ptr_deref_1229_store_0_ack_0;
    ptr_deref_1229_store_0_req_1 <= cp_elements(49);
    cp_elements(50) <= ptr_deref_1229_store_0_ack_1;
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(5 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(17) & cp_elements(23) & cp_elements(29) & cp_elements(40) & cp_elements(50));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(52) <= call_stmt_1233_call_ack_0;
    call_stmt_1233_call_req_1 <= cp_elements(52);
    cp_elements(53) <= call_stmt_1233_call_ack_1;
    simple_obj_ref_1235_load_0_req_0 <= cp_elements(53);
    cp_elements(54) <= simple_obj_ref_1235_load_0_ack_0;
    simple_obj_ref_1235_load_0_req_1 <= cp_elements(54);
    cp_elements(55) <= simple_obj_ref_1235_load_0_ack_1;
    simple_obj_ref_1235_gather_scatter_req_0 <= cp_elements(55);
    cp_elements(56) <= simple_obj_ref_1235_gather_scatter_ack_0;
    simple_obj_ref_1237_inst_req_0 <= cp_elements(56);
    cp_elements(57) <= simple_obj_ref_1237_inst_ack_0;
    simple_obj_ref_1241_load_0_req_0 <= cp_elements(57);
    cp_elements(58) <= simple_obj_ref_1241_load_0_ack_0;
    simple_obj_ref_1241_load_0_req_1 <= cp_elements(58);
    cp_elements(59) <= simple_obj_ref_1241_load_0_ack_1;
    simple_obj_ref_1241_gather_scatter_req_0 <= cp_elements(59);
    cp_elements(60) <= simple_obj_ref_1241_gather_scatter_ack_0;
    simple_obj_ref_1243_inst_req_0 <= cp_elements(60);
    cp_elements(61) <= simple_obj_ref_1243_inst_ack_0;
    simple_obj_ref_1247_load_0_req_0 <= cp_elements(61);
    cp_elements(62) <= simple_obj_ref_1247_load_0_ack_0;
    simple_obj_ref_1247_load_0_req_1 <= cp_elements(62);
    cp_elements(63) <= simple_obj_ref_1247_load_0_ack_1;
    simple_obj_ref_1247_gather_scatter_req_0 <= cp_elements(63);
    cp_elements(64) <= simple_obj_ref_1247_gather_scatter_ack_0;
    simple_obj_ref_1249_inst_req_0 <= cp_elements(64);
    cp_elements(65) <= simple_obj_ref_1249_inst_ack_0;
    cp_elements(66) <= call_stmt_1270_call_ack_0;
    call_stmt_1270_call_req_1 <= cp_elements(66);
    cp_elements(67) <= call_stmt_1270_call_ack_1;
    cp_elements(68) <= cp_elements(67);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(71));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1275_inst_req_0 <= cp_elements(69);
    cp_elements(70) <= cp_elements(68);
    cp_elements(71) <= cp_elements(68);
    cp_elements(72) <= binary_1275_inst_ack_0;
    binary_1275_inst_req_1 <= cp_elements(72);
    cp_elements(73) <= binary_1275_inst_ack_1;
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(73) & cp_elements(75) & cp_elements(76));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1280_inst_req_0 <= cp_elements(74);
    cp_elements(75) <= cp_elements(68);
    cp_elements(76) <= cp_elements(68);
    cp_elements(77) <= binary_1280_inst_ack_0;
    binary_1280_inst_req_1 <= cp_elements(77);
    cp_elements(78) <= binary_1280_inst_ack_1;
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(80) & cp_elements(81));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1285_inst_req_0 <= cp_elements(79);
    cp_elements(80) <= cp_elements(68);
    cp_elements(81) <= cp_elements(68);
    cp_elements(82) <= binary_1285_inst_ack_0;
    binary_1285_inst_req_1 <= cp_elements(82);
    cp_elements(83) <= binary_1285_inst_ack_1;
    cpelement_group_84 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(85) & cp_elements(86));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(84),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1291_inst_req_0 <= cp_elements(84);
    cp_elements(85) <= cp_elements(68);
    cp_elements(86) <= cp_elements(68);
    cp_elements(87) <= binary_1291_inst_ack_0;
    binary_1291_inst_req_1 <= cp_elements(87);
    cp_elements(88) <= binary_1291_inst_ack_1;
    cpelement_group_89 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(88) & cp_elements(90));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(89),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1297_inst_req_0 <= cp_elements(89);
    cp_elements(90) <= cp_elements(68);
    cp_elements(91) <= binary_1297_inst_ack_0;
    binary_1297_inst_req_1 <= cp_elements(91);
    cp_elements(92) <= binary_1297_inst_ack_1;
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(92));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(94) <= cp_elements(3);
    cp_elements(95) <= false;
    cp_elements(96) <= cp_elements(95);
    cp_elements(97) <= cp_elements(3);
    if_stmt_1299_branch_req_0 <= cp_elements(97);
    cp_elements(98) <= cp_elements(97);
    cp_elements(99) <= cp_elements(98);
    cp_elements(100) <= if_stmt_1299_branch_ack_1;
    cp_elements(101) <= cp_elements(98);
    cp_elements(102) <= if_stmt_1299_branch_ack_0;
    cp_elements(103) <= simple_obj_ref_1306_inst_ack_0;
    cp_elements(104) <= cp_elements(102);
    cp_elements(105) <= cp_elements(104);
    type_cast_1260_inst_req_0 <= cp_elements(105);
    cp_elements(106) <= type_cast_1260_inst_ack_0;
    phi_stmt_1254_req_1 <= cp_elements(106);
    cp_elements(107) <= cp_elements(104);
    type_cast_1267_inst_req_0 <= cp_elements(107);
    cp_elements(108) <= type_cast_1267_inst_ack_0;
    phi_stmt_1261_req_1 <= cp_elements(108);
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(110) <= cp_elements(65);
    cp_elements(111) <= cp_elements(110);
    phi_stmt_1254_req_0 <= cp_elements(111);
    cp_elements(112) <= cp_elements(110);
    phi_stmt_1261_req_0 <= cp_elements(112);
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(111) & cp_elements(112));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(114) <= OrReduce(cp_elements(109) & cp_elements(113));
    cp_elements(115) <= cp_elements(114);
    cp_elements(116) <= phi_stmt_1254_ack_0;
    cp_elements(117) <= phi_stmt_1261_ack_0;
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(116) & cp_elements(117));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(119) <= false;
    cp_elements(120) <= cp_elements(119);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal Bx_xnot_1254 : std_logic_vector(31 downto 0);
    signal exitcond_1298 : std_logic_vector(0 downto 0);
    signal iNsTr_12_1242 : std_logic_vector(31 downto 0);
    signal iNsTr_15_1248 : std_logic_vector(31 downto 0);
    signal iNsTr_19_1270 : std_logic_vector(31 downto 0);
    signal iNsTr_20_1276 : std_logic_vector(31 downto 0);
    signal iNsTr_21_1281 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1216 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1227 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1236 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1292 : std_logic_vector(31 downto 0);
    signal outx_x01_1261 : std_logic_vector(31 downto 0);
    signal ptr_deref_1218_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1218_resized_base_address : std_logic_vector(1 downto 0);
    signal ptr_deref_1218_root_address : std_logic_vector(1 downto 0);
    signal ptr_deref_1218_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1218_word_address_0 : std_logic_vector(1 downto 0);
    signal ptr_deref_1218_word_offset_0 : std_logic_vector(1 downto 0);
    signal ptr_deref_1229_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1229_resized_base_address : std_logic_vector(1 downto 0);
    signal ptr_deref_1229_root_address : std_logic_vector(1 downto 0);
    signal ptr_deref_1229_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1229_word_address_0 : std_logic_vector(1 downto 0);
    signal ptr_deref_1229_word_offset_0 : std_logic_vector(1 downto 0);
    signal simple_obj_ref_1195_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1195_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1199_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1199_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1203_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1203_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1207_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1207_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1235_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1235_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1241_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1241_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1247_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1247_word_address_0 : std_logic_vector(0 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1201_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1205_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1209_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1220_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1231_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1258_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1260_wire : std_logic_vector(31 downto 0);
    signal type_cast_1265_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1267_wire : std_logic_vector(31 downto 0);
    signal type_cast_1274_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1290_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1296_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    iNsTr_4_1216 <= "00000000000000000000000000000000";
    iNsTr_6_1227 <= "00000000000000000000000000000001";
    ptr_deref_1218_word_offset_0 <= "00";
    ptr_deref_1229_word_offset_0 <= "00";
    simple_obj_ref_1195_word_address_0 <= "0";
    simple_obj_ref_1199_word_address_0 <= "0";
    simple_obj_ref_1203_word_address_0 <= "0";
    simple_obj_ref_1207_word_address_0 <= "0";
    simple_obj_ref_1235_word_address_0 <= "0";
    simple_obj_ref_1241_word_address_0 <= "0";
    simple_obj_ref_1247_word_address_0 <= "0";
    type_cast_1197_wire_constant <= "00000000000000000000000000000000";
    type_cast_1201_wire_constant <= "00000000000000000000000000000000";
    type_cast_1205_wire_constant <= "00000000000000000000000000000000";
    type_cast_1209_wire_constant <= "00000000000000000000000000000000";
    type_cast_1220_wire_constant <= "11111111111111111111111111111111";
    type_cast_1231_wire_constant <= "11111111111111111111111111111111";
    type_cast_1258_wire_constant <= "00000000000000000000000000000000";
    type_cast_1265_wire_constant <= "00000000000000000000000000000000";
    type_cast_1274_wire_constant <= "00000000000000000000000000011111";
    type_cast_1290_wire_constant <= "00000000000000000000000000000001";
    type_cast_1296_wire_constant <= "00000000000000000000000000100000";
    phi_stmt_1254: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1258_wire_constant & type_cast_1260_wire;
      req <= phi_stmt_1254_req_0 & phi_stmt_1254_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1254_ack_0,
          idata => idata,
          odata => Bx_xnot_1254,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1254
    phi_stmt_1261: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1265_wire_constant & type_cast_1267_wire;
      req <= phi_stmt_1261_req_0 & phi_stmt_1261_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1261_ack_0,
          idata => idata,
          odata => outx_x01_1261,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1261
    ptr_deref_1218_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 2, flow_through => true ) 
      port map( din => iNsTr_4_1216, dout => ptr_deref_1218_resized_base_address, req => ptr_deref_1218_base_resize_req_0, ack => ptr_deref_1218_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1229_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 2, flow_through => true ) 
      port map( din => iNsTr_6_1227, dout => ptr_deref_1229_resized_base_address, req => ptr_deref_1229_base_resize_req_0, ack => ptr_deref_1229_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1260_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnext_1292, dout => type_cast_1260_wire, req => type_cast_1260_inst_req_0, ack => type_cast_1260_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1267_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => ret_val_x_x_buffer, dout => type_cast_1267_wire, req => type_cast_1267_inst_req_0, ack => type_cast_1267_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1218_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      ptr_deref_1218_addr_0_ack_0 <= ptr_deref_1218_addr_0_req_0;
      aggregated_sig <= ptr_deref_1218_root_address;
      ptr_deref_1218_word_address_0 <= aggregated_sig(1 downto 0);
      --
    end Block;
    ptr_deref_1218_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1218_gather_scatter_ack_0 <= ptr_deref_1218_gather_scatter_req_0;
      aggregated_sig <= type_cast_1220_wire_constant;
      ptr_deref_1218_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1218_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      ptr_deref_1218_root_address_inst_ack_0 <= ptr_deref_1218_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1218_resized_base_address;
      ptr_deref_1218_root_address <= aggregated_sig(1 downto 0);
      --
    end Block;
    ptr_deref_1229_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      ptr_deref_1229_addr_0_ack_0 <= ptr_deref_1229_addr_0_req_0;
      aggregated_sig <= ptr_deref_1229_root_address;
      ptr_deref_1229_word_address_0 <= aggregated_sig(1 downto 0);
      --
    end Block;
    ptr_deref_1229_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1229_gather_scatter_ack_0 <= ptr_deref_1229_gather_scatter_req_0;
      aggregated_sig <= type_cast_1231_wire_constant;
      ptr_deref_1229_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1229_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(1 downto 0); --
    begin -- 
      ptr_deref_1229_root_address_inst_ack_0 <= ptr_deref_1229_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1229_resized_base_address;
      ptr_deref_1229_root_address <= aggregated_sig(1 downto 0);
      --
    end Block;
    simple_obj_ref_1195_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1195_gather_scatter_ack_0 <= simple_obj_ref_1195_gather_scatter_req_0;
      aggregated_sig <= type_cast_1197_wire_constant;
      simple_obj_ref_1195_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1199_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1199_gather_scatter_ack_0 <= simple_obj_ref_1199_gather_scatter_req_0;
      aggregated_sig <= type_cast_1201_wire_constant;
      simple_obj_ref_1199_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1203_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1203_gather_scatter_ack_0 <= simple_obj_ref_1203_gather_scatter_req_0;
      aggregated_sig <= type_cast_1205_wire_constant;
      simple_obj_ref_1203_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1207_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1207_gather_scatter_ack_0 <= simple_obj_ref_1207_gather_scatter_req_0;
      aggregated_sig <= type_cast_1209_wire_constant;
      simple_obj_ref_1207_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1235_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1235_gather_scatter_ack_0 <= simple_obj_ref_1235_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_1235_data_0;
      iNsTr_9_1236 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1241_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1241_gather_scatter_ack_0 <= simple_obj_ref_1241_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_1241_data_0;
      iNsTr_12_1242 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1247_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1247_gather_scatter_ack_0 <= simple_obj_ref_1247_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_1247_data_0;
      iNsTr_15_1248 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_1299_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1298;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1299_branch_req_0,
          ack0 => if_stmt_1299_branch_ack_0,
          ack1 => if_stmt_1299_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_1275_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= Bx_xnot_1254;
      iNsTr_20_1276 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000011111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1275_inst_req_0,
          ackL => binary_1275_inst_ack_0,
          reqR => binary_1275_inst_req_1,
          ackR => binary_1275_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_1280_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_19_1270 & iNsTr_20_1276;
      iNsTr_21_1281 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1280_inst_req_0,
          ackL => binary_1280_inst_ack_0,
          reqR => binary_1280_inst_req_1,
          ackR => binary_1280_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1285_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_21_1281 & outx_x01_1261;
      ret_val_x_x_buffer <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1285_inst_req_0,
          ackL => binary_1285_inst_ack_0,
          reqR => binary_1285_inst_req_1,
          ackR => binary_1285_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1291_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= Bx_xnot_1254;
      indvarx_xnext_1292 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1291_inst_req_0,
          ackL => binary_1291_inst_ack_0,
          reqR => binary_1291_inst_req_1,
          ackR => binary_1291_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_1297_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext_1292;
      exitcond_1298 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000100000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1297_inst_req_0,
          ackL => binary_1297_inst_ack_0,
          reqR => binary_1297_inst_req_1,
          ackR => binary_1297_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared load operator group (0) : simple_obj_ref_1235_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1235_load_0_req_0;
      simple_obj_ref_1235_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1235_load_0_req_1;
      simple_obj_ref_1235_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_1235_word_address_0;
      simple_obj_ref_1235_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : simple_obj_ref_1241_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1241_load_0_req_0;
      simple_obj_ref_1241_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1241_load_0_req_1;
      simple_obj_ref_1241_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_1241_word_address_0;
      simple_obj_ref_1241_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : simple_obj_ref_1247_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1247_load_0_req_0;
      simple_obj_ref_1247_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1247_load_0_req_1;
      simple_obj_ref_1247_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_1247_word_address_0;
      simple_obj_ref_1247_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2, min_clock_period => true,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : ptr_deref_1218_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1218_store_0_req_0;
      ptr_deref_1218_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1218_store_0_req_1;
      ptr_deref_1218_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1218_word_address_0;
      data_in <= ptr_deref_1218_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 2,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(1),
          mack => memory_space_3_sr_ack(1),
          maddr => memory_space_3_sr_addr(3 downto 2),
          mdata => memory_space_3_sr_data(63 downto 32),
          mtag => memory_space_3_sr_tag(1 downto 1),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(1),
          mack => memory_space_3_sc_ack(1),
          mtag => memory_space_3_sc_tag(1 downto 1),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1229_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1229_store_0_req_0;
      ptr_deref_1229_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1229_store_0_req_1;
      ptr_deref_1229_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1229_word_address_0;
      data_in <= ptr_deref_1229_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 2,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(1 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : simple_obj_ref_1195_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1195_store_0_req_0;
      simple_obj_ref_1195_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1195_store_0_req_1;
      simple_obj_ref_1195_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_1195_word_address_0;
      data_in <= simple_obj_ref_1195_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : simple_obj_ref_1199_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1199_store_0_req_0;
      simple_obj_ref_1199_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1199_store_0_req_1;
      simple_obj_ref_1199_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_1199_word_address_0;
      data_in <= simple_obj_ref_1199_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : simple_obj_ref_1203_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1203_store_0_req_0;
      simple_obj_ref_1203_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1203_store_0_req_1;
      simple_obj_ref_1203_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_1203_word_address_0;
      data_in <= simple_obj_ref_1203_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : simple_obj_ref_1207_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1207_store_0_req_0;
      simple_obj_ref_1207_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1207_store_0_req_1;
      simple_obj_ref_1207_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_1207_word_address_0;
      data_in <= simple_obj_ref_1207_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => true,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared outport operator group (0) : simple_obj_ref_1237_inst simple_obj_ref_1243_inst simple_obj_ref_1249_inst simple_obj_ref_1306_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal req, ack : BooleanArray( 3 downto 0);
      -- 
    begin -- 
      req(3) <= simple_obj_ref_1237_inst_req_0;
      req(2) <= simple_obj_ref_1243_inst_req_0;
      req(1) <= simple_obj_ref_1249_inst_req_0;
      req(0) <= simple_obj_ref_1306_inst_req_0;
      simple_obj_ref_1237_inst_ack_0 <= ack(3);
      simple_obj_ref_1243_inst_ack_0 <= ack(2);
      simple_obj_ref_1249_inst_ack_0 <= ack(1);
      simple_obj_ref_1306_inst_ack_0 <= ack(0);
      data_in <= iNsTr_9_1236 & iNsTr_12_1242 & iNsTr_15_1248 & ret_val_x_x_buffer;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 4,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => outpipe_pipe_write_req(0),
          oack => outpipe_pipe_write_ack(0),
          odata => outpipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1233_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1233_call_req_0;
      call_stmt_1233_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1233_call_req_1;
      call_stmt_1233_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => a5init_call_reqs(0),
          ackR => a5init_call_acks(0),
          tagR => a5init_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => a5init_return_acks(0), -- cross-over
          ackL => a5init_return_reqs(0), -- cross-over
          tagL => a5init_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1270_call 
    CallGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1270_call_req_0;
      call_stmt_1270_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1270_call_req_1;
      call_stmt_1270_call_ack_1 <= ackR(0);
      iNsTr_19_1270 <= data_out(31 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => a5reg_call_reqs(0),
          ackR => a5reg_call_acks(0),
          tagR => a5reg_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 32, owidth => 32, twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => a5reg_return_acks(0), -- cross-over
          ackL => a5reg_return_reqs(0), -- cross-over
          dataL => a5reg_return_data(31 downto 0),
          tagL => a5reg_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system is  -- system 
  port (-- 
    main_inner_ret_val_x_x : out  std_logic_vector(31 downto 0);
    main_inner_tag_in: in std_logic_vector(0 downto 0);
    main_inner_tag_out: out std_logic_vector(0 downto 0);
    main_inner_start_req : in std_logic;
    main_inner_start_ack : out std_logic;
    main_inner_fin_req   : in std_logic;
    main_inner_fin_ack   : out std_logic;
    clk : in std_logic;
    reset : in std_logic;
    outpipe_pipe_read_data: out std_logic_vector(31 downto 0);
    outpipe_pipe_read_req : in std_logic_vector(0 downto 0);
    outpipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(2 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(95 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(2 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(5 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(2 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(95 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(2 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(5 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(2 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(2 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(95 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(2 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(5 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module a5init
  component a5init is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(1 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      a5reg_call_reqs : out  std_logic_vector(0 downto 0);
      a5reg_call_acks : in   std_logic_vector(0 downto 0);
      a5reg_call_tag  :  out  std_logic_vector(0 downto 0);
      a5reg_return_reqs : out  std_logic_vector(0 downto 0);
      a5reg_return_acks : in   std_logic_vector(0 downto 0);
      a5reg_return_data : in   std_logic_vector(31 downto 0);
      a5reg_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module a5init
  signal a5init_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal a5init_tag_out   : std_logic_vector(0 downto 0);
  signal a5init_start_req : std_logic;
  signal a5init_start_ack : std_logic;
  signal a5init_fin_req   : std_logic;
  signal a5init_fin_ack : std_logic;
  -- caller side aggregated signals for module a5init
  signal a5init_call_reqs: std_logic_vector(0 downto 0);
  signal a5init_call_acks: std_logic_vector(0 downto 0);
  signal a5init_return_reqs: std_logic_vector(0 downto 0);
  signal a5init_return_acks: std_logic_vector(0 downto 0);
  signal a5init_call_tag: std_logic_vector(0 downto 0);
  signal a5init_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module a5reg
  component a5reg is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module a5reg
  signal a5reg_ret_val_x_x :  std_logic_vector(31 downto 0);
  signal a5reg_out_args   : std_logic_vector(31 downto 0);
  signal a5reg_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal a5reg_tag_out   : std_logic_vector(1 downto 0);
  signal a5reg_start_req : std_logic;
  signal a5reg_start_ack : std_logic;
  signal a5reg_fin_req   : std_logic;
  signal a5reg_fin_ack : std_logic;
  -- caller side aggregated signals for module a5reg
  signal a5reg_call_reqs: std_logic_vector(1 downto 0);
  signal a5reg_call_acks: std_logic_vector(1 downto 0);
  signal a5reg_return_reqs: std_logic_vector(1 downto 0);
  signal a5reg_return_acks: std_logic_vector(1 downto 0);
  signal a5reg_call_tag: std_logic_vector(1 downto 0);
  signal a5reg_return_data: std_logic_vector(63 downto 0);
  signal a5reg_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module main_inner
  component main_inner is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(1 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(1 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(1 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(1 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      outpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      outpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      outpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      a5reg_call_reqs : out  std_logic_vector(0 downto 0);
      a5reg_call_acks : in   std_logic_vector(0 downto 0);
      a5reg_call_tag  :  out  std_logic_vector(0 downto 0);
      a5reg_return_reqs : out  std_logic_vector(0 downto 0);
      a5reg_return_acks : in   std_logic_vector(0 downto 0);
      a5reg_return_data : in   std_logic_vector(31 downto 0);
      a5reg_return_tag :  in   std_logic_vector(0 downto 0);
      a5init_call_reqs : out  std_logic_vector(0 downto 0);
      a5init_call_acks : in   std_logic_vector(0 downto 0);
      a5init_call_tag  :  out  std_logic_vector(0 downto 0);
      a5init_return_reqs : out  std_logic_vector(0 downto 0);
      a5init_return_acks : in   std_logic_vector(0 downto 0);
      a5init_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- aggregate signals for write to pipe outpipe
  signal outpipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal outpipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal outpipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module a5init
  -- call arbiter for module a5init
  a5init_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => a5init_call_reqs,
      call_acks => a5init_call_acks,
      return_reqs => a5init_return_reqs,
      return_acks => a5init_return_acks,
      call_tag  => a5init_call_tag,
      return_tag  => a5init_return_tag,
      call_mtag => a5init_tag_in,
      return_mtag => a5init_tag_out,
      call_mreq => a5init_start_req,
      call_mack => a5init_start_ack,
      return_mreq => a5init_fin_req,
      return_mack => a5init_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  a5init_instance:a5init-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => a5init_start_req,
      start_ack => a5init_start_ack,
      fin_req => a5init_fin_req,
      fin_ack => a5init_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(1 downto 1),
      memory_space_0_lr_tag => memory_space_0_lr_tag(3 downto 2),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(1 downto 1),
      memory_space_1_lr_tag => memory_space_1_lr_tag(3 downto 2),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 2),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(1 downto 1),
      memory_space_2_lr_tag => memory_space_2_lr_tag(3 downto 2),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 2),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(1 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(0 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(0 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(1 downto 1),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 32),
      memory_space_0_sr_tag => memory_space_0_sr_tag(3 downto 2),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(1 downto 1),
      memory_space_1_sr_ack => memory_space_1_sr_ack(1 downto 1),
      memory_space_1_sr_addr => memory_space_1_sr_addr(1 downto 1),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 32),
      memory_space_1_sr_tag => memory_space_1_sr_tag(3 downto 2),
      memory_space_1_sc_req => memory_space_1_sc_req(1 downto 1),
      memory_space_1_sc_ack => memory_space_1_sc_ack(1 downto 1),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(1 downto 1),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 32),
      memory_space_2_sr_tag => memory_space_2_sr_tag(3 downto 2),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 2),
      a5reg_call_reqs => a5reg_call_reqs(1 downto 1),
      a5reg_call_acks => a5reg_call_acks(1 downto 1),
      a5reg_call_tag => a5reg_call_tag(1 downto 1),
      a5reg_return_reqs => a5reg_return_reqs(1 downto 1),
      a5reg_return_acks => a5reg_return_acks(1 downto 1),
      a5reg_return_data => a5reg_return_data(63 downto 32),
      a5reg_return_tag => a5reg_return_tag(1 downto 1),
      tag_in => a5init_tag_in,
      tag_out => a5init_tag_out-- 
    ); -- 
  -- module a5reg
  a5reg_out_args <= a5reg_ret_val_x_x ;
  -- call arbiter for module a5reg
  a5reg_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      num_reqs => 2,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => a5reg_call_reqs,
      call_acks => a5reg_call_acks,
      return_reqs => a5reg_return_reqs,
      return_acks => a5reg_return_acks,
      call_tag  => a5reg_call_tag,
      return_tag  => a5reg_return_tag,
      call_mtag => a5reg_tag_in,
      return_mtag => a5reg_tag_out,
      return_data =>a5reg_return_data,
      call_mreq => a5reg_start_req,
      call_mack => a5reg_start_ack,
      return_mreq => a5reg_fin_req,
      return_mack => a5reg_fin_ack,
      return_mdata => a5reg_out_args,
      clk => clk, 
      reset => reset --
    ); --
  a5reg_instance:a5reg-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => a5reg_ret_val_x_x,
      start_req => a5reg_start_req,
      start_ack => a5reg_start_ack,
      fin_req => a5reg_fin_req,
      fin_ack => a5reg_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(2 downto 2),
      memory_space_0_lr_tag => memory_space_0_lr_tag(5 downto 4),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(95 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 4),
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(2 downto 2),
      memory_space_1_lr_tag => memory_space_1_lr_tag(5 downto 4),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 4),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(2 downto 2),
      memory_space_2_lr_tag => memory_space_2_lr_tag(5 downto 4),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(95 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 4),
      memory_space_0_sr_req => memory_space_0_sr_req(2 downto 2),
      memory_space_0_sr_ack => memory_space_0_sr_ack(2 downto 2),
      memory_space_0_sr_addr => memory_space_0_sr_addr(2 downto 2),
      memory_space_0_sr_data => memory_space_0_sr_data(95 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(5 downto 4),
      memory_space_0_sc_req => memory_space_0_sc_req(2 downto 2),
      memory_space_0_sc_ack => memory_space_0_sc_ack(2 downto 2),
      memory_space_0_sc_tag => memory_space_0_sc_tag(5 downto 4),
      memory_space_1_sr_req => memory_space_1_sr_req(2 downto 2),
      memory_space_1_sr_ack => memory_space_1_sr_ack(2 downto 2),
      memory_space_1_sr_addr => memory_space_1_sr_addr(2 downto 2),
      memory_space_1_sr_data => memory_space_1_sr_data(95 downto 64),
      memory_space_1_sr_tag => memory_space_1_sr_tag(5 downto 4),
      memory_space_1_sc_req => memory_space_1_sc_req(2 downto 2),
      memory_space_1_sc_ack => memory_space_1_sc_ack(2 downto 2),
      memory_space_1_sc_tag => memory_space_1_sc_tag(5 downto 4),
      memory_space_2_sr_req => memory_space_2_sr_req(2 downto 2),
      memory_space_2_sr_ack => memory_space_2_sr_ack(2 downto 2),
      memory_space_2_sr_addr => memory_space_2_sr_addr(2 downto 2),
      memory_space_2_sr_data => memory_space_2_sr_data(95 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(5 downto 4),
      memory_space_2_sc_req => memory_space_2_sc_req(2 downto 2),
      memory_space_2_sc_ack => memory_space_2_sc_ack(2 downto 2),
      memory_space_2_sc_tag => memory_space_2_sc_tag(5 downto 4),
      tag_in => a5reg_tag_in,
      tag_out => a5reg_tag_out-- 
    ); -- 
  -- module main_inner
  main_inner_instance:main_inner-- 
    generic map(tag_length => 1)
    port map(-- 
      ret_val_x_x => main_inner_ret_val_x_x,
      start_req => main_inner_start_req,
      start_ack => main_inner_start_ack,
      fin_req => main_inner_fin_req,
      fin_ack => main_inner_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(1 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(0 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(1 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(1 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(0 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(1 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(0 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(1 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(1 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(3 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(1 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(31 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(0 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      outpipe_pipe_write_req => outpipe_pipe_write_req(0 downto 0),
      outpipe_pipe_write_ack => outpipe_pipe_write_ack(0 downto 0),
      outpipe_pipe_write_data => outpipe_pipe_write_data(31 downto 0),
      a5reg_call_reqs => a5reg_call_reqs(0 downto 0),
      a5reg_call_acks => a5reg_call_acks(0 downto 0),
      a5reg_call_tag => a5reg_call_tag(0 downto 0),
      a5reg_return_reqs => a5reg_return_reqs(0 downto 0),
      a5reg_return_acks => a5reg_return_acks(0 downto 0),
      a5reg_return_data => a5reg_return_data(31 downto 0),
      a5reg_return_tag => a5reg_return_tag(0 downto 0),
      a5init_call_reqs => a5init_call_reqs(0 downto 0),
      a5init_call_acks => a5init_call_acks(0 downto 0),
      a5init_call_tag => a5init_call_tag(0 downto 0),
      a5init_return_reqs => a5init_return_reqs(0 downto 0),
      a5init_return_acks => a5init_return_acks(0 downto 0),
      a5init_return_tag => a5init_return_tag(0 downto 0),
      tag_in => main_inner_tag_in,
      tag_out => main_inner_tag_out-- 
    ); -- 
  outpipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => outpipe_pipe_read_req,
      read_ack => outpipe_pipe_read_ack,
      read_data => outpipe_pipe_read_data,
      write_req => outpipe_pipe_write_req,
      write_ack => outpipe_pipe_write_ack,
      write_data => outpipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  RegisterBank_memory_space_0: register_bank -- 
    generic map(-- 
      num_loads => 3,
      num_stores => 3,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_1: register_bank -- 
    generic map(-- 
      num_loads => 3,
      num_stores => 3,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_2: register_bank -- 
    generic map(-- 
      num_loads => 3,
      num_stores => 3,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_3: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 2,
      addr_width => 2,
      data_width => 32,
      tag_width => 1,
      num_registers => 2) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_4: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
