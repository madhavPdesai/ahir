-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant foo_base_address : std_logic_vector(3 downto 0) := "0000";
  constant free_queue_base_address : std_logic_vector(2 downto 0) := "000";
  constant free_queue_ram_base_address : std_logic_vector(10 downto 0) := "00000000000";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  constant xx_xstr10_base_address : std_logic_vector(4 downto 0) := "00000";
  constant xx_xstr11_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr12_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr13_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr14_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr15_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr1_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr2_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr3_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr4_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr5_base_address : std_logic_vector(4 downto 0) := "00000";
  constant xx_xstr6_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr7_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr8_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr9_base_address : std_logic_vector(4 downto 0) := "00000";
  constant xx_xstr_base_address : std_logic_vector(4 downto 0) := "00000";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_foo is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_foo;
architecture Default of default_initializer_foo is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_foo_CP_0_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_92_index_0_resize_req_0 : boolean;
  signal array_obj_ref_92_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_92_index_0_rename_req_0 : boolean;
  signal binary_89_inst_req_0 : boolean;
  signal binary_89_inst_ack_0 : boolean;
  signal binary_89_inst_req_1 : boolean;
  signal binary_89_inst_ack_1 : boolean;
  signal array_obj_ref_92_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_92_offset_inst_req_0 : boolean;
  signal array_obj_ref_92_offset_inst_ack_0 : boolean;
  signal array_obj_ref_92_root_address_inst_req_0 : boolean;
  signal array_obj_ref_92_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_92_addr_0_req_0 : boolean;
  signal array_obj_ref_92_addr_0_ack_0 : boolean;
  signal array_obj_ref_92_gather_scatter_req_0 : boolean;
  signal array_obj_ref_92_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_92_store_0_req_0 : boolean;
  signal array_obj_ref_92_store_0_ack_0 : boolean;
  signal array_obj_ref_92_store_0_req_1 : boolean;
  signal array_obj_ref_92_store_0_ack_1 : boolean;
  signal binary_98_inst_req_0 : boolean;
  signal binary_98_inst_ack_0 : boolean;
  signal binary_98_inst_req_1 : boolean;
  signal binary_98_inst_ack_1 : boolean;
  signal if_stmt_95_branch_req_0 : boolean;
  signal if_stmt_95_branch_ack_1 : boolean;
  signal if_stmt_95_branch_ack_0 : boolean;
  signal phi_stmt_79_req_0 : boolean;
  signal phi_stmt_79_req_1 : boolean;
  signal phi_stmt_79_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_foo_CP_0: Block -- control-path 
    signal cp_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(30) & cp_elements(26));
    binary_89_inst_req_0 <= cp_elements(1);
    cp_elements(2) <= OrReduce(cp_elements(23) & cp_elements(15));
    cp_elements(3) <= binary_89_inst_ack_0;
    binary_89_inst_req_1 <= cp_elements(3);
    cp_elements(4) <= binary_89_inst_ack_1;
    array_obj_ref_92_index_0_resize_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_92_index_0_resize_ack_0;
    array_obj_ref_92_index_0_rename_req_0 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_92_index_0_rename_ack_0;
    array_obj_ref_92_offset_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_92_offset_inst_ack_0;
    array_obj_ref_92_root_address_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_92_root_address_inst_ack_0;
    array_obj_ref_92_addr_0_req_0 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_92_addr_0_ack_0;
    array_obj_ref_92_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_92_gather_scatter_ack_0;
    array_obj_ref_92_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_92_store_0_ack_0;
    array_obj_ref_92_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_92_store_0_ack_1;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= false;
    cp_elements(15) <= cp_elements(14);
    cp_elements(16) <= cp_elements(12);
    binary_98_inst_req_0 <= cp_elements(16);
    cp_elements(17) <= binary_98_inst_ack_0;
    binary_98_inst_req_1 <= cp_elements(17);
    cp_elements(18) <= binary_98_inst_ack_1;
    if_stmt_95_branch_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(18);
    cp_elements(20) <= cp_elements(19);
    cp_elements(21) <= if_stmt_95_branch_ack_1;
    phi_stmt_79_req_1 <= cp_elements(21);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= if_stmt_95_branch_ack_0;
    cp_elements(24) <= cp_elements(0);
    cp_elements(25) <= false;
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(0);
    phi_stmt_79_req_0 <= cp_elements(27);
    cp_elements(28) <= OrReduce(cp_elements(21) & cp_elements(27));
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= phi_stmt_79_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_0_79 : std_logic_vector(3 downto 0);
    signal array_obj_ref_92_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_92_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_92_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_92_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_92_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_92_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_92_word_offset_0 : std_logic_vector(3 downto 0);
    signal binary_98_wire : std_logic_vector(0 downto 0);
    signal expr_88_wire_constant : std_logic_vector(3 downto 0);
    signal expr_93_wire_constant : std_logic_vector(7 downto 0);
    signal expr_97_wire_constant : std_logic_vector(3 downto 0);
    signal next_I_90 : std_logic_vector(3 downto 0);
    signal simple_obj_ref_91_resized : std_logic_vector(3 downto 0);
    signal simple_obj_ref_91_scaled : std_logic_vector(3 downto 0);
    signal type_cast_83_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    array_obj_ref_92_offset_scale_factor_0 <= "0001";
    array_obj_ref_92_resized_base_address <= "0000";
    array_obj_ref_92_word_offset_0 <= "0000";
    expr_88_wire_constant <= "0001";
    expr_93_wire_constant <= "00000000";
    expr_97_wire_constant <= "1010";
    type_cast_83_wire_constant <= "0000";
    phi_stmt_79: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_83_wire_constant & next_I_90;
      req <= phi_stmt_79_req_0 & phi_stmt_79_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_79_ack_0,
          idata => idata,
          odata => I_0_79,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_79
    array_obj_ref_92_index_0_resize: RegisterBase --
      generic map(in_data_width => 4,out_data_width => 4, flow_through => true ) 
      port map( din => I_0_79, dout => simple_obj_ref_91_resized, req => array_obj_ref_92_index_0_resize_req_0, ack => array_obj_ref_92_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_92_offset_inst: RegisterBase --
      generic map(in_data_width => 4,out_data_width => 4, flow_through => true ) 
      port map( din => simple_obj_ref_91_scaled, dout => array_obj_ref_92_final_offset, req => array_obj_ref_92_offset_inst_req_0, ack => array_obj_ref_92_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_92_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(3 downto 0); --
    begin -- 
      array_obj_ref_92_addr_0_ack_0 <= array_obj_ref_92_addr_0_req_0;
      aggregated_sig <= array_obj_ref_92_root_address;
      array_obj_ref_92_word_address_0 <= aggregated_sig(3 downto 0);
      --
    end Block;
    array_obj_ref_92_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_92_gather_scatter_ack_0 <= array_obj_ref_92_gather_scatter_req_0;
      aggregated_sig <= expr_93_wire_constant;
      array_obj_ref_92_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_92_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(3 downto 0); --
    begin -- 
      array_obj_ref_92_index_0_rename_ack_0 <= array_obj_ref_92_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_91_resized;
      simple_obj_ref_91_scaled <= aggregated_sig(3 downto 0);
      --
    end Block;
    array_obj_ref_92_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(3 downto 0); --
    begin -- 
      array_obj_ref_92_root_address_inst_ack_0 <= array_obj_ref_92_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_92_final_offset;
      array_obj_ref_92_root_address <= aggregated_sig(3 downto 0);
      --
    end Block;
    if_stmt_95_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_98_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_95_branch_req_0,
          ack0 => if_stmt_95_branch_ack_0,
          ack1 => if_stmt_95_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_89_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_0_79;
      next_I_90 <= data_out(3 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0001",
          constant_width => 4,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_89_inst_req_0,
          ackL => binary_89_inst_ack_0,
          reqR => binary_89_inst_req_1,
          ackR => binary_89_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_98_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= next_I_90;
      binary_98_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1010",
          constant_width => 4,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_98_inst_req_0,
          ackL => binary_98_inst_ack_0,
          reqR => binary_98_inst_req_1,
          ackR => binary_98_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_92_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_92_store_0_req_0;
      array_obj_ref_92_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_92_store_0_req_1;
      array_obj_ref_92_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_92_word_address_0;
      data_in <= array_obj_ref_92_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(3 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_free_queue is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_free_queue;
architecture Default of default_initializer_free_queue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_free_queue_CP_134_start: Boolean;
  -- links between control-path and data-path
  signal binary_119_inst_req_0 : boolean;
  signal binary_119_inst_ack_0 : boolean;
  signal binary_119_inst_req_1 : boolean;
  signal binary_119_inst_ack_1 : boolean;
  signal array_obj_ref_122_index_0_resize_req_0 : boolean;
  signal array_obj_ref_122_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_122_index_0_rename_req_0 : boolean;
  signal array_obj_ref_122_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_122_offset_inst_req_0 : boolean;
  signal array_obj_ref_122_offset_inst_ack_0 : boolean;
  signal array_obj_ref_122_root_address_inst_req_0 : boolean;
  signal array_obj_ref_122_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_122_addr_0_req_0 : boolean;
  signal array_obj_ref_122_addr_0_ack_0 : boolean;
  signal array_obj_ref_122_gather_scatter_req_0 : boolean;
  signal array_obj_ref_122_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_122_store_0_req_0 : boolean;
  signal array_obj_ref_122_store_0_ack_0 : boolean;
  signal array_obj_ref_122_store_0_req_1 : boolean;
  signal array_obj_ref_122_store_0_ack_1 : boolean;
  signal binary_128_inst_req_0 : boolean;
  signal binary_128_inst_ack_0 : boolean;
  signal binary_128_inst_req_1 : boolean;
  signal binary_128_inst_ack_1 : boolean;
  signal if_stmt_125_branch_req_0 : boolean;
  signal if_stmt_125_branch_ack_1 : boolean;
  signal if_stmt_125_branch_ack_0 : boolean;
  signal phi_stmt_109_req_0 : boolean;
  signal phi_stmt_109_req_1 : boolean;
  signal phi_stmt_109_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_free_queue_CP_134: Block -- control-path 
    signal cp_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(30) & cp_elements(26));
    binary_119_inst_req_0 <= cp_elements(1);
    cp_elements(2) <= OrReduce(cp_elements(23) & cp_elements(15));
    cp_elements(3) <= binary_119_inst_ack_0;
    binary_119_inst_req_1 <= cp_elements(3);
    cp_elements(4) <= binary_119_inst_ack_1;
    array_obj_ref_122_index_0_resize_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_122_index_0_resize_ack_0;
    array_obj_ref_122_index_0_rename_req_0 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_122_index_0_rename_ack_0;
    array_obj_ref_122_offset_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_122_offset_inst_ack_0;
    array_obj_ref_122_root_address_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_122_root_address_inst_ack_0;
    array_obj_ref_122_addr_0_req_0 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_122_addr_0_ack_0;
    array_obj_ref_122_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_122_gather_scatter_ack_0;
    array_obj_ref_122_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_122_store_0_ack_0;
    array_obj_ref_122_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_122_store_0_ack_1;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= false;
    cp_elements(15) <= cp_elements(14);
    cp_elements(16) <= cp_elements(12);
    binary_128_inst_req_0 <= cp_elements(16);
    cp_elements(17) <= binary_128_inst_ack_0;
    binary_128_inst_req_1 <= cp_elements(17);
    cp_elements(18) <= binary_128_inst_ack_1;
    if_stmt_125_branch_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(18);
    cp_elements(20) <= cp_elements(19);
    cp_elements(21) <= if_stmt_125_branch_ack_1;
    phi_stmt_109_req_1 <= cp_elements(21);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= if_stmt_125_branch_ack_0;
    cp_elements(24) <= cp_elements(0);
    cp_elements(25) <= false;
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(0);
    phi_stmt_109_req_0 <= cp_elements(27);
    cp_elements(28) <= OrReduce(cp_elements(21) & cp_elements(27));
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= phi_stmt_109_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_0_109 : std_logic_vector(2 downto 0);
    signal array_obj_ref_122_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_122_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_122_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_122_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_122_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_122_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_122_word_offset_0 : std_logic_vector(2 downto 0);
    signal binary_128_wire : std_logic_vector(0 downto 0);
    signal expr_118_wire_constant : std_logic_vector(2 downto 0);
    signal expr_123_wire_constant : std_logic_vector(7 downto 0);
    signal expr_127_wire_constant : std_logic_vector(2 downto 0);
    signal next_I_120 : std_logic_vector(2 downto 0);
    signal simple_obj_ref_121_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_121_scaled : std_logic_vector(2 downto 0);
    signal type_cast_113_wire_constant : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    array_obj_ref_122_offset_scale_factor_0 <= "001";
    array_obj_ref_122_resized_base_address <= "000";
    array_obj_ref_122_word_offset_0 <= "000";
    expr_118_wire_constant <= "001";
    expr_123_wire_constant <= "00000000";
    expr_127_wire_constant <= "100";
    type_cast_113_wire_constant <= "000";
    phi_stmt_109: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_113_wire_constant & next_I_120;
      req <= phi_stmt_109_req_0 & phi_stmt_109_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_109_ack_0,
          idata => idata,
          odata => I_0_109,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_109
    array_obj_ref_122_index_0_resize: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => I_0_109, dout => simple_obj_ref_121_resized, req => array_obj_ref_122_index_0_resize_req_0, ack => array_obj_ref_122_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_122_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_121_scaled, dout => array_obj_ref_122_final_offset, req => array_obj_ref_122_offset_inst_req_0, ack => array_obj_ref_122_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_122_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_122_addr_0_ack_0 <= array_obj_ref_122_addr_0_req_0;
      aggregated_sig <= array_obj_ref_122_root_address;
      array_obj_ref_122_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_122_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_122_gather_scatter_ack_0 <= array_obj_ref_122_gather_scatter_req_0;
      aggregated_sig <= expr_123_wire_constant;
      array_obj_ref_122_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_122_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_122_index_0_rename_ack_0 <= array_obj_ref_122_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_121_resized;
      simple_obj_ref_121_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_122_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_122_root_address_inst_ack_0 <= array_obj_ref_122_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_122_final_offset;
      array_obj_ref_122_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    if_stmt_125_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_128_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_125_branch_req_0,
          ack0 => if_stmt_125_branch_ack_0,
          ack1 => if_stmt_125_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_119_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_0_109;
      next_I_120 <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "001",
          constant_width => 3,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_119_inst_req_0,
          ackL => binary_119_inst_ack_0,
          reqR => binary_119_inst_req_1,
          ackR => binary_119_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_128_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= next_I_120;
      binary_128_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_128_inst_req_0,
          ackL => binary_128_inst_ack_0,
          reqR => binary_128_inst_req_1,
          ackR => binary_128_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_122_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_122_store_0_req_0;
      array_obj_ref_122_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_122_store_0_req_1;
      array_obj_ref_122_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_122_word_address_0;
      data_in <= array_obj_ref_122_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(2 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_free_queue_ram is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_free_queue_ram;
architecture Default of default_initializer_free_queue_ram is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_free_queue_ram_CP_268_start: Boolean;
  -- links between control-path and data-path
  signal binary_148_inst_req_0 : boolean;
  signal binary_148_inst_ack_0 : boolean;
  signal binary_148_inst_req_1 : boolean;
  signal binary_148_inst_ack_1 : boolean;
  signal array_obj_ref_151_index_0_resize_req_0 : boolean;
  signal array_obj_ref_151_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_151_index_0_rename_req_0 : boolean;
  signal array_obj_ref_151_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_151_offset_inst_req_0 : boolean;
  signal array_obj_ref_151_offset_inst_ack_0 : boolean;
  signal array_obj_ref_151_root_address_inst_req_0 : boolean;
  signal array_obj_ref_151_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_151_addr_0_req_0 : boolean;
  signal array_obj_ref_151_addr_0_ack_0 : boolean;
  signal array_obj_ref_151_gather_scatter_req_0 : boolean;
  signal array_obj_ref_151_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_151_store_0_req_0 : boolean;
  signal array_obj_ref_151_store_0_ack_0 : boolean;
  signal array_obj_ref_151_store_0_req_1 : boolean;
  signal array_obj_ref_151_store_0_ack_1 : boolean;
  signal binary_157_inst_req_0 : boolean;
  signal binary_157_inst_ack_0 : boolean;
  signal binary_157_inst_req_1 : boolean;
  signal binary_157_inst_ack_1 : boolean;
  signal if_stmt_154_branch_req_0 : boolean;
  signal if_stmt_154_branch_ack_1 : boolean;
  signal if_stmt_154_branch_ack_0 : boolean;
  signal phi_stmt_138_req_0 : boolean;
  signal phi_stmt_138_req_1 : boolean;
  signal phi_stmt_138_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_free_queue_ram_CP_268: Block -- control-path 
    signal cp_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(26) & cp_elements(30));
    binary_148_inst_req_0 <= cp_elements(1);
    cp_elements(2) <= OrReduce(cp_elements(15) & cp_elements(23));
    cp_elements(3) <= binary_148_inst_ack_0;
    binary_148_inst_req_1 <= cp_elements(3);
    cp_elements(4) <= binary_148_inst_ack_1;
    array_obj_ref_151_index_0_resize_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_151_index_0_resize_ack_0;
    array_obj_ref_151_index_0_rename_req_0 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_151_index_0_rename_ack_0;
    array_obj_ref_151_offset_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_151_offset_inst_ack_0;
    array_obj_ref_151_root_address_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_151_root_address_inst_ack_0;
    array_obj_ref_151_addr_0_req_0 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_151_addr_0_ack_0;
    array_obj_ref_151_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_151_gather_scatter_ack_0;
    array_obj_ref_151_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_151_store_0_ack_0;
    array_obj_ref_151_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_151_store_0_ack_1;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= false;
    cp_elements(15) <= cp_elements(14);
    cp_elements(16) <= cp_elements(12);
    binary_157_inst_req_0 <= cp_elements(16);
    cp_elements(17) <= binary_157_inst_ack_0;
    binary_157_inst_req_1 <= cp_elements(17);
    cp_elements(18) <= binary_157_inst_ack_1;
    if_stmt_154_branch_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(18);
    cp_elements(20) <= cp_elements(19);
    cp_elements(21) <= if_stmt_154_branch_ack_1;
    phi_stmt_138_req_1 <= cp_elements(21);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= if_stmt_154_branch_ack_0;
    cp_elements(24) <= cp_elements(0);
    cp_elements(25) <= false;
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(0);
    phi_stmt_138_req_0 <= cp_elements(27);
    cp_elements(28) <= OrReduce(cp_elements(21) & cp_elements(27));
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= phi_stmt_138_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_0_138 : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_151_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_word_offset_0 : std_logic_vector(10 downto 0);
    signal binary_157_wire : std_logic_vector(0 downto 0);
    signal expr_147_wire_constant : std_logic_vector(10 downto 0);
    signal expr_152_wire_constant : std_logic_vector(7 downto 0);
    signal expr_156_wire_constant : std_logic_vector(10 downto 0);
    signal next_I_149 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_150_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_150_scaled : std_logic_vector(10 downto 0);
    signal type_cast_142_wire_constant : std_logic_vector(10 downto 0);
    -- 
  begin -- 
    array_obj_ref_151_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_151_resized_base_address <= "00000000000";
    array_obj_ref_151_word_offset_0 <= "00000000000";
    expr_147_wire_constant <= "00000000001";
    expr_152_wire_constant <= "00000000";
    expr_156_wire_constant <= "10000000000";
    type_cast_142_wire_constant <= "00000000000";
    phi_stmt_138: Block -- phi operator 
      signal idata: std_logic_vector(21 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_142_wire_constant & next_I_149;
      req <= phi_stmt_138_req_0 & phi_stmt_138_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 11) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_138_ack_0,
          idata => idata,
          odata => I_0_138,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_138
    array_obj_ref_151_index_0_resize: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => I_0_138, dout => simple_obj_ref_150_resized, req => array_obj_ref_151_index_0_resize_req_0, ack => array_obj_ref_151_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_151_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_150_scaled, dout => array_obj_ref_151_final_offset, req => array_obj_ref_151_offset_inst_req_0, ack => array_obj_ref_151_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_151_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_151_addr_0_ack_0 <= array_obj_ref_151_addr_0_req_0;
      aggregated_sig <= array_obj_ref_151_root_address;
      array_obj_ref_151_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_151_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_151_gather_scatter_ack_0 <= array_obj_ref_151_gather_scatter_req_0;
      aggregated_sig <= expr_152_wire_constant;
      array_obj_ref_151_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_151_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_151_index_0_rename_ack_0 <= array_obj_ref_151_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_150_resized;
      simple_obj_ref_150_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_151_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_151_root_address_inst_ack_0 <= array_obj_ref_151_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_151_final_offset;
      array_obj_ref_151_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_154_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_157_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_154_branch_req_0,
          ack0 => if_stmt_154_branch_ack_0,
          ack1 => if_stmt_154_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_148_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_0_138;
      next_I_149 <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_148_inst_req_0,
          ackL => binary_148_inst_ack_0,
          reqR => binary_148_inst_req_1,
          ackR => binary_148_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_157_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= next_I_149;
      binary_157_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10000000000",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_157_inst_req_0,
          ackL => binary_157_inst_ack_0,
          reqR => binary_157_inst_req_1,
          ackR => binary_157_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_151_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_151_store_0_req_0;
      array_obj_ref_151_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_151_store_0_req_1;
      array_obj_ref_151_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_151_word_address_0;
      data_in <= array_obj_ref_151_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(10 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr;
architecture Default of default_initializer_xx_xstr is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr_CP_402_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_166_gather_scatter_req_0 : boolean;
  signal array_obj_ref_166_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_166_store_0_req_0 : boolean;
  signal array_obj_ref_166_store_0_ack_0 : boolean;
  signal array_obj_ref_166_store_0_req_1 : boolean;
  signal array_obj_ref_166_store_0_ack_1 : boolean;
  signal array_obj_ref_170_gather_scatter_req_0 : boolean;
  signal array_obj_ref_170_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_170_store_0_req_0 : boolean;
  signal array_obj_ref_170_store_0_ack_0 : boolean;
  signal array_obj_ref_170_store_0_req_1 : boolean;
  signal array_obj_ref_170_store_0_ack_1 : boolean;
  signal array_obj_ref_174_gather_scatter_req_0 : boolean;
  signal array_obj_ref_174_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_174_store_0_req_0 : boolean;
  signal array_obj_ref_174_store_0_ack_0 : boolean;
  signal array_obj_ref_174_store_0_req_1 : boolean;
  signal array_obj_ref_174_store_0_ack_1 : boolean;
  signal array_obj_ref_178_gather_scatter_req_0 : boolean;
  signal array_obj_ref_178_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_178_store_0_req_0 : boolean;
  signal array_obj_ref_178_store_0_ack_0 : boolean;
  signal array_obj_ref_178_store_0_req_1 : boolean;
  signal array_obj_ref_178_store_0_ack_1 : boolean;
  signal array_obj_ref_182_gather_scatter_req_0 : boolean;
  signal array_obj_ref_182_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_182_store_0_req_0 : boolean;
  signal array_obj_ref_182_store_0_ack_0 : boolean;
  signal array_obj_ref_182_store_0_req_1 : boolean;
  signal array_obj_ref_182_store_0_ack_1 : boolean;
  signal array_obj_ref_186_gather_scatter_req_0 : boolean;
  signal array_obj_ref_186_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_186_store_0_req_0 : boolean;
  signal array_obj_ref_186_store_0_ack_0 : boolean;
  signal array_obj_ref_186_store_0_req_1 : boolean;
  signal array_obj_ref_186_store_0_ack_1 : boolean;
  signal array_obj_ref_190_gather_scatter_req_0 : boolean;
  signal array_obj_ref_190_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_190_store_0_req_0 : boolean;
  signal array_obj_ref_190_store_0_ack_0 : boolean;
  signal array_obj_ref_190_store_0_req_1 : boolean;
  signal array_obj_ref_190_store_0_ack_1 : boolean;
  signal array_obj_ref_194_gather_scatter_req_0 : boolean;
  signal array_obj_ref_194_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_194_store_0_req_0 : boolean;
  signal array_obj_ref_194_store_0_ack_0 : boolean;
  signal array_obj_ref_194_store_0_req_1 : boolean;
  signal array_obj_ref_194_store_0_ack_1 : boolean;
  signal array_obj_ref_198_gather_scatter_req_0 : boolean;
  signal array_obj_ref_198_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_198_store_0_req_0 : boolean;
  signal array_obj_ref_198_store_0_ack_0 : boolean;
  signal array_obj_ref_198_store_0_req_1 : boolean;
  signal array_obj_ref_198_store_0_ack_1 : boolean;
  signal array_obj_ref_202_gather_scatter_req_0 : boolean;
  signal array_obj_ref_202_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_202_store_0_req_0 : boolean;
  signal array_obj_ref_202_store_0_ack_0 : boolean;
  signal array_obj_ref_202_store_0_req_1 : boolean;
  signal array_obj_ref_202_store_0_ack_1 : boolean;
  signal array_obj_ref_206_gather_scatter_req_0 : boolean;
  signal array_obj_ref_206_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_206_store_0_req_0 : boolean;
  signal array_obj_ref_206_store_0_ack_0 : boolean;
  signal array_obj_ref_206_store_0_req_1 : boolean;
  signal array_obj_ref_206_store_0_ack_1 : boolean;
  signal array_obj_ref_210_gather_scatter_req_0 : boolean;
  signal array_obj_ref_210_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_210_store_0_req_0 : boolean;
  signal array_obj_ref_210_store_0_ack_0 : boolean;
  signal array_obj_ref_210_store_0_req_1 : boolean;
  signal array_obj_ref_210_store_0_ack_1 : boolean;
  signal array_obj_ref_214_gather_scatter_req_0 : boolean;
  signal array_obj_ref_214_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_214_store_0_req_0 : boolean;
  signal array_obj_ref_214_store_0_ack_0 : boolean;
  signal array_obj_ref_214_store_0_req_1 : boolean;
  signal array_obj_ref_214_store_0_ack_1 : boolean;
  signal array_obj_ref_218_gather_scatter_req_0 : boolean;
  signal array_obj_ref_218_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_218_store_0_req_0 : boolean;
  signal array_obj_ref_218_store_0_ack_0 : boolean;
  signal array_obj_ref_218_store_0_req_1 : boolean;
  signal array_obj_ref_218_store_0_ack_1 : boolean;
  signal array_obj_ref_222_gather_scatter_req_0 : boolean;
  signal array_obj_ref_222_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_222_store_0_req_0 : boolean;
  signal array_obj_ref_222_store_0_ack_0 : boolean;
  signal array_obj_ref_222_store_0_req_1 : boolean;
  signal array_obj_ref_222_store_0_ack_1 : boolean;
  signal array_obj_ref_226_gather_scatter_req_0 : boolean;
  signal array_obj_ref_226_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_226_store_0_req_0 : boolean;
  signal array_obj_ref_226_store_0_ack_0 : boolean;
  signal array_obj_ref_226_store_0_req_1 : boolean;
  signal array_obj_ref_226_store_0_ack_1 : boolean;
  signal array_obj_ref_230_gather_scatter_req_0 : boolean;
  signal array_obj_ref_230_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_230_store_0_req_0 : boolean;
  signal array_obj_ref_230_store_0_ack_0 : boolean;
  signal array_obj_ref_230_store_0_req_1 : boolean;
  signal array_obj_ref_230_store_0_ack_1 : boolean;
  signal array_obj_ref_234_gather_scatter_req_0 : boolean;
  signal array_obj_ref_234_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_234_store_0_req_0 : boolean;
  signal array_obj_ref_234_store_0_ack_0 : boolean;
  signal array_obj_ref_234_store_0_req_1 : boolean;
  signal array_obj_ref_234_store_0_ack_1 : boolean;
  signal array_obj_ref_238_gather_scatter_req_0 : boolean;
  signal array_obj_ref_238_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_238_store_0_req_0 : boolean;
  signal array_obj_ref_238_store_0_ack_0 : boolean;
  signal array_obj_ref_238_store_0_req_1 : boolean;
  signal array_obj_ref_238_store_0_ack_1 : boolean;
  signal array_obj_ref_242_gather_scatter_req_0 : boolean;
  signal array_obj_ref_242_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_242_store_0_req_0 : boolean;
  signal array_obj_ref_242_store_0_ack_0 : boolean;
  signal array_obj_ref_242_store_0_req_1 : boolean;
  signal array_obj_ref_242_store_0_ack_1 : boolean;
  signal array_obj_ref_246_gather_scatter_req_0 : boolean;
  signal array_obj_ref_246_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_246_store_0_req_0 : boolean;
  signal array_obj_ref_246_store_0_ack_0 : boolean;
  signal array_obj_ref_246_store_0_req_1 : boolean;
  signal array_obj_ref_246_store_0_ack_1 : boolean;
  signal array_obj_ref_250_gather_scatter_req_0 : boolean;
  signal array_obj_ref_250_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_250_store_0_req_0 : boolean;
  signal array_obj_ref_250_store_0_ack_0 : boolean;
  signal array_obj_ref_250_store_0_req_1 : boolean;
  signal array_obj_ref_250_store_0_ack_1 : boolean;
  signal array_obj_ref_254_gather_scatter_req_0 : boolean;
  signal array_obj_ref_254_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_254_store_0_req_0 : boolean;
  signal array_obj_ref_254_store_0_ack_0 : boolean;
  signal array_obj_ref_254_store_0_req_1 : boolean;
  signal array_obj_ref_254_store_0_ack_1 : boolean;
  signal array_obj_ref_258_gather_scatter_req_0 : boolean;
  signal array_obj_ref_258_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_258_store_0_req_0 : boolean;
  signal array_obj_ref_258_store_0_ack_0 : boolean;
  signal array_obj_ref_258_store_0_req_1 : boolean;
  signal array_obj_ref_258_store_0_ack_1 : boolean;
  signal array_obj_ref_262_gather_scatter_req_0 : boolean;
  signal array_obj_ref_262_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_262_store_0_req_0 : boolean;
  signal array_obj_ref_262_store_0_ack_0 : boolean;
  signal array_obj_ref_262_store_0_req_1 : boolean;
  signal array_obj_ref_262_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 25 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr_CP_402: Block -- control-path 
    signal cp_elements: BooleanArray(75 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(75);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(75), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_166_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_166_gather_scatter_ack_0;
    array_obj_ref_166_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_166_store_0_ack_0;
    array_obj_ref_166_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_166_store_0_ack_1;
    array_obj_ref_170_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_170_gather_scatter_ack_0;
    array_obj_ref_170_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_170_store_0_ack_0;
    array_obj_ref_170_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_170_store_0_ack_1;
    array_obj_ref_174_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_174_gather_scatter_ack_0;
    array_obj_ref_174_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_174_store_0_ack_0;
    array_obj_ref_174_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_174_store_0_ack_1;
    array_obj_ref_178_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_178_gather_scatter_ack_0;
    array_obj_ref_178_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_178_store_0_ack_0;
    array_obj_ref_178_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_178_store_0_ack_1;
    array_obj_ref_182_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_182_gather_scatter_ack_0;
    array_obj_ref_182_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_182_store_0_ack_0;
    array_obj_ref_182_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_182_store_0_ack_1;
    array_obj_ref_186_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_186_gather_scatter_ack_0;
    array_obj_ref_186_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_186_store_0_ack_0;
    array_obj_ref_186_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_186_store_0_ack_1;
    array_obj_ref_190_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_190_gather_scatter_ack_0;
    array_obj_ref_190_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_190_store_0_ack_0;
    array_obj_ref_190_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_190_store_0_ack_1;
    array_obj_ref_194_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_194_gather_scatter_ack_0;
    array_obj_ref_194_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_194_store_0_ack_0;
    array_obj_ref_194_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_194_store_0_ack_1;
    array_obj_ref_198_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_198_gather_scatter_ack_0;
    array_obj_ref_198_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_198_store_0_ack_0;
    array_obj_ref_198_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_198_store_0_ack_1;
    array_obj_ref_202_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_202_gather_scatter_ack_0;
    array_obj_ref_202_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_202_store_0_ack_0;
    array_obj_ref_202_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_202_store_0_ack_1;
    array_obj_ref_206_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_206_gather_scatter_ack_0;
    array_obj_ref_206_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_206_store_0_ack_0;
    array_obj_ref_206_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_206_store_0_ack_1;
    array_obj_ref_210_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_210_gather_scatter_ack_0;
    array_obj_ref_210_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_210_store_0_ack_0;
    array_obj_ref_210_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_210_store_0_ack_1;
    array_obj_ref_214_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_214_gather_scatter_ack_0;
    array_obj_ref_214_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_214_store_0_ack_0;
    array_obj_ref_214_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_214_store_0_ack_1;
    array_obj_ref_218_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_218_gather_scatter_ack_0;
    array_obj_ref_218_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_218_store_0_ack_0;
    array_obj_ref_218_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_218_store_0_ack_1;
    array_obj_ref_222_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_222_gather_scatter_ack_0;
    array_obj_ref_222_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_222_store_0_ack_0;
    array_obj_ref_222_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_222_store_0_ack_1;
    array_obj_ref_226_gather_scatter_req_0 <= cp_elements(45);
    cp_elements(46) <= array_obj_ref_226_gather_scatter_ack_0;
    array_obj_ref_226_store_0_req_0 <= cp_elements(46);
    cp_elements(47) <= array_obj_ref_226_store_0_ack_0;
    array_obj_ref_226_store_0_req_1 <= cp_elements(47);
    cp_elements(48) <= array_obj_ref_226_store_0_ack_1;
    array_obj_ref_230_gather_scatter_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_230_gather_scatter_ack_0;
    array_obj_ref_230_store_0_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_230_store_0_ack_0;
    array_obj_ref_230_store_0_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_230_store_0_ack_1;
    array_obj_ref_234_gather_scatter_req_0 <= cp_elements(51);
    cp_elements(52) <= array_obj_ref_234_gather_scatter_ack_0;
    array_obj_ref_234_store_0_req_0 <= cp_elements(52);
    cp_elements(53) <= array_obj_ref_234_store_0_ack_0;
    array_obj_ref_234_store_0_req_1 <= cp_elements(53);
    cp_elements(54) <= array_obj_ref_234_store_0_ack_1;
    array_obj_ref_238_gather_scatter_req_0 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_238_gather_scatter_ack_0;
    array_obj_ref_238_store_0_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_238_store_0_ack_0;
    array_obj_ref_238_store_0_req_1 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_238_store_0_ack_1;
    array_obj_ref_242_gather_scatter_req_0 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_242_gather_scatter_ack_0;
    array_obj_ref_242_store_0_req_0 <= cp_elements(58);
    cp_elements(59) <= array_obj_ref_242_store_0_ack_0;
    array_obj_ref_242_store_0_req_1 <= cp_elements(59);
    cp_elements(60) <= array_obj_ref_242_store_0_ack_1;
    array_obj_ref_246_gather_scatter_req_0 <= cp_elements(60);
    cp_elements(61) <= array_obj_ref_246_gather_scatter_ack_0;
    array_obj_ref_246_store_0_req_0 <= cp_elements(61);
    cp_elements(62) <= array_obj_ref_246_store_0_ack_0;
    array_obj_ref_246_store_0_req_1 <= cp_elements(62);
    cp_elements(63) <= array_obj_ref_246_store_0_ack_1;
    array_obj_ref_250_gather_scatter_req_0 <= cp_elements(63);
    cp_elements(64) <= array_obj_ref_250_gather_scatter_ack_0;
    array_obj_ref_250_store_0_req_0 <= cp_elements(64);
    cp_elements(65) <= array_obj_ref_250_store_0_ack_0;
    array_obj_ref_250_store_0_req_1 <= cp_elements(65);
    cp_elements(66) <= array_obj_ref_250_store_0_ack_1;
    array_obj_ref_254_gather_scatter_req_0 <= cp_elements(66);
    cp_elements(67) <= array_obj_ref_254_gather_scatter_ack_0;
    array_obj_ref_254_store_0_req_0 <= cp_elements(67);
    cp_elements(68) <= array_obj_ref_254_store_0_ack_0;
    array_obj_ref_254_store_0_req_1 <= cp_elements(68);
    cp_elements(69) <= array_obj_ref_254_store_0_ack_1;
    array_obj_ref_258_gather_scatter_req_0 <= cp_elements(69);
    cp_elements(70) <= array_obj_ref_258_gather_scatter_ack_0;
    array_obj_ref_258_store_0_req_0 <= cp_elements(70);
    cp_elements(71) <= array_obj_ref_258_store_0_ack_0;
    array_obj_ref_258_store_0_req_1 <= cp_elements(71);
    cp_elements(72) <= array_obj_ref_258_store_0_ack_1;
    array_obj_ref_262_gather_scatter_req_0 <= cp_elements(72);
    cp_elements(73) <= array_obj_ref_262_gather_scatter_ack_0;
    array_obj_ref_262_store_0_req_0 <= cp_elements(73);
    cp_elements(74) <= array_obj_ref_262_store_0_ack_0;
    array_obj_ref_262_store_0_req_1 <= cp_elements(74);
    cp_elements(75) <= array_obj_ref_262_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_166_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_170_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_170_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_174_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_174_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_178_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_178_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_182_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_182_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_186_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_186_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_190_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_190_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_194_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_194_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_198_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_198_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_202_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_202_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_206_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_206_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_210_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_210_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_214_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_218_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_218_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_222_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_222_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_226_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_226_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_230_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_230_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_234_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_234_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_238_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_238_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_242_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_242_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_246_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_246_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_250_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_250_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_254_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_254_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_258_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_258_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_262_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_262_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_167_wire_constant : std_logic_vector(7 downto 0);
    signal expr_171_wire_constant : std_logic_vector(7 downto 0);
    signal expr_175_wire_constant : std_logic_vector(7 downto 0);
    signal expr_179_wire_constant : std_logic_vector(7 downto 0);
    signal expr_183_wire_constant : std_logic_vector(7 downto 0);
    signal expr_187_wire_constant : std_logic_vector(7 downto 0);
    signal expr_191_wire_constant : std_logic_vector(7 downto 0);
    signal expr_195_wire_constant : std_logic_vector(7 downto 0);
    signal expr_199_wire_constant : std_logic_vector(7 downto 0);
    signal expr_203_wire_constant : std_logic_vector(7 downto 0);
    signal expr_207_wire_constant : std_logic_vector(7 downto 0);
    signal expr_211_wire_constant : std_logic_vector(7 downto 0);
    signal expr_215_wire_constant : std_logic_vector(7 downto 0);
    signal expr_219_wire_constant : std_logic_vector(7 downto 0);
    signal expr_223_wire_constant : std_logic_vector(7 downto 0);
    signal expr_227_wire_constant : std_logic_vector(7 downto 0);
    signal expr_231_wire_constant : std_logic_vector(7 downto 0);
    signal expr_235_wire_constant : std_logic_vector(7 downto 0);
    signal expr_239_wire_constant : std_logic_vector(7 downto 0);
    signal expr_243_wire_constant : std_logic_vector(7 downto 0);
    signal expr_247_wire_constant : std_logic_vector(7 downto 0);
    signal expr_251_wire_constant : std_logic_vector(7 downto 0);
    signal expr_255_wire_constant : std_logic_vector(7 downto 0);
    signal expr_259_wire_constant : std_logic_vector(7 downto 0);
    signal expr_263_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_166_word_address_0 <= "00000";
    array_obj_ref_170_word_address_0 <= "00001";
    array_obj_ref_174_word_address_0 <= "00010";
    array_obj_ref_178_word_address_0 <= "00011";
    array_obj_ref_182_word_address_0 <= "00100";
    array_obj_ref_186_word_address_0 <= "00101";
    array_obj_ref_190_word_address_0 <= "00110";
    array_obj_ref_194_word_address_0 <= "00111";
    array_obj_ref_198_word_address_0 <= "01000";
    array_obj_ref_202_word_address_0 <= "01001";
    array_obj_ref_206_word_address_0 <= "01010";
    array_obj_ref_210_word_address_0 <= "01011";
    array_obj_ref_214_word_address_0 <= "01100";
    array_obj_ref_218_word_address_0 <= "01101";
    array_obj_ref_222_word_address_0 <= "01110";
    array_obj_ref_226_word_address_0 <= "01111";
    array_obj_ref_230_word_address_0 <= "10000";
    array_obj_ref_234_word_address_0 <= "10001";
    array_obj_ref_238_word_address_0 <= "10010";
    array_obj_ref_242_word_address_0 <= "10011";
    array_obj_ref_246_word_address_0 <= "10100";
    array_obj_ref_250_word_address_0 <= "10101";
    array_obj_ref_254_word_address_0 <= "10110";
    array_obj_ref_258_word_address_0 <= "10111";
    array_obj_ref_262_word_address_0 <= "11000";
    expr_167_wire_constant <= "01110011";
    expr_171_wire_constant <= "01110100";
    expr_175_wire_constant <= "01100001";
    expr_179_wire_constant <= "01110010";
    expr_183_wire_constant <= "01110100";
    expr_187_wire_constant <= "01011111";
    expr_191_wire_constant <= "01101111";
    expr_195_wire_constant <= "01110101";
    expr_199_wire_constant <= "01110100";
    expr_203_wire_constant <= "01110000";
    expr_207_wire_constant <= "01110101";
    expr_211_wire_constant <= "01110100";
    expr_215_wire_constant <= "01011111";
    expr_219_wire_constant <= "01110000";
    expr_223_wire_constant <= "01101111";
    expr_227_wire_constant <= "01110010";
    expr_231_wire_constant <= "01110100";
    expr_235_wire_constant <= "01011111";
    expr_239_wire_constant <= "01101100";
    expr_243_wire_constant <= "01101111";
    expr_247_wire_constant <= "01101111";
    expr_251_wire_constant <= "01101011";
    expr_255_wire_constant <= "01110101";
    expr_259_wire_constant <= "01110000";
    expr_263_wire_constant <= "00000000";
    array_obj_ref_166_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_166_gather_scatter_ack_0 <= array_obj_ref_166_gather_scatter_req_0;
      aggregated_sig <= expr_167_wire_constant;
      array_obj_ref_166_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_170_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_170_gather_scatter_ack_0 <= array_obj_ref_170_gather_scatter_req_0;
      aggregated_sig <= expr_171_wire_constant;
      array_obj_ref_170_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_174_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_174_gather_scatter_ack_0 <= array_obj_ref_174_gather_scatter_req_0;
      aggregated_sig <= expr_175_wire_constant;
      array_obj_ref_174_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_178_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_178_gather_scatter_ack_0 <= array_obj_ref_178_gather_scatter_req_0;
      aggregated_sig <= expr_179_wire_constant;
      array_obj_ref_178_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_182_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_182_gather_scatter_ack_0 <= array_obj_ref_182_gather_scatter_req_0;
      aggregated_sig <= expr_183_wire_constant;
      array_obj_ref_182_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_186_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_186_gather_scatter_ack_0 <= array_obj_ref_186_gather_scatter_req_0;
      aggregated_sig <= expr_187_wire_constant;
      array_obj_ref_186_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_190_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_190_gather_scatter_ack_0 <= array_obj_ref_190_gather_scatter_req_0;
      aggregated_sig <= expr_191_wire_constant;
      array_obj_ref_190_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_194_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_194_gather_scatter_ack_0 <= array_obj_ref_194_gather_scatter_req_0;
      aggregated_sig <= expr_195_wire_constant;
      array_obj_ref_194_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_198_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_198_gather_scatter_ack_0 <= array_obj_ref_198_gather_scatter_req_0;
      aggregated_sig <= expr_199_wire_constant;
      array_obj_ref_198_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_202_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_202_gather_scatter_ack_0 <= array_obj_ref_202_gather_scatter_req_0;
      aggregated_sig <= expr_203_wire_constant;
      array_obj_ref_202_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_206_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_206_gather_scatter_ack_0 <= array_obj_ref_206_gather_scatter_req_0;
      aggregated_sig <= expr_207_wire_constant;
      array_obj_ref_206_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_210_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_210_gather_scatter_ack_0 <= array_obj_ref_210_gather_scatter_req_0;
      aggregated_sig <= expr_211_wire_constant;
      array_obj_ref_210_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_214_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_214_gather_scatter_ack_0 <= array_obj_ref_214_gather_scatter_req_0;
      aggregated_sig <= expr_215_wire_constant;
      array_obj_ref_214_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_218_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_218_gather_scatter_ack_0 <= array_obj_ref_218_gather_scatter_req_0;
      aggregated_sig <= expr_219_wire_constant;
      array_obj_ref_218_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_222_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_222_gather_scatter_ack_0 <= array_obj_ref_222_gather_scatter_req_0;
      aggregated_sig <= expr_223_wire_constant;
      array_obj_ref_222_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_226_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_226_gather_scatter_ack_0 <= array_obj_ref_226_gather_scatter_req_0;
      aggregated_sig <= expr_227_wire_constant;
      array_obj_ref_226_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_230_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_230_gather_scatter_ack_0 <= array_obj_ref_230_gather_scatter_req_0;
      aggregated_sig <= expr_231_wire_constant;
      array_obj_ref_230_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_234_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_234_gather_scatter_ack_0 <= array_obj_ref_234_gather_scatter_req_0;
      aggregated_sig <= expr_235_wire_constant;
      array_obj_ref_234_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_238_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_238_gather_scatter_ack_0 <= array_obj_ref_238_gather_scatter_req_0;
      aggregated_sig <= expr_239_wire_constant;
      array_obj_ref_238_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_242_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_242_gather_scatter_ack_0 <= array_obj_ref_242_gather_scatter_req_0;
      aggregated_sig <= expr_243_wire_constant;
      array_obj_ref_242_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_246_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_246_gather_scatter_ack_0 <= array_obj_ref_246_gather_scatter_req_0;
      aggregated_sig <= expr_247_wire_constant;
      array_obj_ref_246_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_250_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_250_gather_scatter_ack_0 <= array_obj_ref_250_gather_scatter_req_0;
      aggregated_sig <= expr_251_wire_constant;
      array_obj_ref_250_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_254_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_254_gather_scatter_ack_0 <= array_obj_ref_254_gather_scatter_req_0;
      aggregated_sig <= expr_255_wire_constant;
      array_obj_ref_254_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_258_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_258_gather_scatter_ack_0 <= array_obj_ref_258_gather_scatter_req_0;
      aggregated_sig <= expr_259_wire_constant;
      array_obj_ref_258_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_262_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_262_gather_scatter_ack_0 <= array_obj_ref_262_gather_scatter_req_0;
      aggregated_sig <= expr_263_wire_constant;
      array_obj_ref_262_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_234_store_0 array_obj_ref_230_store_0 array_obj_ref_182_store_0 array_obj_ref_250_store_0 array_obj_ref_222_store_0 array_obj_ref_178_store_0 array_obj_ref_218_store_0 array_obj_ref_246_store_0 array_obj_ref_186_store_0 array_obj_ref_214_store_0 array_obj_ref_242_store_0 array_obj_ref_238_store_0 array_obj_ref_210_store_0 array_obj_ref_206_store_0 array_obj_ref_170_store_0 array_obj_ref_254_store_0 array_obj_ref_202_store_0 array_obj_ref_226_store_0 array_obj_ref_166_store_0 array_obj_ref_198_store_0 array_obj_ref_194_store_0 array_obj_ref_174_store_0 array_obj_ref_190_store_0 array_obj_ref_258_store_0 array_obj_ref_262_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(124 downto 0);
      signal data_in: std_logic_vector(199 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 24 downto 0);
      -- 
    begin -- 
      reqL(24) <= array_obj_ref_234_store_0_req_0;
      reqL(23) <= array_obj_ref_230_store_0_req_0;
      reqL(22) <= array_obj_ref_182_store_0_req_0;
      reqL(21) <= array_obj_ref_250_store_0_req_0;
      reqL(20) <= array_obj_ref_222_store_0_req_0;
      reqL(19) <= array_obj_ref_178_store_0_req_0;
      reqL(18) <= array_obj_ref_218_store_0_req_0;
      reqL(17) <= array_obj_ref_246_store_0_req_0;
      reqL(16) <= array_obj_ref_186_store_0_req_0;
      reqL(15) <= array_obj_ref_214_store_0_req_0;
      reqL(14) <= array_obj_ref_242_store_0_req_0;
      reqL(13) <= array_obj_ref_238_store_0_req_0;
      reqL(12) <= array_obj_ref_210_store_0_req_0;
      reqL(11) <= array_obj_ref_206_store_0_req_0;
      reqL(10) <= array_obj_ref_170_store_0_req_0;
      reqL(9) <= array_obj_ref_254_store_0_req_0;
      reqL(8) <= array_obj_ref_202_store_0_req_0;
      reqL(7) <= array_obj_ref_226_store_0_req_0;
      reqL(6) <= array_obj_ref_166_store_0_req_0;
      reqL(5) <= array_obj_ref_198_store_0_req_0;
      reqL(4) <= array_obj_ref_194_store_0_req_0;
      reqL(3) <= array_obj_ref_174_store_0_req_0;
      reqL(2) <= array_obj_ref_190_store_0_req_0;
      reqL(1) <= array_obj_ref_258_store_0_req_0;
      reqL(0) <= array_obj_ref_262_store_0_req_0;
      array_obj_ref_234_store_0_ack_0 <= ackL(24);
      array_obj_ref_230_store_0_ack_0 <= ackL(23);
      array_obj_ref_182_store_0_ack_0 <= ackL(22);
      array_obj_ref_250_store_0_ack_0 <= ackL(21);
      array_obj_ref_222_store_0_ack_0 <= ackL(20);
      array_obj_ref_178_store_0_ack_0 <= ackL(19);
      array_obj_ref_218_store_0_ack_0 <= ackL(18);
      array_obj_ref_246_store_0_ack_0 <= ackL(17);
      array_obj_ref_186_store_0_ack_0 <= ackL(16);
      array_obj_ref_214_store_0_ack_0 <= ackL(15);
      array_obj_ref_242_store_0_ack_0 <= ackL(14);
      array_obj_ref_238_store_0_ack_0 <= ackL(13);
      array_obj_ref_210_store_0_ack_0 <= ackL(12);
      array_obj_ref_206_store_0_ack_0 <= ackL(11);
      array_obj_ref_170_store_0_ack_0 <= ackL(10);
      array_obj_ref_254_store_0_ack_0 <= ackL(9);
      array_obj_ref_202_store_0_ack_0 <= ackL(8);
      array_obj_ref_226_store_0_ack_0 <= ackL(7);
      array_obj_ref_166_store_0_ack_0 <= ackL(6);
      array_obj_ref_198_store_0_ack_0 <= ackL(5);
      array_obj_ref_194_store_0_ack_0 <= ackL(4);
      array_obj_ref_174_store_0_ack_0 <= ackL(3);
      array_obj_ref_190_store_0_ack_0 <= ackL(2);
      array_obj_ref_258_store_0_ack_0 <= ackL(1);
      array_obj_ref_262_store_0_ack_0 <= ackL(0);
      reqR(24) <= array_obj_ref_234_store_0_req_1;
      reqR(23) <= array_obj_ref_230_store_0_req_1;
      reqR(22) <= array_obj_ref_182_store_0_req_1;
      reqR(21) <= array_obj_ref_250_store_0_req_1;
      reqR(20) <= array_obj_ref_222_store_0_req_1;
      reqR(19) <= array_obj_ref_178_store_0_req_1;
      reqR(18) <= array_obj_ref_218_store_0_req_1;
      reqR(17) <= array_obj_ref_246_store_0_req_1;
      reqR(16) <= array_obj_ref_186_store_0_req_1;
      reqR(15) <= array_obj_ref_214_store_0_req_1;
      reqR(14) <= array_obj_ref_242_store_0_req_1;
      reqR(13) <= array_obj_ref_238_store_0_req_1;
      reqR(12) <= array_obj_ref_210_store_0_req_1;
      reqR(11) <= array_obj_ref_206_store_0_req_1;
      reqR(10) <= array_obj_ref_170_store_0_req_1;
      reqR(9) <= array_obj_ref_254_store_0_req_1;
      reqR(8) <= array_obj_ref_202_store_0_req_1;
      reqR(7) <= array_obj_ref_226_store_0_req_1;
      reqR(6) <= array_obj_ref_166_store_0_req_1;
      reqR(5) <= array_obj_ref_198_store_0_req_1;
      reqR(4) <= array_obj_ref_194_store_0_req_1;
      reqR(3) <= array_obj_ref_174_store_0_req_1;
      reqR(2) <= array_obj_ref_190_store_0_req_1;
      reqR(1) <= array_obj_ref_258_store_0_req_1;
      reqR(0) <= array_obj_ref_262_store_0_req_1;
      array_obj_ref_234_store_0_ack_1 <= ackR(24);
      array_obj_ref_230_store_0_ack_1 <= ackR(23);
      array_obj_ref_182_store_0_ack_1 <= ackR(22);
      array_obj_ref_250_store_0_ack_1 <= ackR(21);
      array_obj_ref_222_store_0_ack_1 <= ackR(20);
      array_obj_ref_178_store_0_ack_1 <= ackR(19);
      array_obj_ref_218_store_0_ack_1 <= ackR(18);
      array_obj_ref_246_store_0_ack_1 <= ackR(17);
      array_obj_ref_186_store_0_ack_1 <= ackR(16);
      array_obj_ref_214_store_0_ack_1 <= ackR(15);
      array_obj_ref_242_store_0_ack_1 <= ackR(14);
      array_obj_ref_238_store_0_ack_1 <= ackR(13);
      array_obj_ref_210_store_0_ack_1 <= ackR(12);
      array_obj_ref_206_store_0_ack_1 <= ackR(11);
      array_obj_ref_170_store_0_ack_1 <= ackR(10);
      array_obj_ref_254_store_0_ack_1 <= ackR(9);
      array_obj_ref_202_store_0_ack_1 <= ackR(8);
      array_obj_ref_226_store_0_ack_1 <= ackR(7);
      array_obj_ref_166_store_0_ack_1 <= ackR(6);
      array_obj_ref_198_store_0_ack_1 <= ackR(5);
      array_obj_ref_194_store_0_ack_1 <= ackR(4);
      array_obj_ref_174_store_0_ack_1 <= ackR(3);
      array_obj_ref_190_store_0_ack_1 <= ackR(2);
      array_obj_ref_258_store_0_ack_1 <= ackR(1);
      array_obj_ref_262_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_234_word_address_0 & array_obj_ref_230_word_address_0 & array_obj_ref_182_word_address_0 & array_obj_ref_250_word_address_0 & array_obj_ref_222_word_address_0 & array_obj_ref_178_word_address_0 & array_obj_ref_218_word_address_0 & array_obj_ref_246_word_address_0 & array_obj_ref_186_word_address_0 & array_obj_ref_214_word_address_0 & array_obj_ref_242_word_address_0 & array_obj_ref_238_word_address_0 & array_obj_ref_210_word_address_0 & array_obj_ref_206_word_address_0 & array_obj_ref_170_word_address_0 & array_obj_ref_254_word_address_0 & array_obj_ref_202_word_address_0 & array_obj_ref_226_word_address_0 & array_obj_ref_166_word_address_0 & array_obj_ref_198_word_address_0 & array_obj_ref_194_word_address_0 & array_obj_ref_174_word_address_0 & array_obj_ref_190_word_address_0 & array_obj_ref_258_word_address_0 & array_obj_ref_262_word_address_0;
      data_in <= array_obj_ref_234_data_0 & array_obj_ref_230_data_0 & array_obj_ref_182_data_0 & array_obj_ref_250_data_0 & array_obj_ref_222_data_0 & array_obj_ref_178_data_0 & array_obj_ref_218_data_0 & array_obj_ref_246_data_0 & array_obj_ref_186_data_0 & array_obj_ref_214_data_0 & array_obj_ref_242_data_0 & array_obj_ref_238_data_0 & array_obj_ref_210_data_0 & array_obj_ref_206_data_0 & array_obj_ref_170_data_0 & array_obj_ref_254_data_0 & array_obj_ref_202_data_0 & array_obj_ref_226_data_0 & array_obj_ref_166_data_0 & array_obj_ref_198_data_0 & array_obj_ref_194_data_0 & array_obj_ref_174_data_0 & array_obj_ref_190_data_0 & array_obj_ref_258_data_0 & array_obj_ref_262_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 8,
        num_reqs => 25,
        tag_length => 5,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(4 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 25,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr1;
architecture Default of default_initializer_xx_xstr1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr1_CP_930_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_276_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_0 : boolean;
  signal array_obj_ref_276_store_0_ack_0 : boolean;
  signal array_obj_ref_272_gather_scatter_req_0 : boolean;
  signal array_obj_ref_272_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_268_store_0_req_0 : boolean;
  signal array_obj_ref_268_store_0_ack_0 : boolean;
  signal array_obj_ref_268_store_0_req_1 : boolean;
  signal array_obj_ref_268_store_0_ack_1 : boolean;
  signal array_obj_ref_280_store_0_req_0 : boolean;
  signal array_obj_ref_280_store_0_ack_0 : boolean;
  signal array_obj_ref_280_store_0_req_1 : boolean;
  signal array_obj_ref_280_store_0_ack_1 : boolean;
  signal array_obj_ref_276_store_0_req_1 : boolean;
  signal array_obj_ref_276_store_0_ack_1 : boolean;
  signal array_obj_ref_272_store_0_req_0 : boolean;
  signal array_obj_ref_272_store_0_ack_0 : boolean;
  signal array_obj_ref_272_store_0_req_1 : boolean;
  signal array_obj_ref_272_store_0_ack_1 : boolean;
  signal array_obj_ref_284_gather_scatter_req_0 : boolean;
  signal array_obj_ref_284_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_268_gather_scatter_req_0 : boolean;
  signal array_obj_ref_268_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_280_gather_scatter_req_0 : boolean;
  signal array_obj_ref_280_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_276_gather_scatter_req_0 : boolean;
  signal array_obj_ref_284_store_0_req_0 : boolean;
  signal array_obj_ref_284_store_0_ack_0 : boolean;
  signal array_obj_ref_284_store_0_req_1 : boolean;
  signal array_obj_ref_284_store_0_ack_1 : boolean;
  signal array_obj_ref_288_gather_scatter_req_0 : boolean;
  signal array_obj_ref_288_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_288_store_0_req_0 : boolean;
  signal array_obj_ref_288_store_0_ack_0 : boolean;
  signal array_obj_ref_288_store_0_req_1 : boolean;
  signal array_obj_ref_288_store_0_ack_1 : boolean;
  signal array_obj_ref_292_gather_scatter_req_0 : boolean;
  signal array_obj_ref_292_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_292_store_0_req_0 : boolean;
  signal array_obj_ref_292_store_0_ack_0 : boolean;
  signal array_obj_ref_292_store_0_req_1 : boolean;
  signal array_obj_ref_292_store_0_ack_1 : boolean;
  signal array_obj_ref_296_gather_scatter_req_0 : boolean;
  signal array_obj_ref_296_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_296_store_0_req_0 : boolean;
  signal array_obj_ref_296_store_0_ack_0 : boolean;
  signal array_obj_ref_296_store_0_req_1 : boolean;
  signal array_obj_ref_296_store_0_ack_1 : boolean;
  signal array_obj_ref_300_gather_scatter_req_0 : boolean;
  signal array_obj_ref_300_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_300_store_0_req_0 : boolean;
  signal array_obj_ref_300_store_0_ack_0 : boolean;
  signal array_obj_ref_300_store_0_req_1 : boolean;
  signal array_obj_ref_300_store_0_ack_1 : boolean;
  signal array_obj_ref_304_gather_scatter_req_0 : boolean;
  signal array_obj_ref_304_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_304_store_0_req_0 : boolean;
  signal array_obj_ref_304_store_0_ack_0 : boolean;
  signal array_obj_ref_304_store_0_req_1 : boolean;
  signal array_obj_ref_304_store_0_ack_1 : boolean;
  signal array_obj_ref_308_gather_scatter_req_0 : boolean;
  signal array_obj_ref_308_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_308_store_0_req_0 : boolean;
  signal array_obj_ref_308_store_0_ack_0 : boolean;
  signal array_obj_ref_308_store_0_req_1 : boolean;
  signal array_obj_ref_308_store_0_ack_1 : boolean;
  signal array_obj_ref_312_gather_scatter_req_0 : boolean;
  signal array_obj_ref_312_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_312_store_0_req_0 : boolean;
  signal array_obj_ref_312_store_0_ack_0 : boolean;
  signal array_obj_ref_312_store_0_req_1 : boolean;
  signal array_obj_ref_312_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 12 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr1_CP_930: Block -- control-path 
    signal cp_elements: BooleanArray(36 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(36);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(36), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_268_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_268_gather_scatter_ack_0;
    array_obj_ref_268_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_268_store_0_ack_0;
    array_obj_ref_268_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_268_store_0_ack_1;
    array_obj_ref_272_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_272_gather_scatter_ack_0;
    array_obj_ref_272_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_272_store_0_ack_0;
    array_obj_ref_272_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_272_store_0_ack_1;
    array_obj_ref_276_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_276_gather_scatter_ack_0;
    array_obj_ref_276_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_276_store_0_ack_0;
    array_obj_ref_276_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_276_store_0_ack_1;
    array_obj_ref_280_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_280_gather_scatter_ack_0;
    array_obj_ref_280_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_280_store_0_ack_0;
    array_obj_ref_280_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_280_store_0_ack_1;
    array_obj_ref_284_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_284_gather_scatter_ack_0;
    array_obj_ref_284_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_284_store_0_ack_0;
    array_obj_ref_284_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_284_store_0_ack_1;
    array_obj_ref_288_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_288_gather_scatter_ack_0;
    array_obj_ref_288_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_288_store_0_ack_0;
    array_obj_ref_288_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_288_store_0_ack_1;
    array_obj_ref_292_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_292_gather_scatter_ack_0;
    array_obj_ref_292_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_292_store_0_ack_0;
    array_obj_ref_292_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_292_store_0_ack_1;
    array_obj_ref_296_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_296_gather_scatter_ack_0;
    array_obj_ref_296_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_296_store_0_ack_0;
    array_obj_ref_296_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_296_store_0_ack_1;
    array_obj_ref_300_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_300_gather_scatter_ack_0;
    array_obj_ref_300_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_300_store_0_ack_0;
    array_obj_ref_300_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_300_store_0_ack_1;
    array_obj_ref_304_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_304_gather_scatter_ack_0;
    array_obj_ref_304_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_304_store_0_ack_0;
    array_obj_ref_304_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_304_store_0_ack_1;
    array_obj_ref_308_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_308_gather_scatter_ack_0;
    array_obj_ref_308_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_308_store_0_ack_0;
    array_obj_ref_308_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_308_store_0_ack_1;
    array_obj_ref_312_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_312_gather_scatter_ack_0;
    array_obj_ref_312_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_312_store_0_ack_0;
    array_obj_ref_312_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_312_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_268_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_268_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_272_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_272_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_276_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_276_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_280_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_280_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_284_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_284_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_288_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_288_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_292_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_292_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_296_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_296_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_300_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_300_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_304_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_304_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_308_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_308_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_312_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_312_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_269_wire_constant : std_logic_vector(7 downto 0);
    signal expr_273_wire_constant : std_logic_vector(7 downto 0);
    signal expr_277_wire_constant : std_logic_vector(7 downto 0);
    signal expr_281_wire_constant : std_logic_vector(7 downto 0);
    signal expr_285_wire_constant : std_logic_vector(7 downto 0);
    signal expr_289_wire_constant : std_logic_vector(7 downto 0);
    signal expr_293_wire_constant : std_logic_vector(7 downto 0);
    signal expr_297_wire_constant : std_logic_vector(7 downto 0);
    signal expr_301_wire_constant : std_logic_vector(7 downto 0);
    signal expr_305_wire_constant : std_logic_vector(7 downto 0);
    signal expr_309_wire_constant : std_logic_vector(7 downto 0);
    signal expr_313_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_268_word_address_0 <= "0000";
    array_obj_ref_272_word_address_0 <= "0001";
    array_obj_ref_276_word_address_0 <= "0010";
    array_obj_ref_280_word_address_0 <= "0011";
    array_obj_ref_284_word_address_0 <= "0100";
    array_obj_ref_288_word_address_0 <= "0101";
    array_obj_ref_292_word_address_0 <= "0110";
    array_obj_ref_296_word_address_0 <= "0111";
    array_obj_ref_300_word_address_0 <= "1000";
    array_obj_ref_304_word_address_0 <= "1001";
    array_obj_ref_308_word_address_0 <= "1010";
    array_obj_ref_312_word_address_0 <= "1011";
    expr_269_wire_constant <= "01101111";
    expr_273_wire_constant <= "01110000";
    expr_277_wire_constant <= "01011111";
    expr_281_wire_constant <= "01101100";
    expr_285_wire_constant <= "01110101";
    expr_289_wire_constant <= "01110100";
    expr_293_wire_constant <= "01011111";
    expr_297_wire_constant <= "01100011";
    expr_301_wire_constant <= "01110100";
    expr_305_wire_constant <= "01110010";
    expr_309_wire_constant <= "01101100";
    expr_313_wire_constant <= "00000000";
    array_obj_ref_268_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_268_gather_scatter_ack_0 <= array_obj_ref_268_gather_scatter_req_0;
      aggregated_sig <= expr_269_wire_constant;
      array_obj_ref_268_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_272_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_272_gather_scatter_ack_0 <= array_obj_ref_272_gather_scatter_req_0;
      aggregated_sig <= expr_273_wire_constant;
      array_obj_ref_272_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_276_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_276_gather_scatter_ack_0 <= array_obj_ref_276_gather_scatter_req_0;
      aggregated_sig <= expr_277_wire_constant;
      array_obj_ref_276_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_280_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_280_gather_scatter_ack_0 <= array_obj_ref_280_gather_scatter_req_0;
      aggregated_sig <= expr_281_wire_constant;
      array_obj_ref_280_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_284_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_284_gather_scatter_ack_0 <= array_obj_ref_284_gather_scatter_req_0;
      aggregated_sig <= expr_285_wire_constant;
      array_obj_ref_284_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_288_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_288_gather_scatter_ack_0 <= array_obj_ref_288_gather_scatter_req_0;
      aggregated_sig <= expr_289_wire_constant;
      array_obj_ref_288_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_292_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_292_gather_scatter_ack_0 <= array_obj_ref_292_gather_scatter_req_0;
      aggregated_sig <= expr_293_wire_constant;
      array_obj_ref_292_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_296_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_296_gather_scatter_ack_0 <= array_obj_ref_296_gather_scatter_req_0;
      aggregated_sig <= expr_297_wire_constant;
      array_obj_ref_296_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_300_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_300_gather_scatter_ack_0 <= array_obj_ref_300_gather_scatter_req_0;
      aggregated_sig <= expr_301_wire_constant;
      array_obj_ref_300_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_304_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_304_gather_scatter_ack_0 <= array_obj_ref_304_gather_scatter_req_0;
      aggregated_sig <= expr_305_wire_constant;
      array_obj_ref_304_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_308_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_308_gather_scatter_ack_0 <= array_obj_ref_308_gather_scatter_req_0;
      aggregated_sig <= expr_309_wire_constant;
      array_obj_ref_308_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_312_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_312_gather_scatter_ack_0 <= array_obj_ref_312_gather_scatter_req_0;
      aggregated_sig <= expr_313_wire_constant;
      array_obj_ref_312_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_268_store_0 array_obj_ref_272_store_0 array_obj_ref_276_store_0 array_obj_ref_280_store_0 array_obj_ref_284_store_0 array_obj_ref_288_store_0 array_obj_ref_292_store_0 array_obj_ref_296_store_0 array_obj_ref_300_store_0 array_obj_ref_304_store_0 array_obj_ref_308_store_0 array_obj_ref_312_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(47 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      reqL(11) <= array_obj_ref_268_store_0_req_0;
      reqL(10) <= array_obj_ref_272_store_0_req_0;
      reqL(9) <= array_obj_ref_276_store_0_req_0;
      reqL(8) <= array_obj_ref_280_store_0_req_0;
      reqL(7) <= array_obj_ref_284_store_0_req_0;
      reqL(6) <= array_obj_ref_288_store_0_req_0;
      reqL(5) <= array_obj_ref_292_store_0_req_0;
      reqL(4) <= array_obj_ref_296_store_0_req_0;
      reqL(3) <= array_obj_ref_300_store_0_req_0;
      reqL(2) <= array_obj_ref_304_store_0_req_0;
      reqL(1) <= array_obj_ref_308_store_0_req_0;
      reqL(0) <= array_obj_ref_312_store_0_req_0;
      array_obj_ref_268_store_0_ack_0 <= ackL(11);
      array_obj_ref_272_store_0_ack_0 <= ackL(10);
      array_obj_ref_276_store_0_ack_0 <= ackL(9);
      array_obj_ref_280_store_0_ack_0 <= ackL(8);
      array_obj_ref_284_store_0_ack_0 <= ackL(7);
      array_obj_ref_288_store_0_ack_0 <= ackL(6);
      array_obj_ref_292_store_0_ack_0 <= ackL(5);
      array_obj_ref_296_store_0_ack_0 <= ackL(4);
      array_obj_ref_300_store_0_ack_0 <= ackL(3);
      array_obj_ref_304_store_0_ack_0 <= ackL(2);
      array_obj_ref_308_store_0_ack_0 <= ackL(1);
      array_obj_ref_312_store_0_ack_0 <= ackL(0);
      reqR(11) <= array_obj_ref_268_store_0_req_1;
      reqR(10) <= array_obj_ref_272_store_0_req_1;
      reqR(9) <= array_obj_ref_276_store_0_req_1;
      reqR(8) <= array_obj_ref_280_store_0_req_1;
      reqR(7) <= array_obj_ref_284_store_0_req_1;
      reqR(6) <= array_obj_ref_288_store_0_req_1;
      reqR(5) <= array_obj_ref_292_store_0_req_1;
      reqR(4) <= array_obj_ref_296_store_0_req_1;
      reqR(3) <= array_obj_ref_300_store_0_req_1;
      reqR(2) <= array_obj_ref_304_store_0_req_1;
      reqR(1) <= array_obj_ref_308_store_0_req_1;
      reqR(0) <= array_obj_ref_312_store_0_req_1;
      array_obj_ref_268_store_0_ack_1 <= ackR(11);
      array_obj_ref_272_store_0_ack_1 <= ackR(10);
      array_obj_ref_276_store_0_ack_1 <= ackR(9);
      array_obj_ref_280_store_0_ack_1 <= ackR(8);
      array_obj_ref_284_store_0_ack_1 <= ackR(7);
      array_obj_ref_288_store_0_ack_1 <= ackR(6);
      array_obj_ref_292_store_0_ack_1 <= ackR(5);
      array_obj_ref_296_store_0_ack_1 <= ackR(4);
      array_obj_ref_300_store_0_ack_1 <= ackR(3);
      array_obj_ref_304_store_0_ack_1 <= ackR(2);
      array_obj_ref_308_store_0_ack_1 <= ackR(1);
      array_obj_ref_312_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_268_word_address_0 & array_obj_ref_272_word_address_0 & array_obj_ref_276_word_address_0 & array_obj_ref_280_word_address_0 & array_obj_ref_284_word_address_0 & array_obj_ref_288_word_address_0 & array_obj_ref_292_word_address_0 & array_obj_ref_296_word_address_0 & array_obj_ref_300_word_address_0 & array_obj_ref_304_word_address_0 & array_obj_ref_308_word_address_0 & array_obj_ref_312_word_address_0;
      data_in <= array_obj_ref_268_data_0 & array_obj_ref_272_data_0 & array_obj_ref_276_data_0 & array_obj_ref_280_data_0 & array_obj_ref_284_data_0 & array_obj_ref_288_data_0 & array_obj_ref_292_data_0 & array_obj_ref_296_data_0 & array_obj_ref_300_data_0 & array_obj_ref_304_data_0 & array_obj_ref_308_data_0 & array_obj_ref_312_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 12,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(3 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 12,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr10 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr10;
architecture Default of default_initializer_xx_xstr10 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr10_CP_1185_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_394_store_0_req_1 : boolean;
  signal array_obj_ref_394_store_0_ack_0 : boolean;
  signal array_obj_ref_398_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_398_store_0_ack_1 : boolean;
  signal array_obj_ref_394_store_0_req_0 : boolean;
  signal array_obj_ref_398_gather_scatter_req_0 : boolean;
  signal array_obj_ref_398_store_0_req_0 : boolean;
  signal array_obj_ref_394_store_0_ack_1 : boolean;
  signal array_obj_ref_398_store_0_ack_0 : boolean;
  signal array_obj_ref_398_store_0_req_1 : boolean;
  signal array_obj_ref_318_gather_scatter_req_0 : boolean;
  signal array_obj_ref_318_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_0 : boolean;
  signal array_obj_ref_318_store_0_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_1 : boolean;
  signal array_obj_ref_318_store_0_ack_1 : boolean;
  signal array_obj_ref_322_gather_scatter_req_0 : boolean;
  signal array_obj_ref_322_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_322_store_0_req_0 : boolean;
  signal array_obj_ref_322_store_0_ack_0 : boolean;
  signal array_obj_ref_322_store_0_req_1 : boolean;
  signal array_obj_ref_322_store_0_ack_1 : boolean;
  signal array_obj_ref_326_gather_scatter_req_0 : boolean;
  signal array_obj_ref_326_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_326_store_0_req_0 : boolean;
  signal array_obj_ref_326_store_0_ack_0 : boolean;
  signal array_obj_ref_326_store_0_req_1 : boolean;
  signal array_obj_ref_326_store_0_ack_1 : boolean;
  signal array_obj_ref_330_gather_scatter_req_0 : boolean;
  signal array_obj_ref_330_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_330_store_0_req_0 : boolean;
  signal array_obj_ref_330_store_0_ack_0 : boolean;
  signal array_obj_ref_330_store_0_req_1 : boolean;
  signal array_obj_ref_330_store_0_ack_1 : boolean;
  signal array_obj_ref_334_gather_scatter_req_0 : boolean;
  signal array_obj_ref_334_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_334_store_0_req_0 : boolean;
  signal array_obj_ref_334_store_0_ack_0 : boolean;
  signal array_obj_ref_334_store_0_req_1 : boolean;
  signal array_obj_ref_334_store_0_ack_1 : boolean;
  signal array_obj_ref_338_gather_scatter_req_0 : boolean;
  signal array_obj_ref_338_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_338_store_0_req_0 : boolean;
  signal array_obj_ref_338_store_0_ack_0 : boolean;
  signal array_obj_ref_338_store_0_req_1 : boolean;
  signal array_obj_ref_338_store_0_ack_1 : boolean;
  signal array_obj_ref_342_gather_scatter_req_0 : boolean;
  signal array_obj_ref_342_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_342_store_0_req_0 : boolean;
  signal array_obj_ref_342_store_0_ack_0 : boolean;
  signal array_obj_ref_342_store_0_req_1 : boolean;
  signal array_obj_ref_342_store_0_ack_1 : boolean;
  signal array_obj_ref_346_gather_scatter_req_0 : boolean;
  signal array_obj_ref_346_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_0 : boolean;
  signal array_obj_ref_346_store_0_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_1 : boolean;
  signal array_obj_ref_346_store_0_ack_1 : boolean;
  signal array_obj_ref_350_gather_scatter_req_0 : boolean;
  signal array_obj_ref_350_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_350_store_0_req_0 : boolean;
  signal array_obj_ref_350_store_0_ack_0 : boolean;
  signal array_obj_ref_350_store_0_req_1 : boolean;
  signal array_obj_ref_350_store_0_ack_1 : boolean;
  signal array_obj_ref_354_gather_scatter_req_0 : boolean;
  signal array_obj_ref_354_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_354_store_0_req_0 : boolean;
  signal array_obj_ref_354_store_0_ack_0 : boolean;
  signal array_obj_ref_354_store_0_req_1 : boolean;
  signal array_obj_ref_354_store_0_ack_1 : boolean;
  signal array_obj_ref_358_gather_scatter_req_0 : boolean;
  signal array_obj_ref_358_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_358_store_0_req_0 : boolean;
  signal array_obj_ref_358_store_0_ack_0 : boolean;
  signal array_obj_ref_358_store_0_req_1 : boolean;
  signal array_obj_ref_358_store_0_ack_1 : boolean;
  signal array_obj_ref_362_gather_scatter_req_0 : boolean;
  signal array_obj_ref_362_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_362_store_0_req_0 : boolean;
  signal array_obj_ref_362_store_0_ack_0 : boolean;
  signal array_obj_ref_362_store_0_req_1 : boolean;
  signal array_obj_ref_362_store_0_ack_1 : boolean;
  signal array_obj_ref_366_gather_scatter_req_0 : boolean;
  signal array_obj_ref_366_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_366_store_0_req_0 : boolean;
  signal array_obj_ref_366_store_0_ack_0 : boolean;
  signal array_obj_ref_366_store_0_req_1 : boolean;
  signal array_obj_ref_366_store_0_ack_1 : boolean;
  signal array_obj_ref_370_gather_scatter_req_0 : boolean;
  signal array_obj_ref_370_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_370_store_0_req_0 : boolean;
  signal array_obj_ref_370_store_0_ack_0 : boolean;
  signal array_obj_ref_370_store_0_req_1 : boolean;
  signal array_obj_ref_370_store_0_ack_1 : boolean;
  signal array_obj_ref_374_gather_scatter_req_0 : boolean;
  signal array_obj_ref_374_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_374_store_0_req_0 : boolean;
  signal array_obj_ref_374_store_0_ack_0 : boolean;
  signal array_obj_ref_374_store_0_req_1 : boolean;
  signal array_obj_ref_374_store_0_ack_1 : boolean;
  signal array_obj_ref_378_gather_scatter_req_0 : boolean;
  signal array_obj_ref_378_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_378_store_0_req_0 : boolean;
  signal array_obj_ref_378_store_0_ack_0 : boolean;
  signal array_obj_ref_378_store_0_req_1 : boolean;
  signal array_obj_ref_378_store_0_ack_1 : boolean;
  signal array_obj_ref_382_gather_scatter_req_0 : boolean;
  signal array_obj_ref_382_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_382_store_0_req_0 : boolean;
  signal array_obj_ref_382_store_0_ack_0 : boolean;
  signal array_obj_ref_382_store_0_req_1 : boolean;
  signal array_obj_ref_382_store_0_ack_1 : boolean;
  signal array_obj_ref_386_gather_scatter_req_0 : boolean;
  signal array_obj_ref_386_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_386_store_0_req_0 : boolean;
  signal array_obj_ref_386_store_0_ack_0 : boolean;
  signal array_obj_ref_386_store_0_req_1 : boolean;
  signal array_obj_ref_386_store_0_ack_1 : boolean;
  signal array_obj_ref_390_gather_scatter_req_0 : boolean;
  signal array_obj_ref_390_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_390_store_0_req_0 : boolean;
  signal array_obj_ref_390_store_0_ack_0 : boolean;
  signal array_obj_ref_390_store_0_req_1 : boolean;
  signal array_obj_ref_390_store_0_ack_1 : boolean;
  signal array_obj_ref_394_gather_scatter_req_0 : boolean;
  signal array_obj_ref_394_gather_scatter_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 21 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr10_CP_1185: Block -- control-path 
    signal cp_elements: BooleanArray(63 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(63);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(63), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_318_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_318_gather_scatter_ack_0;
    array_obj_ref_318_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_318_store_0_ack_0;
    array_obj_ref_318_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_318_store_0_ack_1;
    array_obj_ref_322_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_322_gather_scatter_ack_0;
    array_obj_ref_322_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_322_store_0_ack_0;
    array_obj_ref_322_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_322_store_0_ack_1;
    array_obj_ref_326_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_326_gather_scatter_ack_0;
    array_obj_ref_326_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_326_store_0_ack_0;
    array_obj_ref_326_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_326_store_0_ack_1;
    array_obj_ref_330_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_330_gather_scatter_ack_0;
    array_obj_ref_330_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_330_store_0_ack_0;
    array_obj_ref_330_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_330_store_0_ack_1;
    array_obj_ref_334_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_334_gather_scatter_ack_0;
    array_obj_ref_334_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_334_store_0_ack_0;
    array_obj_ref_334_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_334_store_0_ack_1;
    array_obj_ref_338_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_338_gather_scatter_ack_0;
    array_obj_ref_338_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_338_store_0_ack_0;
    array_obj_ref_338_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_338_store_0_ack_1;
    array_obj_ref_342_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_342_gather_scatter_ack_0;
    array_obj_ref_342_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_342_store_0_ack_0;
    array_obj_ref_342_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_342_store_0_ack_1;
    array_obj_ref_346_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_346_gather_scatter_ack_0;
    array_obj_ref_346_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_346_store_0_ack_0;
    array_obj_ref_346_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_346_store_0_ack_1;
    array_obj_ref_350_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_350_gather_scatter_ack_0;
    array_obj_ref_350_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_350_store_0_ack_0;
    array_obj_ref_350_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_350_store_0_ack_1;
    array_obj_ref_354_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_354_gather_scatter_ack_0;
    array_obj_ref_354_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_354_store_0_ack_0;
    array_obj_ref_354_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_354_store_0_ack_1;
    array_obj_ref_358_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_358_gather_scatter_ack_0;
    array_obj_ref_358_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_358_store_0_ack_0;
    array_obj_ref_358_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_358_store_0_ack_1;
    array_obj_ref_362_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_362_gather_scatter_ack_0;
    array_obj_ref_362_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_362_store_0_ack_0;
    array_obj_ref_362_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_362_store_0_ack_1;
    array_obj_ref_366_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_366_gather_scatter_ack_0;
    array_obj_ref_366_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_366_store_0_ack_0;
    array_obj_ref_366_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_366_store_0_ack_1;
    array_obj_ref_370_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_370_gather_scatter_ack_0;
    array_obj_ref_370_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_370_store_0_ack_0;
    array_obj_ref_370_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_370_store_0_ack_1;
    array_obj_ref_374_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_374_gather_scatter_ack_0;
    array_obj_ref_374_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_374_store_0_ack_0;
    array_obj_ref_374_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_374_store_0_ack_1;
    array_obj_ref_378_gather_scatter_req_0 <= cp_elements(45);
    cp_elements(46) <= array_obj_ref_378_gather_scatter_ack_0;
    array_obj_ref_378_store_0_req_0 <= cp_elements(46);
    cp_elements(47) <= array_obj_ref_378_store_0_ack_0;
    array_obj_ref_378_store_0_req_1 <= cp_elements(47);
    cp_elements(48) <= array_obj_ref_378_store_0_ack_1;
    array_obj_ref_382_gather_scatter_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_382_gather_scatter_ack_0;
    array_obj_ref_382_store_0_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_382_store_0_ack_0;
    array_obj_ref_382_store_0_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_382_store_0_ack_1;
    array_obj_ref_386_gather_scatter_req_0 <= cp_elements(51);
    cp_elements(52) <= array_obj_ref_386_gather_scatter_ack_0;
    array_obj_ref_386_store_0_req_0 <= cp_elements(52);
    cp_elements(53) <= array_obj_ref_386_store_0_ack_0;
    array_obj_ref_386_store_0_req_1 <= cp_elements(53);
    cp_elements(54) <= array_obj_ref_386_store_0_ack_1;
    array_obj_ref_390_gather_scatter_req_0 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_390_gather_scatter_ack_0;
    array_obj_ref_390_store_0_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_390_store_0_ack_0;
    array_obj_ref_390_store_0_req_1 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_390_store_0_ack_1;
    array_obj_ref_394_gather_scatter_req_0 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_394_gather_scatter_ack_0;
    array_obj_ref_394_store_0_req_0 <= cp_elements(58);
    cp_elements(59) <= array_obj_ref_394_store_0_ack_0;
    array_obj_ref_394_store_0_req_1 <= cp_elements(59);
    cp_elements(60) <= array_obj_ref_394_store_0_ack_1;
    array_obj_ref_398_gather_scatter_req_0 <= cp_elements(60);
    cp_elements(61) <= array_obj_ref_398_gather_scatter_ack_0;
    array_obj_ref_398_store_0_req_0 <= cp_elements(61);
    cp_elements(62) <= array_obj_ref_398_store_0_ack_0;
    array_obj_ref_398_store_0_req_1 <= cp_elements(62);
    cp_elements(63) <= array_obj_ref_398_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_318_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_318_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_322_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_322_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_326_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_326_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_330_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_330_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_334_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_334_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_338_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_338_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_342_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_342_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_346_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_346_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_350_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_350_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_354_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_354_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_358_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_358_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_362_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_362_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_366_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_366_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_370_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_370_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_374_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_374_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_378_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_378_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_382_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_382_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_386_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_386_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_390_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_390_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_394_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_394_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_398_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_398_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_319_wire_constant : std_logic_vector(7 downto 0);
    signal expr_323_wire_constant : std_logic_vector(7 downto 0);
    signal expr_327_wire_constant : std_logic_vector(7 downto 0);
    signal expr_331_wire_constant : std_logic_vector(7 downto 0);
    signal expr_335_wire_constant : std_logic_vector(7 downto 0);
    signal expr_339_wire_constant : std_logic_vector(7 downto 0);
    signal expr_343_wire_constant : std_logic_vector(7 downto 0);
    signal expr_347_wire_constant : std_logic_vector(7 downto 0);
    signal expr_351_wire_constant : std_logic_vector(7 downto 0);
    signal expr_355_wire_constant : std_logic_vector(7 downto 0);
    signal expr_359_wire_constant : std_logic_vector(7 downto 0);
    signal expr_363_wire_constant : std_logic_vector(7 downto 0);
    signal expr_367_wire_constant : std_logic_vector(7 downto 0);
    signal expr_371_wire_constant : std_logic_vector(7 downto 0);
    signal expr_375_wire_constant : std_logic_vector(7 downto 0);
    signal expr_379_wire_constant : std_logic_vector(7 downto 0);
    signal expr_383_wire_constant : std_logic_vector(7 downto 0);
    signal expr_387_wire_constant : std_logic_vector(7 downto 0);
    signal expr_391_wire_constant : std_logic_vector(7 downto 0);
    signal expr_395_wire_constant : std_logic_vector(7 downto 0);
    signal expr_399_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_318_word_address_0 <= "00000";
    array_obj_ref_322_word_address_0 <= "00001";
    array_obj_ref_326_word_address_0 <= "00010";
    array_obj_ref_330_word_address_0 <= "00011";
    array_obj_ref_334_word_address_0 <= "00100";
    array_obj_ref_338_word_address_0 <= "00101";
    array_obj_ref_342_word_address_0 <= "00110";
    array_obj_ref_346_word_address_0 <= "00111";
    array_obj_ref_350_word_address_0 <= "01000";
    array_obj_ref_354_word_address_0 <= "01001";
    array_obj_ref_358_word_address_0 <= "01010";
    array_obj_ref_362_word_address_0 <= "01011";
    array_obj_ref_366_word_address_0 <= "01100";
    array_obj_ref_370_word_address_0 <= "01101";
    array_obj_ref_374_word_address_0 <= "01110";
    array_obj_ref_378_word_address_0 <= "01111";
    array_obj_ref_382_word_address_0 <= "10000";
    array_obj_ref_386_word_address_0 <= "10001";
    array_obj_ref_390_word_address_0 <= "10010";
    array_obj_ref_394_word_address_0 <= "10011";
    array_obj_ref_398_word_address_0 <= "10100";
    expr_319_wire_constant <= "01110011";
    expr_323_wire_constant <= "01110100";
    expr_327_wire_constant <= "01100001";
    expr_331_wire_constant <= "01110010";
    expr_335_wire_constant <= "01110100";
    expr_339_wire_constant <= "01011111";
    expr_343_wire_constant <= "01110111";
    expr_347_wire_constant <= "01110010";
    expr_351_wire_constant <= "01100001";
    expr_355_wire_constant <= "01110000";
    expr_359_wire_constant <= "01110000";
    expr_363_wire_constant <= "01100101";
    expr_367_wire_constant <= "01110010";
    expr_371_wire_constant <= "01011111";
    expr_375_wire_constant <= "01101111";
    expr_379_wire_constant <= "01110101";
    expr_383_wire_constant <= "01110100";
    expr_387_wire_constant <= "01110000";
    expr_391_wire_constant <= "01110101";
    expr_395_wire_constant <= "01110100";
    expr_399_wire_constant <= "00000000";
    array_obj_ref_318_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_318_gather_scatter_ack_0 <= array_obj_ref_318_gather_scatter_req_0;
      aggregated_sig <= expr_319_wire_constant;
      array_obj_ref_318_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_322_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_322_gather_scatter_ack_0 <= array_obj_ref_322_gather_scatter_req_0;
      aggregated_sig <= expr_323_wire_constant;
      array_obj_ref_322_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_326_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_326_gather_scatter_ack_0 <= array_obj_ref_326_gather_scatter_req_0;
      aggregated_sig <= expr_327_wire_constant;
      array_obj_ref_326_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_330_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_330_gather_scatter_ack_0 <= array_obj_ref_330_gather_scatter_req_0;
      aggregated_sig <= expr_331_wire_constant;
      array_obj_ref_330_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_334_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_334_gather_scatter_ack_0 <= array_obj_ref_334_gather_scatter_req_0;
      aggregated_sig <= expr_335_wire_constant;
      array_obj_ref_334_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_338_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_338_gather_scatter_ack_0 <= array_obj_ref_338_gather_scatter_req_0;
      aggregated_sig <= expr_339_wire_constant;
      array_obj_ref_338_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_342_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_342_gather_scatter_ack_0 <= array_obj_ref_342_gather_scatter_req_0;
      aggregated_sig <= expr_343_wire_constant;
      array_obj_ref_342_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_346_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_346_gather_scatter_ack_0 <= array_obj_ref_346_gather_scatter_req_0;
      aggregated_sig <= expr_347_wire_constant;
      array_obj_ref_346_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_350_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_350_gather_scatter_ack_0 <= array_obj_ref_350_gather_scatter_req_0;
      aggregated_sig <= expr_351_wire_constant;
      array_obj_ref_350_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_354_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_354_gather_scatter_ack_0 <= array_obj_ref_354_gather_scatter_req_0;
      aggregated_sig <= expr_355_wire_constant;
      array_obj_ref_354_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_358_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_358_gather_scatter_ack_0 <= array_obj_ref_358_gather_scatter_req_0;
      aggregated_sig <= expr_359_wire_constant;
      array_obj_ref_358_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_362_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_362_gather_scatter_ack_0 <= array_obj_ref_362_gather_scatter_req_0;
      aggregated_sig <= expr_363_wire_constant;
      array_obj_ref_362_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_366_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_366_gather_scatter_ack_0 <= array_obj_ref_366_gather_scatter_req_0;
      aggregated_sig <= expr_367_wire_constant;
      array_obj_ref_366_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_370_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_370_gather_scatter_ack_0 <= array_obj_ref_370_gather_scatter_req_0;
      aggregated_sig <= expr_371_wire_constant;
      array_obj_ref_370_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_374_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_374_gather_scatter_ack_0 <= array_obj_ref_374_gather_scatter_req_0;
      aggregated_sig <= expr_375_wire_constant;
      array_obj_ref_374_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_378_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_378_gather_scatter_ack_0 <= array_obj_ref_378_gather_scatter_req_0;
      aggregated_sig <= expr_379_wire_constant;
      array_obj_ref_378_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_382_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_382_gather_scatter_ack_0 <= array_obj_ref_382_gather_scatter_req_0;
      aggregated_sig <= expr_383_wire_constant;
      array_obj_ref_382_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_386_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_386_gather_scatter_ack_0 <= array_obj_ref_386_gather_scatter_req_0;
      aggregated_sig <= expr_387_wire_constant;
      array_obj_ref_386_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_390_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_390_gather_scatter_ack_0 <= array_obj_ref_390_gather_scatter_req_0;
      aggregated_sig <= expr_391_wire_constant;
      array_obj_ref_390_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_394_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_394_gather_scatter_ack_0 <= array_obj_ref_394_gather_scatter_req_0;
      aggregated_sig <= expr_395_wire_constant;
      array_obj_ref_394_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_398_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_398_gather_scatter_ack_0 <= array_obj_ref_398_gather_scatter_req_0;
      aggregated_sig <= expr_399_wire_constant;
      array_obj_ref_398_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_338_store_0 array_obj_ref_386_store_0 array_obj_ref_342_store_0 array_obj_ref_398_store_0 array_obj_ref_374_store_0 array_obj_ref_382_store_0 array_obj_ref_390_store_0 array_obj_ref_326_store_0 array_obj_ref_318_store_0 array_obj_ref_394_store_0 array_obj_ref_370_store_0 array_obj_ref_322_store_0 array_obj_ref_346_store_0 array_obj_ref_330_store_0 array_obj_ref_350_store_0 array_obj_ref_334_store_0 array_obj_ref_354_store_0 array_obj_ref_378_store_0 array_obj_ref_358_store_0 array_obj_ref_362_store_0 array_obj_ref_366_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(104 downto 0);
      signal data_in: std_logic_vector(167 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 20 downto 0);
      -- 
    begin -- 
      reqL(20) <= array_obj_ref_338_store_0_req_0;
      reqL(19) <= array_obj_ref_386_store_0_req_0;
      reqL(18) <= array_obj_ref_342_store_0_req_0;
      reqL(17) <= array_obj_ref_398_store_0_req_0;
      reqL(16) <= array_obj_ref_374_store_0_req_0;
      reqL(15) <= array_obj_ref_382_store_0_req_0;
      reqL(14) <= array_obj_ref_390_store_0_req_0;
      reqL(13) <= array_obj_ref_326_store_0_req_0;
      reqL(12) <= array_obj_ref_318_store_0_req_0;
      reqL(11) <= array_obj_ref_394_store_0_req_0;
      reqL(10) <= array_obj_ref_370_store_0_req_0;
      reqL(9) <= array_obj_ref_322_store_0_req_0;
      reqL(8) <= array_obj_ref_346_store_0_req_0;
      reqL(7) <= array_obj_ref_330_store_0_req_0;
      reqL(6) <= array_obj_ref_350_store_0_req_0;
      reqL(5) <= array_obj_ref_334_store_0_req_0;
      reqL(4) <= array_obj_ref_354_store_0_req_0;
      reqL(3) <= array_obj_ref_378_store_0_req_0;
      reqL(2) <= array_obj_ref_358_store_0_req_0;
      reqL(1) <= array_obj_ref_362_store_0_req_0;
      reqL(0) <= array_obj_ref_366_store_0_req_0;
      array_obj_ref_338_store_0_ack_0 <= ackL(20);
      array_obj_ref_386_store_0_ack_0 <= ackL(19);
      array_obj_ref_342_store_0_ack_0 <= ackL(18);
      array_obj_ref_398_store_0_ack_0 <= ackL(17);
      array_obj_ref_374_store_0_ack_0 <= ackL(16);
      array_obj_ref_382_store_0_ack_0 <= ackL(15);
      array_obj_ref_390_store_0_ack_0 <= ackL(14);
      array_obj_ref_326_store_0_ack_0 <= ackL(13);
      array_obj_ref_318_store_0_ack_0 <= ackL(12);
      array_obj_ref_394_store_0_ack_0 <= ackL(11);
      array_obj_ref_370_store_0_ack_0 <= ackL(10);
      array_obj_ref_322_store_0_ack_0 <= ackL(9);
      array_obj_ref_346_store_0_ack_0 <= ackL(8);
      array_obj_ref_330_store_0_ack_0 <= ackL(7);
      array_obj_ref_350_store_0_ack_0 <= ackL(6);
      array_obj_ref_334_store_0_ack_0 <= ackL(5);
      array_obj_ref_354_store_0_ack_0 <= ackL(4);
      array_obj_ref_378_store_0_ack_0 <= ackL(3);
      array_obj_ref_358_store_0_ack_0 <= ackL(2);
      array_obj_ref_362_store_0_ack_0 <= ackL(1);
      array_obj_ref_366_store_0_ack_0 <= ackL(0);
      reqR(20) <= array_obj_ref_338_store_0_req_1;
      reqR(19) <= array_obj_ref_386_store_0_req_1;
      reqR(18) <= array_obj_ref_342_store_0_req_1;
      reqR(17) <= array_obj_ref_398_store_0_req_1;
      reqR(16) <= array_obj_ref_374_store_0_req_1;
      reqR(15) <= array_obj_ref_382_store_0_req_1;
      reqR(14) <= array_obj_ref_390_store_0_req_1;
      reqR(13) <= array_obj_ref_326_store_0_req_1;
      reqR(12) <= array_obj_ref_318_store_0_req_1;
      reqR(11) <= array_obj_ref_394_store_0_req_1;
      reqR(10) <= array_obj_ref_370_store_0_req_1;
      reqR(9) <= array_obj_ref_322_store_0_req_1;
      reqR(8) <= array_obj_ref_346_store_0_req_1;
      reqR(7) <= array_obj_ref_330_store_0_req_1;
      reqR(6) <= array_obj_ref_350_store_0_req_1;
      reqR(5) <= array_obj_ref_334_store_0_req_1;
      reqR(4) <= array_obj_ref_354_store_0_req_1;
      reqR(3) <= array_obj_ref_378_store_0_req_1;
      reqR(2) <= array_obj_ref_358_store_0_req_1;
      reqR(1) <= array_obj_ref_362_store_0_req_1;
      reqR(0) <= array_obj_ref_366_store_0_req_1;
      array_obj_ref_338_store_0_ack_1 <= ackR(20);
      array_obj_ref_386_store_0_ack_1 <= ackR(19);
      array_obj_ref_342_store_0_ack_1 <= ackR(18);
      array_obj_ref_398_store_0_ack_1 <= ackR(17);
      array_obj_ref_374_store_0_ack_1 <= ackR(16);
      array_obj_ref_382_store_0_ack_1 <= ackR(15);
      array_obj_ref_390_store_0_ack_1 <= ackR(14);
      array_obj_ref_326_store_0_ack_1 <= ackR(13);
      array_obj_ref_318_store_0_ack_1 <= ackR(12);
      array_obj_ref_394_store_0_ack_1 <= ackR(11);
      array_obj_ref_370_store_0_ack_1 <= ackR(10);
      array_obj_ref_322_store_0_ack_1 <= ackR(9);
      array_obj_ref_346_store_0_ack_1 <= ackR(8);
      array_obj_ref_330_store_0_ack_1 <= ackR(7);
      array_obj_ref_350_store_0_ack_1 <= ackR(6);
      array_obj_ref_334_store_0_ack_1 <= ackR(5);
      array_obj_ref_354_store_0_ack_1 <= ackR(4);
      array_obj_ref_378_store_0_ack_1 <= ackR(3);
      array_obj_ref_358_store_0_ack_1 <= ackR(2);
      array_obj_ref_362_store_0_ack_1 <= ackR(1);
      array_obj_ref_366_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_338_word_address_0 & array_obj_ref_386_word_address_0 & array_obj_ref_342_word_address_0 & array_obj_ref_398_word_address_0 & array_obj_ref_374_word_address_0 & array_obj_ref_382_word_address_0 & array_obj_ref_390_word_address_0 & array_obj_ref_326_word_address_0 & array_obj_ref_318_word_address_0 & array_obj_ref_394_word_address_0 & array_obj_ref_370_word_address_0 & array_obj_ref_322_word_address_0 & array_obj_ref_346_word_address_0 & array_obj_ref_330_word_address_0 & array_obj_ref_350_word_address_0 & array_obj_ref_334_word_address_0 & array_obj_ref_354_word_address_0 & array_obj_ref_378_word_address_0 & array_obj_ref_358_word_address_0 & array_obj_ref_362_word_address_0 & array_obj_ref_366_word_address_0;
      data_in <= array_obj_ref_338_data_0 & array_obj_ref_386_data_0 & array_obj_ref_342_data_0 & array_obj_ref_398_data_0 & array_obj_ref_374_data_0 & array_obj_ref_382_data_0 & array_obj_ref_390_data_0 & array_obj_ref_326_data_0 & array_obj_ref_318_data_0 & array_obj_ref_394_data_0 & array_obj_ref_370_data_0 & array_obj_ref_322_data_0 & array_obj_ref_346_data_0 & array_obj_ref_330_data_0 & array_obj_ref_350_data_0 & array_obj_ref_334_data_0 & array_obj_ref_354_data_0 & array_obj_ref_378_data_0 & array_obj_ref_358_data_0 & array_obj_ref_362_data_0 & array_obj_ref_366_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 8,
        num_reqs => 21,
        tag_length => 5,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(4 downto 0),
          mdata => memory_space_6_sr_data(7 downto 0),
          mtag => memory_space_6_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 21,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr11 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr11;
architecture Default of default_initializer_xx_xstr11 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr11_CP_1629_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_404_gather_scatter_req_0 : boolean;
  signal array_obj_ref_404_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_404_store_0_req_0 : boolean;
  signal array_obj_ref_404_store_0_ack_0 : boolean;
  signal array_obj_ref_404_store_0_req_1 : boolean;
  signal array_obj_ref_404_store_0_ack_1 : boolean;
  signal array_obj_ref_408_gather_scatter_req_0 : boolean;
  signal array_obj_ref_408_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_408_store_0_req_0 : boolean;
  signal array_obj_ref_408_store_0_ack_0 : boolean;
  signal array_obj_ref_408_store_0_req_1 : boolean;
  signal array_obj_ref_408_store_0_ack_1 : boolean;
  signal array_obj_ref_412_gather_scatter_req_0 : boolean;
  signal array_obj_ref_412_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_412_store_0_req_0 : boolean;
  signal array_obj_ref_412_store_0_ack_0 : boolean;
  signal array_obj_ref_412_store_0_req_1 : boolean;
  signal array_obj_ref_412_store_0_ack_1 : boolean;
  signal array_obj_ref_416_gather_scatter_req_0 : boolean;
  signal array_obj_ref_416_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_416_store_0_req_0 : boolean;
  signal array_obj_ref_416_store_0_ack_0 : boolean;
  signal array_obj_ref_416_store_0_req_1 : boolean;
  signal array_obj_ref_416_store_0_ack_1 : boolean;
  signal array_obj_ref_420_gather_scatter_req_0 : boolean;
  signal array_obj_ref_420_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_420_store_0_req_0 : boolean;
  signal array_obj_ref_420_store_0_ack_0 : boolean;
  signal array_obj_ref_420_store_0_req_1 : boolean;
  signal array_obj_ref_420_store_0_ack_1 : boolean;
  signal array_obj_ref_424_gather_scatter_req_0 : boolean;
  signal array_obj_ref_424_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_424_store_0_req_0 : boolean;
  signal array_obj_ref_424_store_0_ack_0 : boolean;
  signal array_obj_ref_424_store_0_req_1 : boolean;
  signal array_obj_ref_424_store_0_ack_1 : boolean;
  signal array_obj_ref_428_gather_scatter_req_0 : boolean;
  signal array_obj_ref_428_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_428_store_0_req_0 : boolean;
  signal array_obj_ref_428_store_0_ack_0 : boolean;
  signal array_obj_ref_428_store_0_req_1 : boolean;
  signal array_obj_ref_428_store_0_ack_1 : boolean;
  signal array_obj_ref_432_gather_scatter_req_0 : boolean;
  signal array_obj_ref_432_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_432_store_0_req_0 : boolean;
  signal array_obj_ref_432_store_0_ack_0 : boolean;
  signal array_obj_ref_432_store_0_req_1 : boolean;
  signal array_obj_ref_432_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 8 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr11_CP_1629: Block -- control-path 
    signal cp_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(24);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(24), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_404_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_404_gather_scatter_ack_0;
    array_obj_ref_404_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_404_store_0_ack_0;
    array_obj_ref_404_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_404_store_0_ack_1;
    array_obj_ref_408_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_408_gather_scatter_ack_0;
    array_obj_ref_408_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_408_store_0_ack_0;
    array_obj_ref_408_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_408_store_0_ack_1;
    array_obj_ref_412_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_412_gather_scatter_ack_0;
    array_obj_ref_412_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_412_store_0_ack_0;
    array_obj_ref_412_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_412_store_0_ack_1;
    array_obj_ref_416_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_416_gather_scatter_ack_0;
    array_obj_ref_416_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_416_store_0_ack_0;
    array_obj_ref_416_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_416_store_0_ack_1;
    array_obj_ref_420_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_420_gather_scatter_ack_0;
    array_obj_ref_420_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_420_store_0_ack_0;
    array_obj_ref_420_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_420_store_0_ack_1;
    array_obj_ref_424_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_424_gather_scatter_ack_0;
    array_obj_ref_424_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_424_store_0_ack_0;
    array_obj_ref_424_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_424_store_0_ack_1;
    array_obj_ref_428_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_428_gather_scatter_ack_0;
    array_obj_ref_428_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_428_store_0_ack_0;
    array_obj_ref_428_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_428_store_0_ack_1;
    array_obj_ref_432_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_432_gather_scatter_ack_0;
    array_obj_ref_432_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_432_store_0_ack_0;
    array_obj_ref_432_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_432_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_404_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_404_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_408_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_408_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_412_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_412_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_416_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_416_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_420_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_420_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_424_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_424_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_428_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_428_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_432_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_432_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_405_wire_constant : std_logic_vector(7 downto 0);
    signal expr_409_wire_constant : std_logic_vector(7 downto 0);
    signal expr_413_wire_constant : std_logic_vector(7 downto 0);
    signal expr_417_wire_constant : std_logic_vector(7 downto 0);
    signal expr_421_wire_constant : std_logic_vector(7 downto 0);
    signal expr_425_wire_constant : std_logic_vector(7 downto 0);
    signal expr_429_wire_constant : std_logic_vector(7 downto 0);
    signal expr_433_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_404_word_address_0 <= "0000";
    array_obj_ref_408_word_address_0 <= "0001";
    array_obj_ref_412_word_address_0 <= "0010";
    array_obj_ref_416_word_address_0 <= "0011";
    array_obj_ref_420_word_address_0 <= "0100";
    array_obj_ref_424_word_address_0 <= "0101";
    array_obj_ref_428_word_address_0 <= "0110";
    array_obj_ref_432_word_address_0 <= "0111";
    expr_405_wire_constant <= "01101001";
    expr_409_wire_constant <= "01101110";
    expr_413_wire_constant <= "01011111";
    expr_417_wire_constant <= "01100100";
    expr_421_wire_constant <= "01100001";
    expr_425_wire_constant <= "01110100";
    expr_429_wire_constant <= "01100001";
    expr_433_wire_constant <= "00000000";
    array_obj_ref_404_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_404_gather_scatter_ack_0 <= array_obj_ref_404_gather_scatter_req_0;
      aggregated_sig <= expr_405_wire_constant;
      array_obj_ref_404_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_408_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_408_gather_scatter_ack_0 <= array_obj_ref_408_gather_scatter_req_0;
      aggregated_sig <= expr_409_wire_constant;
      array_obj_ref_408_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_412_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_412_gather_scatter_ack_0 <= array_obj_ref_412_gather_scatter_req_0;
      aggregated_sig <= expr_413_wire_constant;
      array_obj_ref_412_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_416_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_416_gather_scatter_ack_0 <= array_obj_ref_416_gather_scatter_req_0;
      aggregated_sig <= expr_417_wire_constant;
      array_obj_ref_416_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_420_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_420_gather_scatter_ack_0 <= array_obj_ref_420_gather_scatter_req_0;
      aggregated_sig <= expr_421_wire_constant;
      array_obj_ref_420_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_424_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_424_gather_scatter_ack_0 <= array_obj_ref_424_gather_scatter_req_0;
      aggregated_sig <= expr_425_wire_constant;
      array_obj_ref_424_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_428_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_428_gather_scatter_ack_0 <= array_obj_ref_428_gather_scatter_req_0;
      aggregated_sig <= expr_429_wire_constant;
      array_obj_ref_428_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_432_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_432_gather_scatter_ack_0 <= array_obj_ref_432_gather_scatter_req_0;
      aggregated_sig <= expr_433_wire_constant;
      array_obj_ref_432_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_404_store_0 array_obj_ref_408_store_0 array_obj_ref_412_store_0 array_obj_ref_416_store_0 array_obj_ref_420_store_0 array_obj_ref_424_store_0 array_obj_ref_428_store_0 array_obj_ref_432_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= array_obj_ref_404_store_0_req_0;
      reqL(6) <= array_obj_ref_408_store_0_req_0;
      reqL(5) <= array_obj_ref_412_store_0_req_0;
      reqL(4) <= array_obj_ref_416_store_0_req_0;
      reqL(3) <= array_obj_ref_420_store_0_req_0;
      reqL(2) <= array_obj_ref_424_store_0_req_0;
      reqL(1) <= array_obj_ref_428_store_0_req_0;
      reqL(0) <= array_obj_ref_432_store_0_req_0;
      array_obj_ref_404_store_0_ack_0 <= ackL(7);
      array_obj_ref_408_store_0_ack_0 <= ackL(6);
      array_obj_ref_412_store_0_ack_0 <= ackL(5);
      array_obj_ref_416_store_0_ack_0 <= ackL(4);
      array_obj_ref_420_store_0_ack_0 <= ackL(3);
      array_obj_ref_424_store_0_ack_0 <= ackL(2);
      array_obj_ref_428_store_0_ack_0 <= ackL(1);
      array_obj_ref_432_store_0_ack_0 <= ackL(0);
      reqR(7) <= array_obj_ref_404_store_0_req_1;
      reqR(6) <= array_obj_ref_408_store_0_req_1;
      reqR(5) <= array_obj_ref_412_store_0_req_1;
      reqR(4) <= array_obj_ref_416_store_0_req_1;
      reqR(3) <= array_obj_ref_420_store_0_req_1;
      reqR(2) <= array_obj_ref_424_store_0_req_1;
      reqR(1) <= array_obj_ref_428_store_0_req_1;
      reqR(0) <= array_obj_ref_432_store_0_req_1;
      array_obj_ref_404_store_0_ack_1 <= ackR(7);
      array_obj_ref_408_store_0_ack_1 <= ackR(6);
      array_obj_ref_412_store_0_ack_1 <= ackR(5);
      array_obj_ref_416_store_0_ack_1 <= ackR(4);
      array_obj_ref_420_store_0_ack_1 <= ackR(3);
      array_obj_ref_424_store_0_ack_1 <= ackR(2);
      array_obj_ref_428_store_0_ack_1 <= ackR(1);
      array_obj_ref_432_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_404_word_address_0 & array_obj_ref_408_word_address_0 & array_obj_ref_412_word_address_0 & array_obj_ref_416_word_address_0 & array_obj_ref_420_word_address_0 & array_obj_ref_424_word_address_0 & array_obj_ref_428_word_address_0 & array_obj_ref_432_word_address_0;
      data_in <= array_obj_ref_404_data_0 & array_obj_ref_408_data_0 & array_obj_ref_412_data_0 & array_obj_ref_416_data_0 & array_obj_ref_420_data_0 & array_obj_ref_424_data_0 & array_obj_ref_428_data_0 & array_obj_ref_432_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(3 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr12 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr12;
architecture Default of default_initializer_xx_xstr12 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr12_CP_1800_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_442_store_0_ack_1 : boolean;
  signal array_obj_ref_438_store_0_ack_1 : boolean;
  signal array_obj_ref_466_store_0_ack_1 : boolean;
  signal array_obj_ref_442_gather_scatter_req_0 : boolean;
  signal array_obj_ref_462_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_0 : boolean;
  signal array_obj_ref_450_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_454_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_446_gather_scatter_req_0 : boolean;
  signal array_obj_ref_458_gather_scatter_req_0 : boolean;
  signal array_obj_ref_458_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_450_gather_scatter_req_0 : boolean;
  signal array_obj_ref_466_gather_scatter_req_0 : boolean;
  signal array_obj_ref_466_store_0_req_1 : boolean;
  signal array_obj_ref_466_store_0_ack_0 : boolean;
  signal array_obj_ref_454_store_0_ack_0 : boolean;
  signal array_obj_ref_450_store_0_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_0 : boolean;
  signal array_obj_ref_438_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_450_store_0_ack_1 : boolean;
  signal array_obj_ref_450_store_0_req_0 : boolean;
  signal array_obj_ref_446_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_446_store_0_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_0 : boolean;
  signal array_obj_ref_446_store_0_ack_1 : boolean;
  signal array_obj_ref_438_store_0_ack_0 : boolean;
  signal array_obj_ref_450_store_0_req_1 : boolean;
  signal array_obj_ref_454_store_0_req_0 : boolean;
  signal array_obj_ref_446_store_0_req_1 : boolean;
  signal array_obj_ref_442_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_438_gather_scatter_req_0 : boolean;
  signal array_obj_ref_446_store_0_req_0 : boolean;
  signal array_obj_ref_462_gather_scatter_req_0 : boolean;
  signal array_obj_ref_454_store_0_req_1 : boolean;
  signal array_obj_ref_466_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_1 : boolean;
  signal array_obj_ref_458_store_0_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_1 : boolean;
  signal array_obj_ref_458_store_0_ack_1 : boolean;
  signal array_obj_ref_442_store_0_req_0 : boolean;
  signal array_obj_ref_442_store_0_ack_0 : boolean;
  signal array_obj_ref_442_store_0_req_1 : boolean;
  signal array_obj_ref_454_gather_scatter_req_0 : boolean;
  signal array_obj_ref_462_store_0_ack_1 : boolean;
  signal array_obj_ref_462_store_0_req_1 : boolean;
  signal array_obj_ref_462_store_0_ack_0 : boolean;
  signal array_obj_ref_462_store_0_req_0 : boolean;
  signal array_obj_ref_454_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 8 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr12_CP_1800: Block -- control-path 
    signal cp_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(24);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(24), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_438_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_438_gather_scatter_ack_0;
    array_obj_ref_438_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_438_store_0_ack_0;
    array_obj_ref_438_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_438_store_0_ack_1;
    array_obj_ref_442_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_442_gather_scatter_ack_0;
    array_obj_ref_442_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_442_store_0_ack_0;
    array_obj_ref_442_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_442_store_0_ack_1;
    array_obj_ref_446_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_446_gather_scatter_ack_0;
    array_obj_ref_446_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_446_store_0_ack_0;
    array_obj_ref_446_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_446_store_0_ack_1;
    array_obj_ref_450_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_450_gather_scatter_ack_0;
    array_obj_ref_450_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_450_store_0_ack_0;
    array_obj_ref_450_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_450_store_0_ack_1;
    array_obj_ref_454_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_454_gather_scatter_ack_0;
    array_obj_ref_454_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_454_store_0_ack_0;
    array_obj_ref_454_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_454_store_0_ack_1;
    array_obj_ref_458_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_458_gather_scatter_ack_0;
    array_obj_ref_458_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_458_store_0_ack_0;
    array_obj_ref_458_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_458_store_0_ack_1;
    array_obj_ref_462_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_462_gather_scatter_ack_0;
    array_obj_ref_462_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_462_store_0_ack_0;
    array_obj_ref_462_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_462_store_0_ack_1;
    array_obj_ref_466_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_466_gather_scatter_ack_0;
    array_obj_ref_466_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_466_store_0_ack_0;
    array_obj_ref_466_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_466_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_438_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_442_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_442_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_446_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_446_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_450_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_454_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_454_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_458_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_458_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_462_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_466_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_466_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_439_wire_constant : std_logic_vector(7 downto 0);
    signal expr_443_wire_constant : std_logic_vector(7 downto 0);
    signal expr_447_wire_constant : std_logic_vector(7 downto 0);
    signal expr_451_wire_constant : std_logic_vector(7 downto 0);
    signal expr_455_wire_constant : std_logic_vector(7 downto 0);
    signal expr_459_wire_constant : std_logic_vector(7 downto 0);
    signal expr_463_wire_constant : std_logic_vector(7 downto 0);
    signal expr_467_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_438_word_address_0 <= "0000";
    array_obj_ref_442_word_address_0 <= "0001";
    array_obj_ref_446_word_address_0 <= "0010";
    array_obj_ref_450_word_address_0 <= "0011";
    array_obj_ref_454_word_address_0 <= "0100";
    array_obj_ref_458_word_address_0 <= "0101";
    array_obj_ref_462_word_address_0 <= "0110";
    array_obj_ref_466_word_address_0 <= "0111";
    expr_439_wire_constant <= "01101001";
    expr_443_wire_constant <= "01101110";
    expr_447_wire_constant <= "01011111";
    expr_451_wire_constant <= "01100011";
    expr_455_wire_constant <= "01110100";
    expr_459_wire_constant <= "01110010";
    expr_463_wire_constant <= "01101100";
    expr_467_wire_constant <= "00000000";
    array_obj_ref_438_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_438_gather_scatter_ack_0 <= array_obj_ref_438_gather_scatter_req_0;
      aggregated_sig <= expr_439_wire_constant;
      array_obj_ref_438_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_442_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_442_gather_scatter_ack_0 <= array_obj_ref_442_gather_scatter_req_0;
      aggregated_sig <= expr_443_wire_constant;
      array_obj_ref_442_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_446_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_446_gather_scatter_ack_0 <= array_obj_ref_446_gather_scatter_req_0;
      aggregated_sig <= expr_447_wire_constant;
      array_obj_ref_446_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_450_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_450_gather_scatter_ack_0 <= array_obj_ref_450_gather_scatter_req_0;
      aggregated_sig <= expr_451_wire_constant;
      array_obj_ref_450_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_454_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_454_gather_scatter_ack_0 <= array_obj_ref_454_gather_scatter_req_0;
      aggregated_sig <= expr_455_wire_constant;
      array_obj_ref_454_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_458_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_458_gather_scatter_ack_0 <= array_obj_ref_458_gather_scatter_req_0;
      aggregated_sig <= expr_459_wire_constant;
      array_obj_ref_458_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_462_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_462_gather_scatter_ack_0 <= array_obj_ref_462_gather_scatter_req_0;
      aggregated_sig <= expr_463_wire_constant;
      array_obj_ref_462_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_466_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_466_gather_scatter_ack_0 <= array_obj_ref_466_gather_scatter_req_0;
      aggregated_sig <= expr_467_wire_constant;
      array_obj_ref_466_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_446_store_0 array_obj_ref_438_store_0 array_obj_ref_450_store_0 array_obj_ref_442_store_0 array_obj_ref_454_store_0 array_obj_ref_466_store_0 array_obj_ref_458_store_0 array_obj_ref_462_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= array_obj_ref_446_store_0_req_0;
      reqL(6) <= array_obj_ref_438_store_0_req_0;
      reqL(5) <= array_obj_ref_450_store_0_req_0;
      reqL(4) <= array_obj_ref_442_store_0_req_0;
      reqL(3) <= array_obj_ref_454_store_0_req_0;
      reqL(2) <= array_obj_ref_466_store_0_req_0;
      reqL(1) <= array_obj_ref_458_store_0_req_0;
      reqL(0) <= array_obj_ref_462_store_0_req_0;
      array_obj_ref_446_store_0_ack_0 <= ackL(7);
      array_obj_ref_438_store_0_ack_0 <= ackL(6);
      array_obj_ref_450_store_0_ack_0 <= ackL(5);
      array_obj_ref_442_store_0_ack_0 <= ackL(4);
      array_obj_ref_454_store_0_ack_0 <= ackL(3);
      array_obj_ref_466_store_0_ack_0 <= ackL(2);
      array_obj_ref_458_store_0_ack_0 <= ackL(1);
      array_obj_ref_462_store_0_ack_0 <= ackL(0);
      reqR(7) <= array_obj_ref_446_store_0_req_1;
      reqR(6) <= array_obj_ref_438_store_0_req_1;
      reqR(5) <= array_obj_ref_450_store_0_req_1;
      reqR(4) <= array_obj_ref_442_store_0_req_1;
      reqR(3) <= array_obj_ref_454_store_0_req_1;
      reqR(2) <= array_obj_ref_466_store_0_req_1;
      reqR(1) <= array_obj_ref_458_store_0_req_1;
      reqR(0) <= array_obj_ref_462_store_0_req_1;
      array_obj_ref_446_store_0_ack_1 <= ackR(7);
      array_obj_ref_438_store_0_ack_1 <= ackR(6);
      array_obj_ref_450_store_0_ack_1 <= ackR(5);
      array_obj_ref_442_store_0_ack_1 <= ackR(4);
      array_obj_ref_454_store_0_ack_1 <= ackR(3);
      array_obj_ref_466_store_0_ack_1 <= ackR(2);
      array_obj_ref_458_store_0_ack_1 <= ackR(1);
      array_obj_ref_462_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_446_word_address_0 & array_obj_ref_438_word_address_0 & array_obj_ref_450_word_address_0 & array_obj_ref_442_word_address_0 & array_obj_ref_454_word_address_0 & array_obj_ref_466_word_address_0 & array_obj_ref_458_word_address_0 & array_obj_ref_462_word_address_0;
      data_in <= array_obj_ref_446_data_0 & array_obj_ref_438_data_0 & array_obj_ref_450_data_0 & array_obj_ref_442_data_0 & array_obj_ref_454_data_0 & array_obj_ref_466_data_0 & array_obj_ref_458_data_0 & array_obj_ref_462_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(3 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr13 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_9_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr13;
architecture Default of default_initializer_xx_xstr13 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr13_CP_1971_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_476_store_0_ack_1 : boolean;
  signal array_obj_ref_480_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_484_store_0_ack_0 : boolean;
  signal array_obj_ref_480_store_0_ack_0 : boolean;
  signal array_obj_ref_500_store_0_ack_1 : boolean;
  signal array_obj_ref_484_store_0_req_0 : boolean;
  signal array_obj_ref_496_gather_scatter_req_0 : boolean;
  signal array_obj_ref_480_store_0_req_1 : boolean;
  signal array_obj_ref_488_store_0_ack_1 : boolean;
  signal array_obj_ref_484_gather_scatter_req_0 : boolean;
  signal array_obj_ref_476_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_472_store_0_req_0 : boolean;
  signal array_obj_ref_500_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_500_gather_scatter_req_0 : boolean;
  signal array_obj_ref_472_store_0_req_1 : boolean;
  signal array_obj_ref_492_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_488_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_492_store_0_req_0 : boolean;
  signal array_obj_ref_476_store_0_req_0 : boolean;
  signal array_obj_ref_500_store_0_req_1 : boolean;
  signal array_obj_ref_484_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_496_store_0_ack_1 : boolean;
  signal array_obj_ref_496_store_0_req_1 : boolean;
  signal array_obj_ref_488_store_0_ack_0 : boolean;
  signal array_obj_ref_472_store_0_ack_0 : boolean;
  signal array_obj_ref_488_gather_scatter_req_0 : boolean;
  signal array_obj_ref_480_store_0_req_0 : boolean;
  signal array_obj_ref_472_store_0_ack_1 : boolean;
  signal array_obj_ref_480_store_0_ack_1 : boolean;
  signal array_obj_ref_492_store_0_req_1 : boolean;
  signal array_obj_ref_492_gather_scatter_req_0 : boolean;
  signal array_obj_ref_500_store_0_req_0 : boolean;
  signal array_obj_ref_476_store_0_req_1 : boolean;
  signal array_obj_ref_496_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_476_store_0_ack_0 : boolean;
  signal array_obj_ref_500_store_0_ack_0 : boolean;
  signal array_obj_ref_480_gather_scatter_req_0 : boolean;
  signal array_obj_ref_488_store_0_req_0 : boolean;
  signal array_obj_ref_476_gather_scatter_req_0 : boolean;
  signal array_obj_ref_492_store_0_ack_1 : boolean;
  signal array_obj_ref_492_store_0_ack_0 : boolean;
  signal array_obj_ref_496_store_0_req_0 : boolean;
  signal array_obj_ref_484_store_0_ack_1 : boolean;
  signal array_obj_ref_472_gather_scatter_req_0 : boolean;
  signal array_obj_ref_472_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_496_store_0_ack_0 : boolean;
  signal array_obj_ref_488_store_0_req_1 : boolean;
  signal array_obj_ref_484_store_0_req_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 8 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr13_CP_1971: Block -- control-path 
    signal cp_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(24);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(24), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_472_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_472_gather_scatter_ack_0;
    array_obj_ref_472_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_472_store_0_ack_0;
    array_obj_ref_472_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_472_store_0_ack_1;
    array_obj_ref_476_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_476_gather_scatter_ack_0;
    array_obj_ref_476_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_476_store_0_ack_0;
    array_obj_ref_476_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_476_store_0_ack_1;
    array_obj_ref_480_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_480_gather_scatter_ack_0;
    array_obj_ref_480_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_480_store_0_ack_0;
    array_obj_ref_480_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_480_store_0_ack_1;
    array_obj_ref_484_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_484_gather_scatter_ack_0;
    array_obj_ref_484_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_484_store_0_ack_0;
    array_obj_ref_484_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_484_store_0_ack_1;
    array_obj_ref_488_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_488_gather_scatter_ack_0;
    array_obj_ref_488_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_488_store_0_ack_0;
    array_obj_ref_488_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_488_store_0_ack_1;
    array_obj_ref_492_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_492_gather_scatter_ack_0;
    array_obj_ref_492_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_492_store_0_ack_0;
    array_obj_ref_492_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_492_store_0_ack_1;
    array_obj_ref_496_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_496_gather_scatter_ack_0;
    array_obj_ref_496_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_496_store_0_ack_0;
    array_obj_ref_496_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_496_store_0_ack_1;
    array_obj_ref_500_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_500_gather_scatter_ack_0;
    array_obj_ref_500_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_500_store_0_ack_0;
    array_obj_ref_500_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_500_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_472_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_472_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_476_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_476_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_480_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_480_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_484_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_484_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_488_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_488_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_492_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_492_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_496_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_496_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_500_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_500_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_473_wire_constant : std_logic_vector(7 downto 0);
    signal expr_477_wire_constant : std_logic_vector(7 downto 0);
    signal expr_481_wire_constant : std_logic_vector(7 downto 0);
    signal expr_485_wire_constant : std_logic_vector(7 downto 0);
    signal expr_489_wire_constant : std_logic_vector(7 downto 0);
    signal expr_493_wire_constant : std_logic_vector(7 downto 0);
    signal expr_497_wire_constant : std_logic_vector(7 downto 0);
    signal expr_501_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_472_word_address_0 <= "0000";
    array_obj_ref_476_word_address_0 <= "0001";
    array_obj_ref_480_word_address_0 <= "0010";
    array_obj_ref_484_word_address_0 <= "0011";
    array_obj_ref_488_word_address_0 <= "0100";
    array_obj_ref_492_word_address_0 <= "0101";
    array_obj_ref_496_word_address_0 <= "0110";
    array_obj_ref_500_word_address_0 <= "0111";
    expr_473_wire_constant <= "01101101";
    expr_477_wire_constant <= "01101001";
    expr_481_wire_constant <= "01100100";
    expr_485_wire_constant <= "01110000";
    expr_489_wire_constant <= "01101001";
    expr_493_wire_constant <= "01110000";
    expr_497_wire_constant <= "01100101";
    expr_501_wire_constant <= "00000000";
    array_obj_ref_472_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_472_gather_scatter_ack_0 <= array_obj_ref_472_gather_scatter_req_0;
      aggregated_sig <= expr_473_wire_constant;
      array_obj_ref_472_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_476_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_476_gather_scatter_ack_0 <= array_obj_ref_476_gather_scatter_req_0;
      aggregated_sig <= expr_477_wire_constant;
      array_obj_ref_476_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_480_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_480_gather_scatter_ack_0 <= array_obj_ref_480_gather_scatter_req_0;
      aggregated_sig <= expr_481_wire_constant;
      array_obj_ref_480_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_484_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_484_gather_scatter_ack_0 <= array_obj_ref_484_gather_scatter_req_0;
      aggregated_sig <= expr_485_wire_constant;
      array_obj_ref_484_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_488_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_488_gather_scatter_ack_0 <= array_obj_ref_488_gather_scatter_req_0;
      aggregated_sig <= expr_489_wire_constant;
      array_obj_ref_488_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_492_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_492_gather_scatter_ack_0 <= array_obj_ref_492_gather_scatter_req_0;
      aggregated_sig <= expr_493_wire_constant;
      array_obj_ref_492_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_496_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_496_gather_scatter_ack_0 <= array_obj_ref_496_gather_scatter_req_0;
      aggregated_sig <= expr_497_wire_constant;
      array_obj_ref_496_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_500_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_500_gather_scatter_ack_0 <= array_obj_ref_500_gather_scatter_req_0;
      aggregated_sig <= expr_501_wire_constant;
      array_obj_ref_500_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_472_store_0 array_obj_ref_496_store_0 array_obj_ref_484_store_0 array_obj_ref_480_store_0 array_obj_ref_476_store_0 array_obj_ref_500_store_0 array_obj_ref_492_store_0 array_obj_ref_488_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= array_obj_ref_472_store_0_req_0;
      reqL(6) <= array_obj_ref_496_store_0_req_0;
      reqL(5) <= array_obj_ref_484_store_0_req_0;
      reqL(4) <= array_obj_ref_480_store_0_req_0;
      reqL(3) <= array_obj_ref_476_store_0_req_0;
      reqL(2) <= array_obj_ref_500_store_0_req_0;
      reqL(1) <= array_obj_ref_492_store_0_req_0;
      reqL(0) <= array_obj_ref_488_store_0_req_0;
      array_obj_ref_472_store_0_ack_0 <= ackL(7);
      array_obj_ref_496_store_0_ack_0 <= ackL(6);
      array_obj_ref_484_store_0_ack_0 <= ackL(5);
      array_obj_ref_480_store_0_ack_0 <= ackL(4);
      array_obj_ref_476_store_0_ack_0 <= ackL(3);
      array_obj_ref_500_store_0_ack_0 <= ackL(2);
      array_obj_ref_492_store_0_ack_0 <= ackL(1);
      array_obj_ref_488_store_0_ack_0 <= ackL(0);
      reqR(7) <= array_obj_ref_472_store_0_req_1;
      reqR(6) <= array_obj_ref_496_store_0_req_1;
      reqR(5) <= array_obj_ref_484_store_0_req_1;
      reqR(4) <= array_obj_ref_480_store_0_req_1;
      reqR(3) <= array_obj_ref_476_store_0_req_1;
      reqR(2) <= array_obj_ref_500_store_0_req_1;
      reqR(1) <= array_obj_ref_492_store_0_req_1;
      reqR(0) <= array_obj_ref_488_store_0_req_1;
      array_obj_ref_472_store_0_ack_1 <= ackR(7);
      array_obj_ref_496_store_0_ack_1 <= ackR(6);
      array_obj_ref_484_store_0_ack_1 <= ackR(5);
      array_obj_ref_480_store_0_ack_1 <= ackR(4);
      array_obj_ref_476_store_0_ack_1 <= ackR(3);
      array_obj_ref_500_store_0_ack_1 <= ackR(2);
      array_obj_ref_492_store_0_ack_1 <= ackR(1);
      array_obj_ref_488_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_472_word_address_0 & array_obj_ref_496_word_address_0 & array_obj_ref_484_word_address_0 & array_obj_ref_480_word_address_0 & array_obj_ref_476_word_address_0 & array_obj_ref_500_word_address_0 & array_obj_ref_492_word_address_0 & array_obj_ref_488_word_address_0;
      data_in <= array_obj_ref_472_data_0 & array_obj_ref_496_data_0 & array_obj_ref_484_data_0 & array_obj_ref_480_data_0 & array_obj_ref_476_data_0 & array_obj_ref_500_data_0 & array_obj_ref_492_data_0 & array_obj_ref_488_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(3 downto 0),
          mdata => memory_space_9_sr_data(7 downto 0),
          mtag => memory_space_9_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr14 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_10_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr14;
architecture Default of default_initializer_xx_xstr14 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr14_CP_2142_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_506_gather_scatter_req_0 : boolean;
  signal array_obj_ref_506_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_506_store_0_req_0 : boolean;
  signal array_obj_ref_506_store_0_ack_0 : boolean;
  signal array_obj_ref_506_store_0_req_1 : boolean;
  signal array_obj_ref_506_store_0_ack_1 : boolean;
  signal array_obj_ref_510_gather_scatter_req_0 : boolean;
  signal array_obj_ref_510_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_510_store_0_req_0 : boolean;
  signal array_obj_ref_510_store_0_ack_0 : boolean;
  signal array_obj_ref_510_store_0_req_1 : boolean;
  signal array_obj_ref_510_store_0_ack_1 : boolean;
  signal array_obj_ref_514_gather_scatter_req_0 : boolean;
  signal array_obj_ref_514_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_514_store_0_req_0 : boolean;
  signal array_obj_ref_514_store_0_ack_0 : boolean;
  signal array_obj_ref_514_store_0_req_1 : boolean;
  signal array_obj_ref_514_store_0_ack_1 : boolean;
  signal array_obj_ref_518_gather_scatter_req_0 : boolean;
  signal array_obj_ref_518_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_518_store_0_req_0 : boolean;
  signal array_obj_ref_518_store_0_ack_0 : boolean;
  signal array_obj_ref_518_store_0_req_1 : boolean;
  signal array_obj_ref_518_store_0_ack_1 : boolean;
  signal array_obj_ref_522_gather_scatter_req_0 : boolean;
  signal array_obj_ref_522_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_522_store_0_req_0 : boolean;
  signal array_obj_ref_522_store_0_ack_0 : boolean;
  signal array_obj_ref_522_store_0_req_1 : boolean;
  signal array_obj_ref_522_store_0_ack_1 : boolean;
  signal array_obj_ref_526_gather_scatter_req_0 : boolean;
  signal array_obj_ref_526_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_526_store_0_req_0 : boolean;
  signal array_obj_ref_526_store_0_ack_0 : boolean;
  signal array_obj_ref_526_store_0_req_1 : boolean;
  signal array_obj_ref_526_store_0_ack_1 : boolean;
  signal array_obj_ref_530_gather_scatter_req_0 : boolean;
  signal array_obj_ref_530_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_530_store_0_req_0 : boolean;
  signal array_obj_ref_530_store_0_ack_0 : boolean;
  signal array_obj_ref_530_store_0_req_1 : boolean;
  signal array_obj_ref_530_store_0_ack_1 : boolean;
  signal array_obj_ref_534_gather_scatter_req_0 : boolean;
  signal array_obj_ref_534_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_534_store_0_req_0 : boolean;
  signal array_obj_ref_534_store_0_ack_0 : boolean;
  signal array_obj_ref_534_store_0_req_1 : boolean;
  signal array_obj_ref_534_store_0_ack_1 : boolean;
  signal array_obj_ref_538_gather_scatter_req_0 : boolean;
  signal array_obj_ref_538_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_538_store_0_req_0 : boolean;
  signal array_obj_ref_538_store_0_ack_0 : boolean;
  signal array_obj_ref_538_store_0_req_1 : boolean;
  signal array_obj_ref_538_store_0_ack_1 : boolean;
  signal array_obj_ref_542_gather_scatter_req_0 : boolean;
  signal array_obj_ref_542_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_542_store_0_req_0 : boolean;
  signal array_obj_ref_542_store_0_ack_0 : boolean;
  signal array_obj_ref_542_store_0_req_1 : boolean;
  signal array_obj_ref_542_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 10 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr14_CP_2142: Block -- control-path 
    signal cp_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(30);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(30), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_506_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_506_gather_scatter_ack_0;
    array_obj_ref_506_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_506_store_0_ack_0;
    array_obj_ref_506_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_506_store_0_ack_1;
    array_obj_ref_510_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_510_gather_scatter_ack_0;
    array_obj_ref_510_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_510_store_0_ack_0;
    array_obj_ref_510_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_510_store_0_ack_1;
    array_obj_ref_514_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_514_gather_scatter_ack_0;
    array_obj_ref_514_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_514_store_0_ack_0;
    array_obj_ref_514_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_514_store_0_ack_1;
    array_obj_ref_518_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_518_gather_scatter_ack_0;
    array_obj_ref_518_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_518_store_0_ack_0;
    array_obj_ref_518_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_518_store_0_ack_1;
    array_obj_ref_522_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_522_gather_scatter_ack_0;
    array_obj_ref_522_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_522_store_0_ack_0;
    array_obj_ref_522_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_522_store_0_ack_1;
    array_obj_ref_526_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_526_gather_scatter_ack_0;
    array_obj_ref_526_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_526_store_0_ack_0;
    array_obj_ref_526_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_526_store_0_ack_1;
    array_obj_ref_530_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_530_gather_scatter_ack_0;
    array_obj_ref_530_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_530_store_0_ack_0;
    array_obj_ref_530_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_530_store_0_ack_1;
    array_obj_ref_534_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_534_gather_scatter_ack_0;
    array_obj_ref_534_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_534_store_0_ack_0;
    array_obj_ref_534_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_534_store_0_ack_1;
    array_obj_ref_538_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_538_gather_scatter_ack_0;
    array_obj_ref_538_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_538_store_0_ack_0;
    array_obj_ref_538_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_538_store_0_ack_1;
    array_obj_ref_542_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_542_gather_scatter_ack_0;
    array_obj_ref_542_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_542_store_0_ack_0;
    array_obj_ref_542_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_542_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_506_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_506_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_510_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_510_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_514_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_514_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_518_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_518_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_522_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_522_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_526_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_526_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_530_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_530_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_534_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_534_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_538_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_538_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_542_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_542_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_507_wire_constant : std_logic_vector(7 downto 0);
    signal expr_511_wire_constant : std_logic_vector(7 downto 0);
    signal expr_515_wire_constant : std_logic_vector(7 downto 0);
    signal expr_519_wire_constant : std_logic_vector(7 downto 0);
    signal expr_523_wire_constant : std_logic_vector(7 downto 0);
    signal expr_527_wire_constant : std_logic_vector(7 downto 0);
    signal expr_531_wire_constant : std_logic_vector(7 downto 0);
    signal expr_535_wire_constant : std_logic_vector(7 downto 0);
    signal expr_539_wire_constant : std_logic_vector(7 downto 0);
    signal expr_543_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_506_word_address_0 <= "0000";
    array_obj_ref_510_word_address_0 <= "0001";
    array_obj_ref_514_word_address_0 <= "0010";
    array_obj_ref_518_word_address_0 <= "0011";
    array_obj_ref_522_word_address_0 <= "0100";
    array_obj_ref_526_word_address_0 <= "0101";
    array_obj_ref_530_word_address_0 <= "0110";
    array_obj_ref_534_word_address_0 <= "0111";
    array_obj_ref_538_word_address_0 <= "1000";
    array_obj_ref_542_word_address_0 <= "1001";
    expr_507_wire_constant <= "01101100";
    expr_511_wire_constant <= "01100001";
    expr_515_wire_constant <= "01110011";
    expr_519_wire_constant <= "01110100";
    expr_523_wire_constant <= "01011111";
    expr_527_wire_constant <= "01100011";
    expr_531_wire_constant <= "01110100";
    expr_535_wire_constant <= "01110010";
    expr_539_wire_constant <= "01101100";
    expr_543_wire_constant <= "00000000";
    array_obj_ref_506_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_506_gather_scatter_ack_0 <= array_obj_ref_506_gather_scatter_req_0;
      aggregated_sig <= expr_507_wire_constant;
      array_obj_ref_506_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_510_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_510_gather_scatter_ack_0 <= array_obj_ref_510_gather_scatter_req_0;
      aggregated_sig <= expr_511_wire_constant;
      array_obj_ref_510_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_514_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_514_gather_scatter_ack_0 <= array_obj_ref_514_gather_scatter_req_0;
      aggregated_sig <= expr_515_wire_constant;
      array_obj_ref_514_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_518_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_518_gather_scatter_ack_0 <= array_obj_ref_518_gather_scatter_req_0;
      aggregated_sig <= expr_519_wire_constant;
      array_obj_ref_518_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_522_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_522_gather_scatter_ack_0 <= array_obj_ref_522_gather_scatter_req_0;
      aggregated_sig <= expr_523_wire_constant;
      array_obj_ref_522_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_526_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_526_gather_scatter_ack_0 <= array_obj_ref_526_gather_scatter_req_0;
      aggregated_sig <= expr_527_wire_constant;
      array_obj_ref_526_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_530_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_530_gather_scatter_ack_0 <= array_obj_ref_530_gather_scatter_req_0;
      aggregated_sig <= expr_531_wire_constant;
      array_obj_ref_530_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_534_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_534_gather_scatter_ack_0 <= array_obj_ref_534_gather_scatter_req_0;
      aggregated_sig <= expr_535_wire_constant;
      array_obj_ref_534_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_538_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_538_gather_scatter_ack_0 <= array_obj_ref_538_gather_scatter_req_0;
      aggregated_sig <= expr_539_wire_constant;
      array_obj_ref_538_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_542_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_542_gather_scatter_ack_0 <= array_obj_ref_542_gather_scatter_req_0;
      aggregated_sig <= expr_543_wire_constant;
      array_obj_ref_542_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_506_store_0 array_obj_ref_510_store_0 array_obj_ref_514_store_0 array_obj_ref_518_store_0 array_obj_ref_522_store_0 array_obj_ref_526_store_0 array_obj_ref_530_store_0 array_obj_ref_534_store_0 array_obj_ref_538_store_0 array_obj_ref_542_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(39 downto 0);
      signal data_in: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 9 downto 0);
      -- 
    begin -- 
      reqL(9) <= array_obj_ref_506_store_0_req_0;
      reqL(8) <= array_obj_ref_510_store_0_req_0;
      reqL(7) <= array_obj_ref_514_store_0_req_0;
      reqL(6) <= array_obj_ref_518_store_0_req_0;
      reqL(5) <= array_obj_ref_522_store_0_req_0;
      reqL(4) <= array_obj_ref_526_store_0_req_0;
      reqL(3) <= array_obj_ref_530_store_0_req_0;
      reqL(2) <= array_obj_ref_534_store_0_req_0;
      reqL(1) <= array_obj_ref_538_store_0_req_0;
      reqL(0) <= array_obj_ref_542_store_0_req_0;
      array_obj_ref_506_store_0_ack_0 <= ackL(9);
      array_obj_ref_510_store_0_ack_0 <= ackL(8);
      array_obj_ref_514_store_0_ack_0 <= ackL(7);
      array_obj_ref_518_store_0_ack_0 <= ackL(6);
      array_obj_ref_522_store_0_ack_0 <= ackL(5);
      array_obj_ref_526_store_0_ack_0 <= ackL(4);
      array_obj_ref_530_store_0_ack_0 <= ackL(3);
      array_obj_ref_534_store_0_ack_0 <= ackL(2);
      array_obj_ref_538_store_0_ack_0 <= ackL(1);
      array_obj_ref_542_store_0_ack_0 <= ackL(0);
      reqR(9) <= array_obj_ref_506_store_0_req_1;
      reqR(8) <= array_obj_ref_510_store_0_req_1;
      reqR(7) <= array_obj_ref_514_store_0_req_1;
      reqR(6) <= array_obj_ref_518_store_0_req_1;
      reqR(5) <= array_obj_ref_522_store_0_req_1;
      reqR(4) <= array_obj_ref_526_store_0_req_1;
      reqR(3) <= array_obj_ref_530_store_0_req_1;
      reqR(2) <= array_obj_ref_534_store_0_req_1;
      reqR(1) <= array_obj_ref_538_store_0_req_1;
      reqR(0) <= array_obj_ref_542_store_0_req_1;
      array_obj_ref_506_store_0_ack_1 <= ackR(9);
      array_obj_ref_510_store_0_ack_1 <= ackR(8);
      array_obj_ref_514_store_0_ack_1 <= ackR(7);
      array_obj_ref_518_store_0_ack_1 <= ackR(6);
      array_obj_ref_522_store_0_ack_1 <= ackR(5);
      array_obj_ref_526_store_0_ack_1 <= ackR(4);
      array_obj_ref_530_store_0_ack_1 <= ackR(3);
      array_obj_ref_534_store_0_ack_1 <= ackR(2);
      array_obj_ref_538_store_0_ack_1 <= ackR(1);
      array_obj_ref_542_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_506_word_address_0 & array_obj_ref_510_word_address_0 & array_obj_ref_514_word_address_0 & array_obj_ref_518_word_address_0 & array_obj_ref_522_word_address_0 & array_obj_ref_526_word_address_0 & array_obj_ref_530_word_address_0 & array_obj_ref_534_word_address_0 & array_obj_ref_538_word_address_0 & array_obj_ref_542_word_address_0;
      data_in <= array_obj_ref_506_data_0 & array_obj_ref_510_data_0 & array_obj_ref_514_data_0 & array_obj_ref_518_data_0 & array_obj_ref_522_data_0 & array_obj_ref_526_data_0 & array_obj_ref_530_data_0 & array_obj_ref_534_data_0 & array_obj_ref_538_data_0 & array_obj_ref_542_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 10,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(3 downto 0),
          mdata => memory_space_10_sr_data(7 downto 0),
          mtag => memory_space_10_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 10,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr15 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_11_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_11_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr15;
architecture Default of default_initializer_xx_xstr15 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr15_CP_2355_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_548_gather_scatter_req_0 : boolean;
  signal array_obj_ref_548_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_548_store_0_req_0 : boolean;
  signal array_obj_ref_548_store_0_ack_0 : boolean;
  signal array_obj_ref_548_store_0_req_1 : boolean;
  signal array_obj_ref_548_store_0_ack_1 : boolean;
  signal array_obj_ref_552_gather_scatter_req_0 : boolean;
  signal array_obj_ref_552_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_552_store_0_req_0 : boolean;
  signal array_obj_ref_552_store_0_ack_0 : boolean;
  signal array_obj_ref_552_store_0_req_1 : boolean;
  signal array_obj_ref_552_store_0_ack_1 : boolean;
  signal array_obj_ref_556_gather_scatter_req_0 : boolean;
  signal array_obj_ref_556_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_556_store_0_req_0 : boolean;
  signal array_obj_ref_556_store_0_ack_0 : boolean;
  signal array_obj_ref_556_store_0_req_1 : boolean;
  signal array_obj_ref_556_store_0_ack_1 : boolean;
  signal array_obj_ref_560_gather_scatter_req_0 : boolean;
  signal array_obj_ref_560_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_560_store_0_req_0 : boolean;
  signal array_obj_ref_560_store_0_ack_0 : boolean;
  signal array_obj_ref_560_store_0_req_1 : boolean;
  signal array_obj_ref_560_store_0_ack_1 : boolean;
  signal array_obj_ref_564_gather_scatter_req_0 : boolean;
  signal array_obj_ref_564_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_564_store_0_req_0 : boolean;
  signal array_obj_ref_564_store_0_ack_0 : boolean;
  signal array_obj_ref_564_store_0_req_1 : boolean;
  signal array_obj_ref_564_store_0_ack_1 : boolean;
  signal array_obj_ref_568_gather_scatter_req_0 : boolean;
  signal array_obj_ref_568_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_568_store_0_req_0 : boolean;
  signal array_obj_ref_568_store_0_ack_0 : boolean;
  signal array_obj_ref_568_store_0_req_1 : boolean;
  signal array_obj_ref_568_store_0_ack_1 : boolean;
  signal array_obj_ref_572_gather_scatter_req_0 : boolean;
  signal array_obj_ref_572_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_572_store_0_req_0 : boolean;
  signal array_obj_ref_572_store_0_ack_0 : boolean;
  signal array_obj_ref_572_store_0_req_1 : boolean;
  signal array_obj_ref_572_store_0_ack_1 : boolean;
  signal array_obj_ref_576_gather_scatter_req_0 : boolean;
  signal array_obj_ref_576_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_576_store_0_req_0 : boolean;
  signal array_obj_ref_576_store_0_ack_0 : boolean;
  signal array_obj_ref_576_store_0_req_1 : boolean;
  signal array_obj_ref_576_store_0_ack_1 : boolean;
  signal array_obj_ref_580_gather_scatter_req_0 : boolean;
  signal array_obj_ref_580_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_580_store_0_req_0 : boolean;
  signal array_obj_ref_580_store_0_ack_0 : boolean;
  signal array_obj_ref_580_store_0_req_1 : boolean;
  signal array_obj_ref_580_store_0_ack_1 : boolean;
  signal array_obj_ref_584_gather_scatter_req_0 : boolean;
  signal array_obj_ref_584_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_584_store_0_req_0 : boolean;
  signal array_obj_ref_584_store_0_ack_0 : boolean;
  signal array_obj_ref_584_store_0_req_1 : boolean;
  signal array_obj_ref_584_store_0_ack_1 : boolean;
  signal array_obj_ref_588_gather_scatter_req_0 : boolean;
  signal array_obj_ref_588_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_588_store_0_req_0 : boolean;
  signal array_obj_ref_588_store_0_ack_0 : boolean;
  signal array_obj_ref_588_store_0_req_1 : boolean;
  signal array_obj_ref_588_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 11 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr15_CP_2355: Block -- control-path 
    signal cp_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(33);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(33), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_548_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_548_gather_scatter_ack_0;
    array_obj_ref_548_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_548_store_0_ack_0;
    array_obj_ref_548_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_548_store_0_ack_1;
    array_obj_ref_552_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_552_gather_scatter_ack_0;
    array_obj_ref_552_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_552_store_0_ack_0;
    array_obj_ref_552_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_552_store_0_ack_1;
    array_obj_ref_556_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_556_gather_scatter_ack_0;
    array_obj_ref_556_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_556_store_0_ack_0;
    array_obj_ref_556_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_556_store_0_ack_1;
    array_obj_ref_560_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_560_gather_scatter_ack_0;
    array_obj_ref_560_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_560_store_0_ack_0;
    array_obj_ref_560_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_560_store_0_ack_1;
    array_obj_ref_564_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_564_gather_scatter_ack_0;
    array_obj_ref_564_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_564_store_0_ack_0;
    array_obj_ref_564_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_564_store_0_ack_1;
    array_obj_ref_568_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_568_gather_scatter_ack_0;
    array_obj_ref_568_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_568_store_0_ack_0;
    array_obj_ref_568_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_568_store_0_ack_1;
    array_obj_ref_572_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_572_gather_scatter_ack_0;
    array_obj_ref_572_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_572_store_0_ack_0;
    array_obj_ref_572_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_572_store_0_ack_1;
    array_obj_ref_576_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_576_gather_scatter_ack_0;
    array_obj_ref_576_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_576_store_0_ack_0;
    array_obj_ref_576_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_576_store_0_ack_1;
    array_obj_ref_580_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_580_gather_scatter_ack_0;
    array_obj_ref_580_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_580_store_0_ack_0;
    array_obj_ref_580_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_580_store_0_ack_1;
    array_obj_ref_584_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_584_gather_scatter_ack_0;
    array_obj_ref_584_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_584_store_0_ack_0;
    array_obj_ref_584_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_584_store_0_ack_1;
    array_obj_ref_588_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_588_gather_scatter_ack_0;
    array_obj_ref_588_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_588_store_0_ack_0;
    array_obj_ref_588_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_588_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_548_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_548_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_552_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_552_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_556_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_556_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_560_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_564_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_564_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_568_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_568_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_572_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_572_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_576_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_576_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_580_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_580_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_584_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_584_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_588_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_588_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_549_wire_constant : std_logic_vector(7 downto 0);
    signal expr_553_wire_constant : std_logic_vector(7 downto 0);
    signal expr_557_wire_constant : std_logic_vector(7 downto 0);
    signal expr_561_wire_constant : std_logic_vector(7 downto 0);
    signal expr_565_wire_constant : std_logic_vector(7 downto 0);
    signal expr_569_wire_constant : std_logic_vector(7 downto 0);
    signal expr_573_wire_constant : std_logic_vector(7 downto 0);
    signal expr_577_wire_constant : std_logic_vector(7 downto 0);
    signal expr_581_wire_constant : std_logic_vector(7 downto 0);
    signal expr_585_wire_constant : std_logic_vector(7 downto 0);
    signal expr_589_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_548_word_address_0 <= "0000";
    array_obj_ref_552_word_address_0 <= "0001";
    array_obj_ref_556_word_address_0 <= "0010";
    array_obj_ref_560_word_address_0 <= "0011";
    array_obj_ref_564_word_address_0 <= "0100";
    array_obj_ref_568_word_address_0 <= "0101";
    array_obj_ref_572_word_address_0 <= "0110";
    array_obj_ref_576_word_address_0 <= "0111";
    array_obj_ref_580_word_address_0 <= "1000";
    array_obj_ref_584_word_address_0 <= "1001";
    array_obj_ref_588_word_address_0 <= "1010";
    expr_549_wire_constant <= "01110000";
    expr_553_wire_constant <= "01101011";
    expr_557_wire_constant <= "01110100";
    expr_561_wire_constant <= "01011111";
    expr_565_wire_constant <= "01101100";
    expr_569_wire_constant <= "01100101";
    expr_573_wire_constant <= "01101110";
    expr_577_wire_constant <= "01100111";
    expr_581_wire_constant <= "01110100";
    expr_585_wire_constant <= "01101000";
    expr_589_wire_constant <= "00000000";
    array_obj_ref_548_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_548_gather_scatter_ack_0 <= array_obj_ref_548_gather_scatter_req_0;
      aggregated_sig <= expr_549_wire_constant;
      array_obj_ref_548_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_552_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_552_gather_scatter_ack_0 <= array_obj_ref_552_gather_scatter_req_0;
      aggregated_sig <= expr_553_wire_constant;
      array_obj_ref_552_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_556_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_556_gather_scatter_ack_0 <= array_obj_ref_556_gather_scatter_req_0;
      aggregated_sig <= expr_557_wire_constant;
      array_obj_ref_556_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_560_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_560_gather_scatter_ack_0 <= array_obj_ref_560_gather_scatter_req_0;
      aggregated_sig <= expr_561_wire_constant;
      array_obj_ref_560_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_564_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_564_gather_scatter_ack_0 <= array_obj_ref_564_gather_scatter_req_0;
      aggregated_sig <= expr_565_wire_constant;
      array_obj_ref_564_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_568_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_568_gather_scatter_ack_0 <= array_obj_ref_568_gather_scatter_req_0;
      aggregated_sig <= expr_569_wire_constant;
      array_obj_ref_568_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_572_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_572_gather_scatter_ack_0 <= array_obj_ref_572_gather_scatter_req_0;
      aggregated_sig <= expr_573_wire_constant;
      array_obj_ref_572_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_576_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_576_gather_scatter_ack_0 <= array_obj_ref_576_gather_scatter_req_0;
      aggregated_sig <= expr_577_wire_constant;
      array_obj_ref_576_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_580_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_580_gather_scatter_ack_0 <= array_obj_ref_580_gather_scatter_req_0;
      aggregated_sig <= expr_581_wire_constant;
      array_obj_ref_580_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_584_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_584_gather_scatter_ack_0 <= array_obj_ref_584_gather_scatter_req_0;
      aggregated_sig <= expr_585_wire_constant;
      array_obj_ref_584_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_588_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_588_gather_scatter_ack_0 <= array_obj_ref_588_gather_scatter_req_0;
      aggregated_sig <= expr_589_wire_constant;
      array_obj_ref_588_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_576_store_0 array_obj_ref_584_store_0 array_obj_ref_564_store_0 array_obj_ref_560_store_0 array_obj_ref_572_store_0 array_obj_ref_588_store_0 array_obj_ref_580_store_0 array_obj_ref_556_store_0 array_obj_ref_552_store_0 array_obj_ref_568_store_0 array_obj_ref_548_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(43 downto 0);
      signal data_in: std_logic_vector(87 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 10 downto 0);
      -- 
    begin -- 
      reqL(10) <= array_obj_ref_576_store_0_req_0;
      reqL(9) <= array_obj_ref_584_store_0_req_0;
      reqL(8) <= array_obj_ref_564_store_0_req_0;
      reqL(7) <= array_obj_ref_560_store_0_req_0;
      reqL(6) <= array_obj_ref_572_store_0_req_0;
      reqL(5) <= array_obj_ref_588_store_0_req_0;
      reqL(4) <= array_obj_ref_580_store_0_req_0;
      reqL(3) <= array_obj_ref_556_store_0_req_0;
      reqL(2) <= array_obj_ref_552_store_0_req_0;
      reqL(1) <= array_obj_ref_568_store_0_req_0;
      reqL(0) <= array_obj_ref_548_store_0_req_0;
      array_obj_ref_576_store_0_ack_0 <= ackL(10);
      array_obj_ref_584_store_0_ack_0 <= ackL(9);
      array_obj_ref_564_store_0_ack_0 <= ackL(8);
      array_obj_ref_560_store_0_ack_0 <= ackL(7);
      array_obj_ref_572_store_0_ack_0 <= ackL(6);
      array_obj_ref_588_store_0_ack_0 <= ackL(5);
      array_obj_ref_580_store_0_ack_0 <= ackL(4);
      array_obj_ref_556_store_0_ack_0 <= ackL(3);
      array_obj_ref_552_store_0_ack_0 <= ackL(2);
      array_obj_ref_568_store_0_ack_0 <= ackL(1);
      array_obj_ref_548_store_0_ack_0 <= ackL(0);
      reqR(10) <= array_obj_ref_576_store_0_req_1;
      reqR(9) <= array_obj_ref_584_store_0_req_1;
      reqR(8) <= array_obj_ref_564_store_0_req_1;
      reqR(7) <= array_obj_ref_560_store_0_req_1;
      reqR(6) <= array_obj_ref_572_store_0_req_1;
      reqR(5) <= array_obj_ref_588_store_0_req_1;
      reqR(4) <= array_obj_ref_580_store_0_req_1;
      reqR(3) <= array_obj_ref_556_store_0_req_1;
      reqR(2) <= array_obj_ref_552_store_0_req_1;
      reqR(1) <= array_obj_ref_568_store_0_req_1;
      reqR(0) <= array_obj_ref_548_store_0_req_1;
      array_obj_ref_576_store_0_ack_1 <= ackR(10);
      array_obj_ref_584_store_0_ack_1 <= ackR(9);
      array_obj_ref_564_store_0_ack_1 <= ackR(8);
      array_obj_ref_560_store_0_ack_1 <= ackR(7);
      array_obj_ref_572_store_0_ack_1 <= ackR(6);
      array_obj_ref_588_store_0_ack_1 <= ackR(5);
      array_obj_ref_580_store_0_ack_1 <= ackR(4);
      array_obj_ref_556_store_0_ack_1 <= ackR(3);
      array_obj_ref_552_store_0_ack_1 <= ackR(2);
      array_obj_ref_568_store_0_ack_1 <= ackR(1);
      array_obj_ref_548_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_576_word_address_0 & array_obj_ref_584_word_address_0 & array_obj_ref_564_word_address_0 & array_obj_ref_560_word_address_0 & array_obj_ref_572_word_address_0 & array_obj_ref_588_word_address_0 & array_obj_ref_580_word_address_0 & array_obj_ref_556_word_address_0 & array_obj_ref_552_word_address_0 & array_obj_ref_568_word_address_0 & array_obj_ref_548_word_address_0;
      data_in <= array_obj_ref_576_data_0 & array_obj_ref_584_data_0 & array_obj_ref_564_data_0 & array_obj_ref_560_data_0 & array_obj_ref_572_data_0 & array_obj_ref_588_data_0 & array_obj_ref_580_data_0 & array_obj_ref_556_data_0 & array_obj_ref_552_data_0 & array_obj_ref_568_data_0 & array_obj_ref_548_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 11,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_11_sr_req(0),
          mack => memory_space_11_sr_ack(0),
          maddr => memory_space_11_sr_addr(3 downto 0),
          mdata => memory_space_11_sr_data(7 downto 0),
          mtag => memory_space_11_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 11,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_11_sc_req(0),
          mack => memory_space_11_sc_ack(0),
          mtag => memory_space_11_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_12_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_12_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_12_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_12_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_12_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_12_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr2;
architecture Default of default_initializer_xx_xstr2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr2_CP_2589_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_622_store_0_req_0 : boolean;
  signal array_obj_ref_626_gather_scatter_req_0 : boolean;
  signal array_obj_ref_614_store_0_req_1 : boolean;
  signal array_obj_ref_610_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_602_store_0_ack_1 : boolean;
  signal array_obj_ref_638_store_0_req_1 : boolean;
  signal array_obj_ref_614_store_0_req_0 : boolean;
  signal array_obj_ref_598_store_0_req_1 : boolean;
  signal array_obj_ref_634_gather_scatter_req_0 : boolean;
  signal array_obj_ref_634_store_0_ack_1 : boolean;
  signal array_obj_ref_622_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_630_store_0_req_1 : boolean;
  signal array_obj_ref_638_gather_scatter_req_0 : boolean;
  signal array_obj_ref_638_store_0_ack_0 : boolean;
  signal array_obj_ref_594_gather_scatter_req_0 : boolean;
  signal array_obj_ref_594_store_0_ack_0 : boolean;
  signal array_obj_ref_606_store_0_ack_1 : boolean;
  signal array_obj_ref_622_store_0_ack_0 : boolean;
  signal array_obj_ref_630_store_0_ack_1 : boolean;
  signal array_obj_ref_610_store_0_ack_1 : boolean;
  signal array_obj_ref_606_store_0_req_0 : boolean;
  signal array_obj_ref_610_store_0_req_1 : boolean;
  signal array_obj_ref_614_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_606_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_610_gather_scatter_req_0 : boolean;
  signal array_obj_ref_626_store_0_ack_1 : boolean;
  signal array_obj_ref_634_store_0_ack_0 : boolean;
  signal array_obj_ref_622_store_0_req_1 : boolean;
  signal array_obj_ref_614_gather_scatter_req_0 : boolean;
  signal array_obj_ref_594_store_0_ack_1 : boolean;
  signal array_obj_ref_598_store_0_req_0 : boolean;
  signal array_obj_ref_602_store_0_req_0 : boolean;
  signal array_obj_ref_638_store_0_ack_1 : boolean;
  signal array_obj_ref_598_store_0_ack_1 : boolean;
  signal array_obj_ref_602_store_0_ack_0 : boolean;
  signal array_obj_ref_634_store_0_req_0 : boolean;
  signal array_obj_ref_614_store_0_ack_0 : boolean;
  signal array_obj_ref_614_store_0_ack_1 : boolean;
  signal array_obj_ref_634_store_0_req_1 : boolean;
  signal array_obj_ref_622_gather_scatter_req_0 : boolean;
  signal array_obj_ref_626_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_638_store_0_req_0 : boolean;
  signal array_obj_ref_602_gather_scatter_req_0 : boolean;
  signal array_obj_ref_626_store_0_req_0 : boolean;
  signal array_obj_ref_606_store_0_req_1 : boolean;
  signal array_obj_ref_602_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_594_store_0_req_0 : boolean;
  signal array_obj_ref_618_store_0_req_0 : boolean;
  signal array_obj_ref_610_store_0_ack_0 : boolean;
  signal array_obj_ref_626_store_0_req_1 : boolean;
  signal array_obj_ref_598_store_0_ack_0 : boolean;
  signal array_obj_ref_630_store_0_ack_0 : boolean;
  signal array_obj_ref_610_store_0_req_0 : boolean;
  signal array_obj_ref_594_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_618_gather_scatter_req_0 : boolean;
  signal array_obj_ref_618_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_630_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_634_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_598_gather_scatter_req_0 : boolean;
  signal array_obj_ref_618_store_0_ack_1 : boolean;
  signal array_obj_ref_626_store_0_ack_0 : boolean;
  signal array_obj_ref_618_store_0_ack_0 : boolean;
  signal array_obj_ref_598_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_606_gather_scatter_req_0 : boolean;
  signal array_obj_ref_618_store_0_req_1 : boolean;
  signal array_obj_ref_630_gather_scatter_req_0 : boolean;
  signal array_obj_ref_594_store_0_req_1 : boolean;
  signal array_obj_ref_630_store_0_req_0 : boolean;
  signal array_obj_ref_638_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_606_store_0_ack_0 : boolean;
  signal array_obj_ref_602_store_0_req_1 : boolean;
  signal array_obj_ref_622_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 12 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr2_CP_2589: Block -- control-path 
    signal cp_elements: BooleanArray(36 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(36);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(36), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_594_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_594_gather_scatter_ack_0;
    array_obj_ref_594_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_594_store_0_ack_0;
    array_obj_ref_594_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_594_store_0_ack_1;
    array_obj_ref_598_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_598_gather_scatter_ack_0;
    array_obj_ref_598_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_598_store_0_ack_0;
    array_obj_ref_598_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_598_store_0_ack_1;
    array_obj_ref_602_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_602_gather_scatter_ack_0;
    array_obj_ref_602_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_602_store_0_ack_0;
    array_obj_ref_602_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_602_store_0_ack_1;
    array_obj_ref_606_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_606_gather_scatter_ack_0;
    array_obj_ref_606_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_606_store_0_ack_0;
    array_obj_ref_606_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_606_store_0_ack_1;
    array_obj_ref_610_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_610_gather_scatter_ack_0;
    array_obj_ref_610_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_610_store_0_ack_0;
    array_obj_ref_610_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_610_store_0_ack_1;
    array_obj_ref_614_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_614_gather_scatter_ack_0;
    array_obj_ref_614_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_614_store_0_ack_0;
    array_obj_ref_614_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_614_store_0_ack_1;
    array_obj_ref_618_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_618_gather_scatter_ack_0;
    array_obj_ref_618_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_618_store_0_ack_0;
    array_obj_ref_618_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_618_store_0_ack_1;
    array_obj_ref_622_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_622_gather_scatter_ack_0;
    array_obj_ref_622_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_622_store_0_ack_0;
    array_obj_ref_622_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_622_store_0_ack_1;
    array_obj_ref_626_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_626_gather_scatter_ack_0;
    array_obj_ref_626_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_626_store_0_ack_0;
    array_obj_ref_626_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_626_store_0_ack_1;
    array_obj_ref_630_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_630_gather_scatter_ack_0;
    array_obj_ref_630_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_630_store_0_ack_0;
    array_obj_ref_630_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_630_store_0_ack_1;
    array_obj_ref_634_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_634_gather_scatter_ack_0;
    array_obj_ref_634_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_634_store_0_ack_0;
    array_obj_ref_634_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_634_store_0_ack_1;
    array_obj_ref_638_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_638_gather_scatter_ack_0;
    array_obj_ref_638_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_638_store_0_ack_0;
    array_obj_ref_638_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_638_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_594_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_594_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_598_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_598_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_602_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_602_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_606_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_606_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_610_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_610_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_614_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_614_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_618_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_618_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_622_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_622_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_626_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_626_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_630_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_630_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_634_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_634_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_638_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_638_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_595_wire_constant : std_logic_vector(7 downto 0);
    signal expr_599_wire_constant : std_logic_vector(7 downto 0);
    signal expr_603_wire_constant : std_logic_vector(7 downto 0);
    signal expr_607_wire_constant : std_logic_vector(7 downto 0);
    signal expr_611_wire_constant : std_logic_vector(7 downto 0);
    signal expr_615_wire_constant : std_logic_vector(7 downto 0);
    signal expr_619_wire_constant : std_logic_vector(7 downto 0);
    signal expr_623_wire_constant : std_logic_vector(7 downto 0);
    signal expr_627_wire_constant : std_logic_vector(7 downto 0);
    signal expr_631_wire_constant : std_logic_vector(7 downto 0);
    signal expr_635_wire_constant : std_logic_vector(7 downto 0);
    signal expr_639_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_594_word_address_0 <= "0000";
    array_obj_ref_598_word_address_0 <= "0001";
    array_obj_ref_602_word_address_0 <= "0010";
    array_obj_ref_606_word_address_0 <= "0011";
    array_obj_ref_610_word_address_0 <= "0100";
    array_obj_ref_614_word_address_0 <= "0101";
    array_obj_ref_618_word_address_0 <= "0110";
    array_obj_ref_622_word_address_0 <= "0111";
    array_obj_ref_626_word_address_0 <= "1000";
    array_obj_ref_630_word_address_0 <= "1001";
    array_obj_ref_634_word_address_0 <= "1010";
    array_obj_ref_638_word_address_0 <= "1011";
    expr_595_wire_constant <= "01101111";
    expr_599_wire_constant <= "01110000";
    expr_603_wire_constant <= "01011111";
    expr_607_wire_constant <= "01101100";
    expr_611_wire_constant <= "01110101";
    expr_615_wire_constant <= "01110100";
    expr_619_wire_constant <= "01011111";
    expr_623_wire_constant <= "01100100";
    expr_627_wire_constant <= "01100001";
    expr_631_wire_constant <= "01110100";
    expr_635_wire_constant <= "01100001";
    expr_639_wire_constant <= "00000000";
    array_obj_ref_594_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_594_gather_scatter_ack_0 <= array_obj_ref_594_gather_scatter_req_0;
      aggregated_sig <= expr_595_wire_constant;
      array_obj_ref_594_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_598_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_598_gather_scatter_ack_0 <= array_obj_ref_598_gather_scatter_req_0;
      aggregated_sig <= expr_599_wire_constant;
      array_obj_ref_598_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_602_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_602_gather_scatter_ack_0 <= array_obj_ref_602_gather_scatter_req_0;
      aggregated_sig <= expr_603_wire_constant;
      array_obj_ref_602_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_606_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_606_gather_scatter_ack_0 <= array_obj_ref_606_gather_scatter_req_0;
      aggregated_sig <= expr_607_wire_constant;
      array_obj_ref_606_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_610_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_610_gather_scatter_ack_0 <= array_obj_ref_610_gather_scatter_req_0;
      aggregated_sig <= expr_611_wire_constant;
      array_obj_ref_610_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_614_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_614_gather_scatter_ack_0 <= array_obj_ref_614_gather_scatter_req_0;
      aggregated_sig <= expr_615_wire_constant;
      array_obj_ref_614_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_618_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_618_gather_scatter_ack_0 <= array_obj_ref_618_gather_scatter_req_0;
      aggregated_sig <= expr_619_wire_constant;
      array_obj_ref_618_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_622_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_622_gather_scatter_ack_0 <= array_obj_ref_622_gather_scatter_req_0;
      aggregated_sig <= expr_623_wire_constant;
      array_obj_ref_622_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_626_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_626_gather_scatter_ack_0 <= array_obj_ref_626_gather_scatter_req_0;
      aggregated_sig <= expr_627_wire_constant;
      array_obj_ref_626_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_630_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_630_gather_scatter_ack_0 <= array_obj_ref_630_gather_scatter_req_0;
      aggregated_sig <= expr_631_wire_constant;
      array_obj_ref_630_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_634_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_634_gather_scatter_ack_0 <= array_obj_ref_634_gather_scatter_req_0;
      aggregated_sig <= expr_635_wire_constant;
      array_obj_ref_634_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_638_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_638_gather_scatter_ack_0 <= array_obj_ref_638_gather_scatter_req_0;
      aggregated_sig <= expr_639_wire_constant;
      array_obj_ref_638_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_618_store_0 array_obj_ref_614_store_0 array_obj_ref_594_store_0 array_obj_ref_602_store_0 array_obj_ref_598_store_0 array_obj_ref_622_store_0 array_obj_ref_606_store_0 array_obj_ref_610_store_0 array_obj_ref_626_store_0 array_obj_ref_630_store_0 array_obj_ref_634_store_0 array_obj_ref_638_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(47 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      reqL(11) <= array_obj_ref_618_store_0_req_0;
      reqL(10) <= array_obj_ref_614_store_0_req_0;
      reqL(9) <= array_obj_ref_594_store_0_req_0;
      reqL(8) <= array_obj_ref_602_store_0_req_0;
      reqL(7) <= array_obj_ref_598_store_0_req_0;
      reqL(6) <= array_obj_ref_622_store_0_req_0;
      reqL(5) <= array_obj_ref_606_store_0_req_0;
      reqL(4) <= array_obj_ref_610_store_0_req_0;
      reqL(3) <= array_obj_ref_626_store_0_req_0;
      reqL(2) <= array_obj_ref_630_store_0_req_0;
      reqL(1) <= array_obj_ref_634_store_0_req_0;
      reqL(0) <= array_obj_ref_638_store_0_req_0;
      array_obj_ref_618_store_0_ack_0 <= ackL(11);
      array_obj_ref_614_store_0_ack_0 <= ackL(10);
      array_obj_ref_594_store_0_ack_0 <= ackL(9);
      array_obj_ref_602_store_0_ack_0 <= ackL(8);
      array_obj_ref_598_store_0_ack_0 <= ackL(7);
      array_obj_ref_622_store_0_ack_0 <= ackL(6);
      array_obj_ref_606_store_0_ack_0 <= ackL(5);
      array_obj_ref_610_store_0_ack_0 <= ackL(4);
      array_obj_ref_626_store_0_ack_0 <= ackL(3);
      array_obj_ref_630_store_0_ack_0 <= ackL(2);
      array_obj_ref_634_store_0_ack_0 <= ackL(1);
      array_obj_ref_638_store_0_ack_0 <= ackL(0);
      reqR(11) <= array_obj_ref_618_store_0_req_1;
      reqR(10) <= array_obj_ref_614_store_0_req_1;
      reqR(9) <= array_obj_ref_594_store_0_req_1;
      reqR(8) <= array_obj_ref_602_store_0_req_1;
      reqR(7) <= array_obj_ref_598_store_0_req_1;
      reqR(6) <= array_obj_ref_622_store_0_req_1;
      reqR(5) <= array_obj_ref_606_store_0_req_1;
      reqR(4) <= array_obj_ref_610_store_0_req_1;
      reqR(3) <= array_obj_ref_626_store_0_req_1;
      reqR(2) <= array_obj_ref_630_store_0_req_1;
      reqR(1) <= array_obj_ref_634_store_0_req_1;
      reqR(0) <= array_obj_ref_638_store_0_req_1;
      array_obj_ref_618_store_0_ack_1 <= ackR(11);
      array_obj_ref_614_store_0_ack_1 <= ackR(10);
      array_obj_ref_594_store_0_ack_1 <= ackR(9);
      array_obj_ref_602_store_0_ack_1 <= ackR(8);
      array_obj_ref_598_store_0_ack_1 <= ackR(7);
      array_obj_ref_622_store_0_ack_1 <= ackR(6);
      array_obj_ref_606_store_0_ack_1 <= ackR(5);
      array_obj_ref_610_store_0_ack_1 <= ackR(4);
      array_obj_ref_626_store_0_ack_1 <= ackR(3);
      array_obj_ref_630_store_0_ack_1 <= ackR(2);
      array_obj_ref_634_store_0_ack_1 <= ackR(1);
      array_obj_ref_638_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_618_word_address_0 & array_obj_ref_614_word_address_0 & array_obj_ref_594_word_address_0 & array_obj_ref_602_word_address_0 & array_obj_ref_598_word_address_0 & array_obj_ref_622_word_address_0 & array_obj_ref_606_word_address_0 & array_obj_ref_610_word_address_0 & array_obj_ref_626_word_address_0 & array_obj_ref_630_word_address_0 & array_obj_ref_634_word_address_0 & array_obj_ref_638_word_address_0;
      data_in <= array_obj_ref_618_data_0 & array_obj_ref_614_data_0 & array_obj_ref_594_data_0 & array_obj_ref_602_data_0 & array_obj_ref_598_data_0 & array_obj_ref_622_data_0 & array_obj_ref_606_data_0 & array_obj_ref_610_data_0 & array_obj_ref_626_data_0 & array_obj_ref_630_data_0 & array_obj_ref_634_data_0 & array_obj_ref_638_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 12,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_12_sr_req(0),
          mack => memory_space_12_sr_ack(0),
          maddr => memory_space_12_sr_addr(3 downto 0),
          mdata => memory_space_12_sr_data(7 downto 0),
          mtag => memory_space_12_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 12,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_12_sc_req(0),
          mack => memory_space_12_sc_ack(0),
          mtag => memory_space_12_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr3 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_13_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_13_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_13_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_13_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_13_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_13_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_13_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_13_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr3;
architecture Default of default_initializer_xx_xstr3 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr3_CP_2844_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_644_gather_scatter_req_0 : boolean;
  signal array_obj_ref_644_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_644_store_0_req_0 : boolean;
  signal array_obj_ref_644_store_0_ack_0 : boolean;
  signal array_obj_ref_644_store_0_req_1 : boolean;
  signal array_obj_ref_644_store_0_ack_1 : boolean;
  signal array_obj_ref_648_gather_scatter_req_0 : boolean;
  signal array_obj_ref_648_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_648_store_0_req_0 : boolean;
  signal array_obj_ref_648_store_0_ack_0 : boolean;
  signal array_obj_ref_648_store_0_req_1 : boolean;
  signal array_obj_ref_648_store_0_ack_1 : boolean;
  signal array_obj_ref_652_gather_scatter_req_0 : boolean;
  signal array_obj_ref_652_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_652_store_0_req_0 : boolean;
  signal array_obj_ref_652_store_0_ack_0 : boolean;
  signal array_obj_ref_652_store_0_req_1 : boolean;
  signal array_obj_ref_652_store_0_ack_1 : boolean;
  signal array_obj_ref_656_gather_scatter_req_0 : boolean;
  signal array_obj_ref_656_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_656_store_0_req_0 : boolean;
  signal array_obj_ref_656_store_0_ack_0 : boolean;
  signal array_obj_ref_656_store_0_req_1 : boolean;
  signal array_obj_ref_656_store_0_ack_1 : boolean;
  signal array_obj_ref_660_gather_scatter_req_0 : boolean;
  signal array_obj_ref_660_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_660_store_0_req_0 : boolean;
  signal array_obj_ref_660_store_0_ack_0 : boolean;
  signal array_obj_ref_660_store_0_req_1 : boolean;
  signal array_obj_ref_660_store_0_ack_1 : boolean;
  signal array_obj_ref_664_gather_scatter_req_0 : boolean;
  signal array_obj_ref_664_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_664_store_0_req_0 : boolean;
  signal array_obj_ref_664_store_0_ack_0 : boolean;
  signal array_obj_ref_664_store_0_req_1 : boolean;
  signal array_obj_ref_664_store_0_ack_1 : boolean;
  signal array_obj_ref_668_gather_scatter_req_0 : boolean;
  signal array_obj_ref_668_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_668_store_0_req_0 : boolean;
  signal array_obj_ref_668_store_0_ack_0 : boolean;
  signal array_obj_ref_668_store_0_req_1 : boolean;
  signal array_obj_ref_668_store_0_ack_1 : boolean;
  signal array_obj_ref_672_gather_scatter_req_0 : boolean;
  signal array_obj_ref_672_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_672_store_0_req_0 : boolean;
  signal array_obj_ref_672_store_0_ack_0 : boolean;
  signal array_obj_ref_672_store_0_req_1 : boolean;
  signal array_obj_ref_672_store_0_ack_1 : boolean;
  signal array_obj_ref_676_gather_scatter_req_0 : boolean;
  signal array_obj_ref_676_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_676_store_0_req_0 : boolean;
  signal array_obj_ref_676_store_0_ack_0 : boolean;
  signal array_obj_ref_676_store_0_req_1 : boolean;
  signal array_obj_ref_676_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 9 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr3_CP_2844: Block -- control-path 
    signal cp_elements: BooleanArray(27 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(27);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(27), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_644_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_644_gather_scatter_ack_0;
    array_obj_ref_644_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_644_store_0_ack_0;
    array_obj_ref_644_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_644_store_0_ack_1;
    array_obj_ref_648_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_648_gather_scatter_ack_0;
    array_obj_ref_648_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_648_store_0_ack_0;
    array_obj_ref_648_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_648_store_0_ack_1;
    array_obj_ref_652_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_652_gather_scatter_ack_0;
    array_obj_ref_652_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_652_store_0_ack_0;
    array_obj_ref_652_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_652_store_0_ack_1;
    array_obj_ref_656_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_656_gather_scatter_ack_0;
    array_obj_ref_656_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_656_store_0_ack_0;
    array_obj_ref_656_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_656_store_0_ack_1;
    array_obj_ref_660_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_660_gather_scatter_ack_0;
    array_obj_ref_660_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_660_store_0_ack_0;
    array_obj_ref_660_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_660_store_0_ack_1;
    array_obj_ref_664_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_664_gather_scatter_ack_0;
    array_obj_ref_664_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_664_store_0_ack_0;
    array_obj_ref_664_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_664_store_0_ack_1;
    array_obj_ref_668_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_668_gather_scatter_ack_0;
    array_obj_ref_668_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_668_store_0_ack_0;
    array_obj_ref_668_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_668_store_0_ack_1;
    array_obj_ref_672_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_672_gather_scatter_ack_0;
    array_obj_ref_672_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_672_store_0_ack_0;
    array_obj_ref_672_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_672_store_0_ack_1;
    array_obj_ref_676_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_676_gather_scatter_ack_0;
    array_obj_ref_676_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_676_store_0_ack_0;
    array_obj_ref_676_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_676_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_644_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_644_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_648_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_648_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_652_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_652_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_656_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_656_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_660_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_660_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_664_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_664_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_668_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_668_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_672_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_676_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_676_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_645_wire_constant : std_logic_vector(7 downto 0);
    signal expr_649_wire_constant : std_logic_vector(7 downto 0);
    signal expr_653_wire_constant : std_logic_vector(7 downto 0);
    signal expr_657_wire_constant : std_logic_vector(7 downto 0);
    signal expr_661_wire_constant : std_logic_vector(7 downto 0);
    signal expr_665_wire_constant : std_logic_vector(7 downto 0);
    signal expr_669_wire_constant : std_logic_vector(7 downto 0);
    signal expr_673_wire_constant : std_logic_vector(7 downto 0);
    signal expr_677_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_644_word_address_0 <= "0000";
    array_obj_ref_648_word_address_0 <= "0001";
    array_obj_ref_652_word_address_0 <= "0010";
    array_obj_ref_656_word_address_0 <= "0011";
    array_obj_ref_660_word_address_0 <= "0100";
    array_obj_ref_664_word_address_0 <= "0101";
    array_obj_ref_668_word_address_0 <= "0110";
    array_obj_ref_672_word_address_0 <= "0111";
    array_obj_ref_676_word_address_0 <= "1000";
    expr_645_wire_constant <= "01101111";
    expr_649_wire_constant <= "01110101";
    expr_653_wire_constant <= "01110100";
    expr_657_wire_constant <= "01011111";
    expr_661_wire_constant <= "01100011";
    expr_665_wire_constant <= "01110100";
    expr_669_wire_constant <= "01110010";
    expr_673_wire_constant <= "01101100";
    expr_677_wire_constant <= "00000000";
    array_obj_ref_644_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_644_gather_scatter_ack_0 <= array_obj_ref_644_gather_scatter_req_0;
      aggregated_sig <= expr_645_wire_constant;
      array_obj_ref_644_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_648_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_648_gather_scatter_ack_0 <= array_obj_ref_648_gather_scatter_req_0;
      aggregated_sig <= expr_649_wire_constant;
      array_obj_ref_648_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_652_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_652_gather_scatter_ack_0 <= array_obj_ref_652_gather_scatter_req_0;
      aggregated_sig <= expr_653_wire_constant;
      array_obj_ref_652_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_656_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_656_gather_scatter_ack_0 <= array_obj_ref_656_gather_scatter_req_0;
      aggregated_sig <= expr_657_wire_constant;
      array_obj_ref_656_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_660_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_660_gather_scatter_ack_0 <= array_obj_ref_660_gather_scatter_req_0;
      aggregated_sig <= expr_661_wire_constant;
      array_obj_ref_660_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_664_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_664_gather_scatter_ack_0 <= array_obj_ref_664_gather_scatter_req_0;
      aggregated_sig <= expr_665_wire_constant;
      array_obj_ref_664_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_668_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_668_gather_scatter_ack_0 <= array_obj_ref_668_gather_scatter_req_0;
      aggregated_sig <= expr_669_wire_constant;
      array_obj_ref_668_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_672_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_672_gather_scatter_ack_0 <= array_obj_ref_672_gather_scatter_req_0;
      aggregated_sig <= expr_673_wire_constant;
      array_obj_ref_672_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_676_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_676_gather_scatter_ack_0 <= array_obj_ref_676_gather_scatter_req_0;
      aggregated_sig <= expr_677_wire_constant;
      array_obj_ref_676_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_652_store_0 array_obj_ref_648_store_0 array_obj_ref_668_store_0 array_obj_ref_664_store_0 array_obj_ref_672_store_0 array_obj_ref_676_store_0 array_obj_ref_656_store_0 array_obj_ref_644_store_0 array_obj_ref_660_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(35 downto 0);
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 8 downto 0);
      -- 
    begin -- 
      reqL(8) <= array_obj_ref_652_store_0_req_0;
      reqL(7) <= array_obj_ref_648_store_0_req_0;
      reqL(6) <= array_obj_ref_668_store_0_req_0;
      reqL(5) <= array_obj_ref_664_store_0_req_0;
      reqL(4) <= array_obj_ref_672_store_0_req_0;
      reqL(3) <= array_obj_ref_676_store_0_req_0;
      reqL(2) <= array_obj_ref_656_store_0_req_0;
      reqL(1) <= array_obj_ref_644_store_0_req_0;
      reqL(0) <= array_obj_ref_660_store_0_req_0;
      array_obj_ref_652_store_0_ack_0 <= ackL(8);
      array_obj_ref_648_store_0_ack_0 <= ackL(7);
      array_obj_ref_668_store_0_ack_0 <= ackL(6);
      array_obj_ref_664_store_0_ack_0 <= ackL(5);
      array_obj_ref_672_store_0_ack_0 <= ackL(4);
      array_obj_ref_676_store_0_ack_0 <= ackL(3);
      array_obj_ref_656_store_0_ack_0 <= ackL(2);
      array_obj_ref_644_store_0_ack_0 <= ackL(1);
      array_obj_ref_660_store_0_ack_0 <= ackL(0);
      reqR(8) <= array_obj_ref_652_store_0_req_1;
      reqR(7) <= array_obj_ref_648_store_0_req_1;
      reqR(6) <= array_obj_ref_668_store_0_req_1;
      reqR(5) <= array_obj_ref_664_store_0_req_1;
      reqR(4) <= array_obj_ref_672_store_0_req_1;
      reqR(3) <= array_obj_ref_676_store_0_req_1;
      reqR(2) <= array_obj_ref_656_store_0_req_1;
      reqR(1) <= array_obj_ref_644_store_0_req_1;
      reqR(0) <= array_obj_ref_660_store_0_req_1;
      array_obj_ref_652_store_0_ack_1 <= ackR(8);
      array_obj_ref_648_store_0_ack_1 <= ackR(7);
      array_obj_ref_668_store_0_ack_1 <= ackR(6);
      array_obj_ref_664_store_0_ack_1 <= ackR(5);
      array_obj_ref_672_store_0_ack_1 <= ackR(4);
      array_obj_ref_676_store_0_ack_1 <= ackR(3);
      array_obj_ref_656_store_0_ack_1 <= ackR(2);
      array_obj_ref_644_store_0_ack_1 <= ackR(1);
      array_obj_ref_660_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_652_word_address_0 & array_obj_ref_648_word_address_0 & array_obj_ref_668_word_address_0 & array_obj_ref_664_word_address_0 & array_obj_ref_672_word_address_0 & array_obj_ref_676_word_address_0 & array_obj_ref_656_word_address_0 & array_obj_ref_644_word_address_0 & array_obj_ref_660_word_address_0;
      data_in <= array_obj_ref_652_data_0 & array_obj_ref_648_data_0 & array_obj_ref_668_data_0 & array_obj_ref_664_data_0 & array_obj_ref_672_data_0 & array_obj_ref_676_data_0 & array_obj_ref_656_data_0 & array_obj_ref_644_data_0 & array_obj_ref_660_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 9,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_13_sr_req(0),
          mack => memory_space_13_sr_ack(0),
          maddr => memory_space_13_sr_addr(3 downto 0),
          mdata => memory_space_13_sr_data(7 downto 0),
          mtag => memory_space_13_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 9,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_13_sc_req(0),
          mack => memory_space_13_sc_ack(0),
          mtag => memory_space_13_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_14_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_14_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_14_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_14_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_14_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_14_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_14_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_14_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr4;
architecture Default of default_initializer_xx_xstr4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr4_CP_3036_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_706_gather_scatter_req_0 : boolean;
  signal array_obj_ref_686_store_0_req_1 : boolean;
  signal array_obj_ref_698_store_0_req_0 : boolean;
  signal array_obj_ref_702_store_0_ack_1 : boolean;
  signal array_obj_ref_686_gather_scatter_req_0 : boolean;
  signal array_obj_ref_690_store_0_req_0 : boolean;
  signal array_obj_ref_714_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_682_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_682_store_0_ack_0 : boolean;
  signal array_obj_ref_702_store_0_ack_0 : boolean;
  signal array_obj_ref_714_store_0_ack_0 : boolean;
  signal array_obj_ref_682_store_0_req_1 : boolean;
  signal array_obj_ref_714_store_0_req_1 : boolean;
  signal array_obj_ref_714_store_0_req_0 : boolean;
  signal array_obj_ref_714_gather_scatter_req_0 : boolean;
  signal array_obj_ref_706_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_686_store_0_ack_0 : boolean;
  signal array_obj_ref_690_gather_scatter_req_0 : boolean;
  signal array_obj_ref_702_store_0_req_1 : boolean;
  signal array_obj_ref_702_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_686_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_694_store_0_ack_1 : boolean;
  signal array_obj_ref_698_gather_scatter_req_0 : boolean;
  signal array_obj_ref_682_store_0_req_0 : boolean;
  signal array_obj_ref_702_store_0_req_0 : boolean;
  signal array_obj_ref_682_gather_scatter_req_0 : boolean;
  signal array_obj_ref_682_store_0_ack_1 : boolean;
  signal array_obj_ref_698_store_0_ack_0 : boolean;
  signal array_obj_ref_702_gather_scatter_req_0 : boolean;
  signal array_obj_ref_690_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_698_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_690_store_0_ack_0 : boolean;
  signal array_obj_ref_714_store_0_ack_1 : boolean;
  signal array_obj_ref_686_store_0_req_0 : boolean;
  signal array_obj_ref_698_store_0_ack_1 : boolean;
  signal array_obj_ref_686_store_0_ack_1 : boolean;
  signal array_obj_ref_698_store_0_req_1 : boolean;
  signal array_obj_ref_706_store_0_req_0 : boolean;
  signal array_obj_ref_706_store_0_ack_0 : boolean;
  signal array_obj_ref_690_store_0_req_1 : boolean;
  signal array_obj_ref_706_store_0_req_1 : boolean;
  signal array_obj_ref_706_store_0_ack_1 : boolean;
  signal array_obj_ref_690_store_0_ack_1 : boolean;
  signal array_obj_ref_710_gather_scatter_req_0 : boolean;
  signal array_obj_ref_710_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_694_gather_scatter_req_0 : boolean;
  signal array_obj_ref_694_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_710_store_0_req_0 : boolean;
  signal array_obj_ref_710_store_0_ack_0 : boolean;
  signal array_obj_ref_710_store_0_req_1 : boolean;
  signal array_obj_ref_710_store_0_ack_1 : boolean;
  signal array_obj_ref_694_store_0_req_0 : boolean;
  signal array_obj_ref_694_store_0_ack_0 : boolean;
  signal array_obj_ref_694_store_0_req_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 9 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr4_CP_3036: Block -- control-path 
    signal cp_elements: BooleanArray(27 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(27);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(27), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_682_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_682_gather_scatter_ack_0;
    array_obj_ref_682_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_682_store_0_ack_0;
    array_obj_ref_682_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_682_store_0_ack_1;
    array_obj_ref_686_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_686_gather_scatter_ack_0;
    array_obj_ref_686_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_686_store_0_ack_0;
    array_obj_ref_686_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_686_store_0_ack_1;
    array_obj_ref_690_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_690_gather_scatter_ack_0;
    array_obj_ref_690_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_690_store_0_ack_0;
    array_obj_ref_690_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_690_store_0_ack_1;
    array_obj_ref_694_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_694_gather_scatter_ack_0;
    array_obj_ref_694_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_694_store_0_ack_0;
    array_obj_ref_694_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_694_store_0_ack_1;
    array_obj_ref_698_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_698_gather_scatter_ack_0;
    array_obj_ref_698_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_698_store_0_ack_0;
    array_obj_ref_698_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_698_store_0_ack_1;
    array_obj_ref_702_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_702_gather_scatter_ack_0;
    array_obj_ref_702_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_702_store_0_ack_0;
    array_obj_ref_702_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_702_store_0_ack_1;
    array_obj_ref_706_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_706_gather_scatter_ack_0;
    array_obj_ref_706_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_706_store_0_ack_0;
    array_obj_ref_706_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_706_store_0_ack_1;
    array_obj_ref_710_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_710_gather_scatter_ack_0;
    array_obj_ref_710_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_710_store_0_ack_0;
    array_obj_ref_710_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_710_store_0_ack_1;
    array_obj_ref_714_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_714_gather_scatter_ack_0;
    array_obj_ref_714_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_714_store_0_ack_0;
    array_obj_ref_714_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_714_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_682_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_682_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_686_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_686_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_690_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_690_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_694_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_694_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_698_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_702_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_702_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_706_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_706_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_710_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_710_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_714_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_714_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_683_wire_constant : std_logic_vector(7 downto 0);
    signal expr_687_wire_constant : std_logic_vector(7 downto 0);
    signal expr_691_wire_constant : std_logic_vector(7 downto 0);
    signal expr_695_wire_constant : std_logic_vector(7 downto 0);
    signal expr_699_wire_constant : std_logic_vector(7 downto 0);
    signal expr_703_wire_constant : std_logic_vector(7 downto 0);
    signal expr_707_wire_constant : std_logic_vector(7 downto 0);
    signal expr_711_wire_constant : std_logic_vector(7 downto 0);
    signal expr_715_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_682_word_address_0 <= "0000";
    array_obj_ref_686_word_address_0 <= "0001";
    array_obj_ref_690_word_address_0 <= "0010";
    array_obj_ref_694_word_address_0 <= "0011";
    array_obj_ref_698_word_address_0 <= "0100";
    array_obj_ref_702_word_address_0 <= "0101";
    array_obj_ref_706_word_address_0 <= "0110";
    array_obj_ref_710_word_address_0 <= "0111";
    array_obj_ref_714_word_address_0 <= "1000";
    expr_683_wire_constant <= "01101111";
    expr_687_wire_constant <= "01110101";
    expr_691_wire_constant <= "01110100";
    expr_695_wire_constant <= "01011111";
    expr_699_wire_constant <= "01100100";
    expr_703_wire_constant <= "01100001";
    expr_707_wire_constant <= "01110100";
    expr_711_wire_constant <= "01100001";
    expr_715_wire_constant <= "00000000";
    array_obj_ref_682_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_682_gather_scatter_ack_0 <= array_obj_ref_682_gather_scatter_req_0;
      aggregated_sig <= expr_683_wire_constant;
      array_obj_ref_682_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_686_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_686_gather_scatter_ack_0 <= array_obj_ref_686_gather_scatter_req_0;
      aggregated_sig <= expr_687_wire_constant;
      array_obj_ref_686_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_690_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_690_gather_scatter_ack_0 <= array_obj_ref_690_gather_scatter_req_0;
      aggregated_sig <= expr_691_wire_constant;
      array_obj_ref_690_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_694_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_694_gather_scatter_ack_0 <= array_obj_ref_694_gather_scatter_req_0;
      aggregated_sig <= expr_695_wire_constant;
      array_obj_ref_694_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_698_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_698_gather_scatter_ack_0 <= array_obj_ref_698_gather_scatter_req_0;
      aggregated_sig <= expr_699_wire_constant;
      array_obj_ref_698_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_702_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_702_gather_scatter_ack_0 <= array_obj_ref_702_gather_scatter_req_0;
      aggregated_sig <= expr_703_wire_constant;
      array_obj_ref_702_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_706_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_706_gather_scatter_ack_0 <= array_obj_ref_706_gather_scatter_req_0;
      aggregated_sig <= expr_707_wire_constant;
      array_obj_ref_706_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_710_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_710_gather_scatter_ack_0 <= array_obj_ref_710_gather_scatter_req_0;
      aggregated_sig <= expr_711_wire_constant;
      array_obj_ref_710_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_714_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_714_gather_scatter_ack_0 <= array_obj_ref_714_gather_scatter_req_0;
      aggregated_sig <= expr_715_wire_constant;
      array_obj_ref_714_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_702_store_0 array_obj_ref_706_store_0 array_obj_ref_694_store_0 array_obj_ref_698_store_0 array_obj_ref_714_store_0 array_obj_ref_682_store_0 array_obj_ref_686_store_0 array_obj_ref_690_store_0 array_obj_ref_710_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(35 downto 0);
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 8 downto 0);
      -- 
    begin -- 
      reqL(8) <= array_obj_ref_702_store_0_req_0;
      reqL(7) <= array_obj_ref_706_store_0_req_0;
      reqL(6) <= array_obj_ref_694_store_0_req_0;
      reqL(5) <= array_obj_ref_698_store_0_req_0;
      reqL(4) <= array_obj_ref_714_store_0_req_0;
      reqL(3) <= array_obj_ref_682_store_0_req_0;
      reqL(2) <= array_obj_ref_686_store_0_req_0;
      reqL(1) <= array_obj_ref_690_store_0_req_0;
      reqL(0) <= array_obj_ref_710_store_0_req_0;
      array_obj_ref_702_store_0_ack_0 <= ackL(8);
      array_obj_ref_706_store_0_ack_0 <= ackL(7);
      array_obj_ref_694_store_0_ack_0 <= ackL(6);
      array_obj_ref_698_store_0_ack_0 <= ackL(5);
      array_obj_ref_714_store_0_ack_0 <= ackL(4);
      array_obj_ref_682_store_0_ack_0 <= ackL(3);
      array_obj_ref_686_store_0_ack_0 <= ackL(2);
      array_obj_ref_690_store_0_ack_0 <= ackL(1);
      array_obj_ref_710_store_0_ack_0 <= ackL(0);
      reqR(8) <= array_obj_ref_702_store_0_req_1;
      reqR(7) <= array_obj_ref_706_store_0_req_1;
      reqR(6) <= array_obj_ref_694_store_0_req_1;
      reqR(5) <= array_obj_ref_698_store_0_req_1;
      reqR(4) <= array_obj_ref_714_store_0_req_1;
      reqR(3) <= array_obj_ref_682_store_0_req_1;
      reqR(2) <= array_obj_ref_686_store_0_req_1;
      reqR(1) <= array_obj_ref_690_store_0_req_1;
      reqR(0) <= array_obj_ref_710_store_0_req_1;
      array_obj_ref_702_store_0_ack_1 <= ackR(8);
      array_obj_ref_706_store_0_ack_1 <= ackR(7);
      array_obj_ref_694_store_0_ack_1 <= ackR(6);
      array_obj_ref_698_store_0_ack_1 <= ackR(5);
      array_obj_ref_714_store_0_ack_1 <= ackR(4);
      array_obj_ref_682_store_0_ack_1 <= ackR(3);
      array_obj_ref_686_store_0_ack_1 <= ackR(2);
      array_obj_ref_690_store_0_ack_1 <= ackR(1);
      array_obj_ref_710_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_702_word_address_0 & array_obj_ref_706_word_address_0 & array_obj_ref_694_word_address_0 & array_obj_ref_698_word_address_0 & array_obj_ref_714_word_address_0 & array_obj_ref_682_word_address_0 & array_obj_ref_686_word_address_0 & array_obj_ref_690_word_address_0 & array_obj_ref_710_word_address_0;
      data_in <= array_obj_ref_702_data_0 & array_obj_ref_706_data_0 & array_obj_ref_694_data_0 & array_obj_ref_698_data_0 & array_obj_ref_714_data_0 & array_obj_ref_682_data_0 & array_obj_ref_686_data_0 & array_obj_ref_690_data_0 & array_obj_ref_710_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 9,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_14_sr_req(0),
          mack => memory_space_14_sr_ack(0),
          maddr => memory_space_14_sr_addr(3 downto 0),
          mdata => memory_space_14_sr_data(7 downto 0),
          mtag => memory_space_14_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 9,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_14_sc_req(0),
          mack => memory_space_14_sc_ack(0),
          mtag => memory_space_14_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr5 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_15_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_15_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_15_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_15_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_15_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_15_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_15_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_15_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr5;
architecture Default of default_initializer_xx_xstr5 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr5_CP_3228_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_728_store_0_req_1 : boolean;
  signal array_obj_ref_728_store_0_ack_1 : boolean;
  signal array_obj_ref_724_store_0_req_1 : boolean;
  signal array_obj_ref_728_store_0_req_0 : boolean;
  signal array_obj_ref_720_store_0_ack_1 : boolean;
  signal array_obj_ref_720_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_720_store_0_req_0 : boolean;
  signal array_obj_ref_720_store_0_ack_0 : boolean;
  signal array_obj_ref_724_gather_scatter_req_0 : boolean;
  signal array_obj_ref_728_store_0_ack_0 : boolean;
  signal array_obj_ref_724_store_0_ack_1 : boolean;
  signal array_obj_ref_720_gather_scatter_req_0 : boolean;
  signal array_obj_ref_724_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_736_store_0_req_0 : boolean;
  signal array_obj_ref_736_store_0_ack_0 : boolean;
  signal array_obj_ref_736_store_0_req_1 : boolean;
  signal array_obj_ref_736_store_0_ack_1 : boolean;
  signal array_obj_ref_724_store_0_req_0 : boolean;
  signal array_obj_ref_724_store_0_ack_0 : boolean;
  signal array_obj_ref_728_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_728_gather_scatter_req_0 : boolean;
  signal array_obj_ref_748_gather_scatter_req_0 : boolean;
  signal array_obj_ref_748_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_764_store_0_req_0 : boolean;
  signal array_obj_ref_764_store_0_ack_0 : boolean;
  signal array_obj_ref_764_store_0_req_1 : boolean;
  signal array_obj_ref_764_store_0_ack_1 : boolean;
  signal array_obj_ref_736_gather_scatter_req_0 : boolean;
  signal array_obj_ref_736_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_744_store_0_req_1 : boolean;
  signal array_obj_ref_744_store_0_ack_1 : boolean;
  signal array_obj_ref_764_gather_scatter_req_0 : boolean;
  signal array_obj_ref_764_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_744_store_0_req_0 : boolean;
  signal array_obj_ref_744_store_0_ack_0 : boolean;
  signal array_obj_ref_760_store_0_req_0 : boolean;
  signal array_obj_ref_760_store_0_ack_0 : boolean;
  signal array_obj_ref_760_store_0_req_1 : boolean;
  signal array_obj_ref_760_store_0_ack_1 : boolean;
  signal array_obj_ref_744_gather_scatter_req_0 : boolean;
  signal array_obj_ref_744_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_760_gather_scatter_req_0 : boolean;
  signal array_obj_ref_760_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_756_store_0_ack_0 : boolean;
  signal array_obj_ref_756_store_0_req_1 : boolean;
  signal array_obj_ref_756_store_0_ack_1 : boolean;
  signal array_obj_ref_732_store_0_req_1 : boolean;
  signal array_obj_ref_732_store_0_ack_1 : boolean;
  signal array_obj_ref_740_store_0_ack_1 : boolean;
  signal array_obj_ref_756_gather_scatter_req_0 : boolean;
  signal array_obj_ref_756_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_756_store_0_req_0 : boolean;
  signal array_obj_ref_732_store_0_req_0 : boolean;
  signal array_obj_ref_732_store_0_ack_0 : boolean;
  signal array_obj_ref_740_store_0_req_0 : boolean;
  signal array_obj_ref_740_store_0_ack_0 : boolean;
  signal array_obj_ref_740_store_0_req_1 : boolean;
  signal array_obj_ref_752_store_0_ack_1 : boolean;
  signal array_obj_ref_740_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_752_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_752_store_0_req_0 : boolean;
  signal array_obj_ref_752_store_0_ack_0 : boolean;
  signal array_obj_ref_752_store_0_req_1 : boolean;
  signal array_obj_ref_740_gather_scatter_req_0 : boolean;
  signal array_obj_ref_752_gather_scatter_req_0 : boolean;
  signal array_obj_ref_732_gather_scatter_req_0 : boolean;
  signal array_obj_ref_732_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_748_store_0_req_0 : boolean;
  signal array_obj_ref_748_store_0_ack_0 : boolean;
  signal array_obj_ref_748_store_0_req_1 : boolean;
  signal array_obj_ref_748_store_0_ack_1 : boolean;
  signal array_obj_ref_768_gather_scatter_req_0 : boolean;
  signal array_obj_ref_768_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_720_store_0_req_1 : boolean;
  signal array_obj_ref_768_store_0_req_0 : boolean;
  signal array_obj_ref_768_store_0_ack_0 : boolean;
  signal array_obj_ref_768_store_0_req_1 : boolean;
  signal array_obj_ref_768_store_0_ack_1 : boolean;
  signal array_obj_ref_772_gather_scatter_req_0 : boolean;
  signal array_obj_ref_772_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_772_store_0_req_0 : boolean;
  signal array_obj_ref_772_store_0_ack_0 : boolean;
  signal array_obj_ref_772_store_0_req_1 : boolean;
  signal array_obj_ref_772_store_0_ack_1 : boolean;
  signal array_obj_ref_776_gather_scatter_req_0 : boolean;
  signal array_obj_ref_776_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_776_store_0_req_0 : boolean;
  signal array_obj_ref_776_store_0_ack_0 : boolean;
  signal array_obj_ref_776_store_0_req_1 : boolean;
  signal array_obj_ref_776_store_0_ack_1 : boolean;
  signal array_obj_ref_780_gather_scatter_req_0 : boolean;
  signal array_obj_ref_780_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_780_store_0_req_0 : boolean;
  signal array_obj_ref_780_store_0_ack_0 : boolean;
  signal array_obj_ref_780_store_0_req_1 : boolean;
  signal array_obj_ref_780_store_0_ack_1 : boolean;
  signal array_obj_ref_784_gather_scatter_req_0 : boolean;
  signal array_obj_ref_784_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_784_store_0_req_0 : boolean;
  signal array_obj_ref_784_store_0_ack_0 : boolean;
  signal array_obj_ref_784_store_0_req_1 : boolean;
  signal array_obj_ref_784_store_0_ack_1 : boolean;
  signal array_obj_ref_788_gather_scatter_req_0 : boolean;
  signal array_obj_ref_788_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_788_store_0_req_0 : boolean;
  signal array_obj_ref_788_store_0_ack_0 : boolean;
  signal array_obj_ref_788_store_0_req_1 : boolean;
  signal array_obj_ref_788_store_0_ack_1 : boolean;
  signal array_obj_ref_792_gather_scatter_req_0 : boolean;
  signal array_obj_ref_792_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_792_store_0_req_0 : boolean;
  signal array_obj_ref_792_store_0_ack_0 : boolean;
  signal array_obj_ref_792_store_0_req_1 : boolean;
  signal array_obj_ref_792_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 19 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr5_CP_3228: Block -- control-path 
    signal cp_elements: BooleanArray(57 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(57);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(57), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_720_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_720_gather_scatter_ack_0;
    array_obj_ref_720_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_720_store_0_ack_0;
    array_obj_ref_720_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_720_store_0_ack_1;
    array_obj_ref_724_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_724_gather_scatter_ack_0;
    array_obj_ref_724_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_724_store_0_ack_0;
    array_obj_ref_724_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_724_store_0_ack_1;
    array_obj_ref_728_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_728_gather_scatter_ack_0;
    array_obj_ref_728_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_728_store_0_ack_0;
    array_obj_ref_728_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_728_store_0_ack_1;
    array_obj_ref_732_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_732_gather_scatter_ack_0;
    array_obj_ref_732_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_732_store_0_ack_0;
    array_obj_ref_732_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_732_store_0_ack_1;
    array_obj_ref_736_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_736_gather_scatter_ack_0;
    array_obj_ref_736_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_736_store_0_ack_0;
    array_obj_ref_736_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_736_store_0_ack_1;
    array_obj_ref_740_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_740_gather_scatter_ack_0;
    array_obj_ref_740_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_740_store_0_ack_0;
    array_obj_ref_740_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_740_store_0_ack_1;
    array_obj_ref_744_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_744_gather_scatter_ack_0;
    array_obj_ref_744_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_744_store_0_ack_0;
    array_obj_ref_744_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_744_store_0_ack_1;
    array_obj_ref_748_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_748_gather_scatter_ack_0;
    array_obj_ref_748_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_748_store_0_ack_0;
    array_obj_ref_748_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_748_store_0_ack_1;
    array_obj_ref_752_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_752_gather_scatter_ack_0;
    array_obj_ref_752_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_752_store_0_ack_0;
    array_obj_ref_752_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_752_store_0_ack_1;
    array_obj_ref_756_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_756_gather_scatter_ack_0;
    array_obj_ref_756_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_756_store_0_ack_0;
    array_obj_ref_756_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_756_store_0_ack_1;
    array_obj_ref_760_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_760_gather_scatter_ack_0;
    array_obj_ref_760_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_760_store_0_ack_0;
    array_obj_ref_760_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_760_store_0_ack_1;
    array_obj_ref_764_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_764_gather_scatter_ack_0;
    array_obj_ref_764_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_764_store_0_ack_0;
    array_obj_ref_764_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_764_store_0_ack_1;
    array_obj_ref_768_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_768_gather_scatter_ack_0;
    array_obj_ref_768_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_768_store_0_ack_0;
    array_obj_ref_768_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_768_store_0_ack_1;
    array_obj_ref_772_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_772_gather_scatter_ack_0;
    array_obj_ref_772_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_772_store_0_ack_0;
    array_obj_ref_772_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_772_store_0_ack_1;
    array_obj_ref_776_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_776_gather_scatter_ack_0;
    array_obj_ref_776_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_776_store_0_ack_0;
    array_obj_ref_776_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_776_store_0_ack_1;
    array_obj_ref_780_gather_scatter_req_0 <= cp_elements(45);
    cp_elements(46) <= array_obj_ref_780_gather_scatter_ack_0;
    array_obj_ref_780_store_0_req_0 <= cp_elements(46);
    cp_elements(47) <= array_obj_ref_780_store_0_ack_0;
    array_obj_ref_780_store_0_req_1 <= cp_elements(47);
    cp_elements(48) <= array_obj_ref_780_store_0_ack_1;
    array_obj_ref_784_gather_scatter_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_784_gather_scatter_ack_0;
    array_obj_ref_784_store_0_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_784_store_0_ack_0;
    array_obj_ref_784_store_0_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_784_store_0_ack_1;
    array_obj_ref_788_gather_scatter_req_0 <= cp_elements(51);
    cp_elements(52) <= array_obj_ref_788_gather_scatter_ack_0;
    array_obj_ref_788_store_0_req_0 <= cp_elements(52);
    cp_elements(53) <= array_obj_ref_788_store_0_ack_0;
    array_obj_ref_788_store_0_req_1 <= cp_elements(53);
    cp_elements(54) <= array_obj_ref_788_store_0_ack_1;
    array_obj_ref_792_gather_scatter_req_0 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_792_gather_scatter_ack_0;
    array_obj_ref_792_store_0_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_792_store_0_ack_0;
    array_obj_ref_792_store_0_req_1 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_792_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_720_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_720_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_724_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_724_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_728_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_728_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_732_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_732_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_736_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_736_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_740_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_740_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_744_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_744_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_748_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_748_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_752_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_752_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_756_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_756_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_760_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_760_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_764_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_764_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_768_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_768_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_772_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_772_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_776_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_776_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_780_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_780_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_784_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_784_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_788_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_788_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_792_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_792_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_721_wire_constant : std_logic_vector(7 downto 0);
    signal expr_725_wire_constant : std_logic_vector(7 downto 0);
    signal expr_729_wire_constant : std_logic_vector(7 downto 0);
    signal expr_733_wire_constant : std_logic_vector(7 downto 0);
    signal expr_737_wire_constant : std_logic_vector(7 downto 0);
    signal expr_741_wire_constant : std_logic_vector(7 downto 0);
    signal expr_745_wire_constant : std_logic_vector(7 downto 0);
    signal expr_749_wire_constant : std_logic_vector(7 downto 0);
    signal expr_753_wire_constant : std_logic_vector(7 downto 0);
    signal expr_757_wire_constant : std_logic_vector(7 downto 0);
    signal expr_761_wire_constant : std_logic_vector(7 downto 0);
    signal expr_765_wire_constant : std_logic_vector(7 downto 0);
    signal expr_769_wire_constant : std_logic_vector(7 downto 0);
    signal expr_773_wire_constant : std_logic_vector(7 downto 0);
    signal expr_777_wire_constant : std_logic_vector(7 downto 0);
    signal expr_781_wire_constant : std_logic_vector(7 downto 0);
    signal expr_785_wire_constant : std_logic_vector(7 downto 0);
    signal expr_789_wire_constant : std_logic_vector(7 downto 0);
    signal expr_793_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_720_word_address_0 <= "00000";
    array_obj_ref_724_word_address_0 <= "00001";
    array_obj_ref_728_word_address_0 <= "00010";
    array_obj_ref_732_word_address_0 <= "00011";
    array_obj_ref_736_word_address_0 <= "00100";
    array_obj_ref_740_word_address_0 <= "00101";
    array_obj_ref_744_word_address_0 <= "00110";
    array_obj_ref_748_word_address_0 <= "00111";
    array_obj_ref_752_word_address_0 <= "01000";
    array_obj_ref_756_word_address_0 <= "01001";
    array_obj_ref_760_word_address_0 <= "01010";
    array_obj_ref_764_word_address_0 <= "01011";
    array_obj_ref_768_word_address_0 <= "01100";
    array_obj_ref_772_word_address_0 <= "01101";
    array_obj_ref_776_word_address_0 <= "01110";
    array_obj_ref_780_word_address_0 <= "01111";
    array_obj_ref_784_word_address_0 <= "10000";
    array_obj_ref_788_word_address_0 <= "10001";
    array_obj_ref_792_word_address_0 <= "10010";
    expr_721_wire_constant <= "01100110";
    expr_725_wire_constant <= "01110010";
    expr_729_wire_constant <= "01100101";
    expr_733_wire_constant <= "01100101";
    expr_737_wire_constant <= "01011111";
    expr_741_wire_constant <= "01110001";
    expr_745_wire_constant <= "01110101";
    expr_749_wire_constant <= "01100101";
    expr_753_wire_constant <= "01110101";
    expr_757_wire_constant <= "01100101";
    expr_761_wire_constant <= "01011111";
    expr_765_wire_constant <= "01110010";
    expr_769_wire_constant <= "01100101";
    expr_773_wire_constant <= "01110001";
    expr_777_wire_constant <= "01110101";
    expr_781_wire_constant <= "01100101";
    expr_785_wire_constant <= "01110011";
    expr_789_wire_constant <= "01110100";
    expr_793_wire_constant <= "00000000";
    array_obj_ref_720_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_720_gather_scatter_ack_0 <= array_obj_ref_720_gather_scatter_req_0;
      aggregated_sig <= expr_721_wire_constant;
      array_obj_ref_720_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_724_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_724_gather_scatter_ack_0 <= array_obj_ref_724_gather_scatter_req_0;
      aggregated_sig <= expr_725_wire_constant;
      array_obj_ref_724_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_728_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_728_gather_scatter_ack_0 <= array_obj_ref_728_gather_scatter_req_0;
      aggregated_sig <= expr_729_wire_constant;
      array_obj_ref_728_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_732_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_732_gather_scatter_ack_0 <= array_obj_ref_732_gather_scatter_req_0;
      aggregated_sig <= expr_733_wire_constant;
      array_obj_ref_732_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_736_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_736_gather_scatter_ack_0 <= array_obj_ref_736_gather_scatter_req_0;
      aggregated_sig <= expr_737_wire_constant;
      array_obj_ref_736_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_740_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_740_gather_scatter_ack_0 <= array_obj_ref_740_gather_scatter_req_0;
      aggregated_sig <= expr_741_wire_constant;
      array_obj_ref_740_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_744_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_744_gather_scatter_ack_0 <= array_obj_ref_744_gather_scatter_req_0;
      aggregated_sig <= expr_745_wire_constant;
      array_obj_ref_744_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_748_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_748_gather_scatter_ack_0 <= array_obj_ref_748_gather_scatter_req_0;
      aggregated_sig <= expr_749_wire_constant;
      array_obj_ref_748_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_752_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_752_gather_scatter_ack_0 <= array_obj_ref_752_gather_scatter_req_0;
      aggregated_sig <= expr_753_wire_constant;
      array_obj_ref_752_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_756_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_756_gather_scatter_ack_0 <= array_obj_ref_756_gather_scatter_req_0;
      aggregated_sig <= expr_757_wire_constant;
      array_obj_ref_756_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_760_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_760_gather_scatter_ack_0 <= array_obj_ref_760_gather_scatter_req_0;
      aggregated_sig <= expr_761_wire_constant;
      array_obj_ref_760_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_764_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_764_gather_scatter_ack_0 <= array_obj_ref_764_gather_scatter_req_0;
      aggregated_sig <= expr_765_wire_constant;
      array_obj_ref_764_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_768_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_768_gather_scatter_ack_0 <= array_obj_ref_768_gather_scatter_req_0;
      aggregated_sig <= expr_769_wire_constant;
      array_obj_ref_768_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_772_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_772_gather_scatter_ack_0 <= array_obj_ref_772_gather_scatter_req_0;
      aggregated_sig <= expr_773_wire_constant;
      array_obj_ref_772_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_776_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_776_gather_scatter_ack_0 <= array_obj_ref_776_gather_scatter_req_0;
      aggregated_sig <= expr_777_wire_constant;
      array_obj_ref_776_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_780_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_780_gather_scatter_ack_0 <= array_obj_ref_780_gather_scatter_req_0;
      aggregated_sig <= expr_781_wire_constant;
      array_obj_ref_780_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_784_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_784_gather_scatter_ack_0 <= array_obj_ref_784_gather_scatter_req_0;
      aggregated_sig <= expr_785_wire_constant;
      array_obj_ref_784_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_788_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_788_gather_scatter_ack_0 <= array_obj_ref_788_gather_scatter_req_0;
      aggregated_sig <= expr_789_wire_constant;
      array_obj_ref_788_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_792_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_792_gather_scatter_ack_0 <= array_obj_ref_792_gather_scatter_req_0;
      aggregated_sig <= expr_793_wire_constant;
      array_obj_ref_792_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_720_store_0 array_obj_ref_724_store_0 array_obj_ref_728_store_0 array_obj_ref_732_store_0 array_obj_ref_736_store_0 array_obj_ref_740_store_0 array_obj_ref_744_store_0 array_obj_ref_748_store_0 array_obj_ref_752_store_0 array_obj_ref_756_store_0 array_obj_ref_760_store_0 array_obj_ref_764_store_0 array_obj_ref_768_store_0 array_obj_ref_772_store_0 array_obj_ref_776_store_0 array_obj_ref_780_store_0 array_obj_ref_784_store_0 array_obj_ref_788_store_0 array_obj_ref_792_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(94 downto 0);
      signal data_in: std_logic_vector(151 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 18 downto 0);
      -- 
    begin -- 
      reqL(18) <= array_obj_ref_720_store_0_req_0;
      reqL(17) <= array_obj_ref_724_store_0_req_0;
      reqL(16) <= array_obj_ref_728_store_0_req_0;
      reqL(15) <= array_obj_ref_732_store_0_req_0;
      reqL(14) <= array_obj_ref_736_store_0_req_0;
      reqL(13) <= array_obj_ref_740_store_0_req_0;
      reqL(12) <= array_obj_ref_744_store_0_req_0;
      reqL(11) <= array_obj_ref_748_store_0_req_0;
      reqL(10) <= array_obj_ref_752_store_0_req_0;
      reqL(9) <= array_obj_ref_756_store_0_req_0;
      reqL(8) <= array_obj_ref_760_store_0_req_0;
      reqL(7) <= array_obj_ref_764_store_0_req_0;
      reqL(6) <= array_obj_ref_768_store_0_req_0;
      reqL(5) <= array_obj_ref_772_store_0_req_0;
      reqL(4) <= array_obj_ref_776_store_0_req_0;
      reqL(3) <= array_obj_ref_780_store_0_req_0;
      reqL(2) <= array_obj_ref_784_store_0_req_0;
      reqL(1) <= array_obj_ref_788_store_0_req_0;
      reqL(0) <= array_obj_ref_792_store_0_req_0;
      array_obj_ref_720_store_0_ack_0 <= ackL(18);
      array_obj_ref_724_store_0_ack_0 <= ackL(17);
      array_obj_ref_728_store_0_ack_0 <= ackL(16);
      array_obj_ref_732_store_0_ack_0 <= ackL(15);
      array_obj_ref_736_store_0_ack_0 <= ackL(14);
      array_obj_ref_740_store_0_ack_0 <= ackL(13);
      array_obj_ref_744_store_0_ack_0 <= ackL(12);
      array_obj_ref_748_store_0_ack_0 <= ackL(11);
      array_obj_ref_752_store_0_ack_0 <= ackL(10);
      array_obj_ref_756_store_0_ack_0 <= ackL(9);
      array_obj_ref_760_store_0_ack_0 <= ackL(8);
      array_obj_ref_764_store_0_ack_0 <= ackL(7);
      array_obj_ref_768_store_0_ack_0 <= ackL(6);
      array_obj_ref_772_store_0_ack_0 <= ackL(5);
      array_obj_ref_776_store_0_ack_0 <= ackL(4);
      array_obj_ref_780_store_0_ack_0 <= ackL(3);
      array_obj_ref_784_store_0_ack_0 <= ackL(2);
      array_obj_ref_788_store_0_ack_0 <= ackL(1);
      array_obj_ref_792_store_0_ack_0 <= ackL(0);
      reqR(18) <= array_obj_ref_720_store_0_req_1;
      reqR(17) <= array_obj_ref_724_store_0_req_1;
      reqR(16) <= array_obj_ref_728_store_0_req_1;
      reqR(15) <= array_obj_ref_732_store_0_req_1;
      reqR(14) <= array_obj_ref_736_store_0_req_1;
      reqR(13) <= array_obj_ref_740_store_0_req_1;
      reqR(12) <= array_obj_ref_744_store_0_req_1;
      reqR(11) <= array_obj_ref_748_store_0_req_1;
      reqR(10) <= array_obj_ref_752_store_0_req_1;
      reqR(9) <= array_obj_ref_756_store_0_req_1;
      reqR(8) <= array_obj_ref_760_store_0_req_1;
      reqR(7) <= array_obj_ref_764_store_0_req_1;
      reqR(6) <= array_obj_ref_768_store_0_req_1;
      reqR(5) <= array_obj_ref_772_store_0_req_1;
      reqR(4) <= array_obj_ref_776_store_0_req_1;
      reqR(3) <= array_obj_ref_780_store_0_req_1;
      reqR(2) <= array_obj_ref_784_store_0_req_1;
      reqR(1) <= array_obj_ref_788_store_0_req_1;
      reqR(0) <= array_obj_ref_792_store_0_req_1;
      array_obj_ref_720_store_0_ack_1 <= ackR(18);
      array_obj_ref_724_store_0_ack_1 <= ackR(17);
      array_obj_ref_728_store_0_ack_1 <= ackR(16);
      array_obj_ref_732_store_0_ack_1 <= ackR(15);
      array_obj_ref_736_store_0_ack_1 <= ackR(14);
      array_obj_ref_740_store_0_ack_1 <= ackR(13);
      array_obj_ref_744_store_0_ack_1 <= ackR(12);
      array_obj_ref_748_store_0_ack_1 <= ackR(11);
      array_obj_ref_752_store_0_ack_1 <= ackR(10);
      array_obj_ref_756_store_0_ack_1 <= ackR(9);
      array_obj_ref_760_store_0_ack_1 <= ackR(8);
      array_obj_ref_764_store_0_ack_1 <= ackR(7);
      array_obj_ref_768_store_0_ack_1 <= ackR(6);
      array_obj_ref_772_store_0_ack_1 <= ackR(5);
      array_obj_ref_776_store_0_ack_1 <= ackR(4);
      array_obj_ref_780_store_0_ack_1 <= ackR(3);
      array_obj_ref_784_store_0_ack_1 <= ackR(2);
      array_obj_ref_788_store_0_ack_1 <= ackR(1);
      array_obj_ref_792_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_720_word_address_0 & array_obj_ref_724_word_address_0 & array_obj_ref_728_word_address_0 & array_obj_ref_732_word_address_0 & array_obj_ref_736_word_address_0 & array_obj_ref_740_word_address_0 & array_obj_ref_744_word_address_0 & array_obj_ref_748_word_address_0 & array_obj_ref_752_word_address_0 & array_obj_ref_756_word_address_0 & array_obj_ref_760_word_address_0 & array_obj_ref_764_word_address_0 & array_obj_ref_768_word_address_0 & array_obj_ref_772_word_address_0 & array_obj_ref_776_word_address_0 & array_obj_ref_780_word_address_0 & array_obj_ref_784_word_address_0 & array_obj_ref_788_word_address_0 & array_obj_ref_792_word_address_0;
      data_in <= array_obj_ref_720_data_0 & array_obj_ref_724_data_0 & array_obj_ref_728_data_0 & array_obj_ref_732_data_0 & array_obj_ref_736_data_0 & array_obj_ref_740_data_0 & array_obj_ref_744_data_0 & array_obj_ref_748_data_0 & array_obj_ref_752_data_0 & array_obj_ref_756_data_0 & array_obj_ref_760_data_0 & array_obj_ref_764_data_0 & array_obj_ref_768_data_0 & array_obj_ref_772_data_0 & array_obj_ref_776_data_0 & array_obj_ref_780_data_0 & array_obj_ref_784_data_0 & array_obj_ref_788_data_0 & array_obj_ref_792_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 8,
        num_reqs => 19,
        tag_length => 5,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_15_sr_req(0),
          mack => memory_space_15_sr_ack(0),
          maddr => memory_space_15_sr_addr(4 downto 0),
          mdata => memory_space_15_sr_data(7 downto 0),
          mtag => memory_space_15_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 19,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_15_sc_req(0),
          mack => memory_space_15_sc_ack(0),
          mtag => memory_space_15_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr6 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_16_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_16_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_16_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_16_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_16_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_16_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_16_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_16_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr6;
architecture Default of default_initializer_xx_xstr6 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr6_CP_3630_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_798_gather_scatter_req_0 : boolean;
  signal array_obj_ref_798_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_798_store_0_req_0 : boolean;
  signal array_obj_ref_798_store_0_ack_0 : boolean;
  signal array_obj_ref_798_store_0_req_1 : boolean;
  signal array_obj_ref_798_store_0_ack_1 : boolean;
  signal array_obj_ref_802_gather_scatter_req_0 : boolean;
  signal array_obj_ref_802_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_802_store_0_req_0 : boolean;
  signal array_obj_ref_802_store_0_ack_0 : boolean;
  signal array_obj_ref_802_store_0_req_1 : boolean;
  signal array_obj_ref_802_store_0_ack_1 : boolean;
  signal array_obj_ref_806_gather_scatter_req_0 : boolean;
  signal array_obj_ref_806_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_806_store_0_req_0 : boolean;
  signal array_obj_ref_806_store_0_ack_0 : boolean;
  signal array_obj_ref_806_store_0_req_1 : boolean;
  signal array_obj_ref_806_store_0_ack_1 : boolean;
  signal array_obj_ref_810_gather_scatter_req_0 : boolean;
  signal array_obj_ref_810_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_810_store_0_req_0 : boolean;
  signal array_obj_ref_810_store_0_ack_0 : boolean;
  signal array_obj_ref_810_store_0_req_1 : boolean;
  signal array_obj_ref_810_store_0_ack_1 : boolean;
  signal array_obj_ref_814_gather_scatter_req_0 : boolean;
  signal array_obj_ref_814_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_814_store_0_req_0 : boolean;
  signal array_obj_ref_814_store_0_ack_0 : boolean;
  signal array_obj_ref_814_store_0_req_1 : boolean;
  signal array_obj_ref_814_store_0_ack_1 : boolean;
  signal array_obj_ref_818_gather_scatter_req_0 : boolean;
  signal array_obj_ref_818_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_818_store_0_req_0 : boolean;
  signal array_obj_ref_818_store_0_ack_0 : boolean;
  signal array_obj_ref_818_store_0_req_1 : boolean;
  signal array_obj_ref_818_store_0_ack_1 : boolean;
  signal array_obj_ref_822_gather_scatter_req_0 : boolean;
  signal array_obj_ref_822_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_822_store_0_req_0 : boolean;
  signal array_obj_ref_822_store_0_ack_0 : boolean;
  signal array_obj_ref_822_store_0_req_1 : boolean;
  signal array_obj_ref_822_store_0_ack_1 : boolean;
  signal array_obj_ref_826_gather_scatter_req_0 : boolean;
  signal array_obj_ref_826_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_826_store_0_req_0 : boolean;
  signal array_obj_ref_826_store_0_ack_0 : boolean;
  signal array_obj_ref_826_store_0_req_1 : boolean;
  signal array_obj_ref_826_store_0_ack_1 : boolean;
  signal array_obj_ref_830_gather_scatter_req_0 : boolean;
  signal array_obj_ref_830_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_830_store_0_req_0 : boolean;
  signal array_obj_ref_830_store_0_ack_0 : boolean;
  signal array_obj_ref_830_store_0_req_1 : boolean;
  signal array_obj_ref_830_store_0_ack_1 : boolean;
  signal array_obj_ref_834_gather_scatter_req_0 : boolean;
  signal array_obj_ref_834_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_834_store_0_req_0 : boolean;
  signal array_obj_ref_834_store_0_ack_0 : boolean;
  signal array_obj_ref_834_store_0_req_1 : boolean;
  signal array_obj_ref_834_store_0_ack_1 : boolean;
  signal array_obj_ref_838_gather_scatter_req_0 : boolean;
  signal array_obj_ref_838_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_838_store_0_req_0 : boolean;
  signal array_obj_ref_838_store_0_ack_0 : boolean;
  signal array_obj_ref_838_store_0_req_1 : boolean;
  signal array_obj_ref_838_store_0_ack_1 : boolean;
  signal array_obj_ref_842_gather_scatter_req_0 : boolean;
  signal array_obj_ref_842_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_842_store_0_req_0 : boolean;
  signal array_obj_ref_842_store_0_ack_0 : boolean;
  signal array_obj_ref_842_store_0_req_1 : boolean;
  signal array_obj_ref_842_store_0_ack_1 : boolean;
  signal array_obj_ref_846_gather_scatter_req_0 : boolean;
  signal array_obj_ref_846_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_846_store_0_req_0 : boolean;
  signal array_obj_ref_846_store_0_ack_0 : boolean;
  signal array_obj_ref_846_store_0_req_1 : boolean;
  signal array_obj_ref_846_store_0_ack_1 : boolean;
  signal array_obj_ref_850_gather_scatter_req_0 : boolean;
  signal array_obj_ref_850_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_850_store_0_req_0 : boolean;
  signal array_obj_ref_850_store_0_ack_0 : boolean;
  signal array_obj_ref_850_store_0_req_1 : boolean;
  signal array_obj_ref_850_store_0_ack_1 : boolean;
  signal array_obj_ref_854_gather_scatter_req_0 : boolean;
  signal array_obj_ref_854_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_854_store_0_req_0 : boolean;
  signal array_obj_ref_854_store_0_ack_0 : boolean;
  signal array_obj_ref_854_store_0_req_1 : boolean;
  signal array_obj_ref_854_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 15 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr6_CP_3630: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_798_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_798_gather_scatter_ack_0;
    array_obj_ref_798_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_798_store_0_ack_0;
    array_obj_ref_798_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_798_store_0_ack_1;
    array_obj_ref_802_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_802_gather_scatter_ack_0;
    array_obj_ref_802_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_802_store_0_ack_0;
    array_obj_ref_802_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_802_store_0_ack_1;
    array_obj_ref_806_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_806_gather_scatter_ack_0;
    array_obj_ref_806_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_806_store_0_ack_0;
    array_obj_ref_806_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_806_store_0_ack_1;
    array_obj_ref_810_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_810_gather_scatter_ack_0;
    array_obj_ref_810_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_810_store_0_ack_0;
    array_obj_ref_810_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_810_store_0_ack_1;
    array_obj_ref_814_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_814_gather_scatter_ack_0;
    array_obj_ref_814_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_814_store_0_ack_0;
    array_obj_ref_814_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_814_store_0_ack_1;
    array_obj_ref_818_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_818_gather_scatter_ack_0;
    array_obj_ref_818_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_818_store_0_ack_0;
    array_obj_ref_818_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_818_store_0_ack_1;
    array_obj_ref_822_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_822_gather_scatter_ack_0;
    array_obj_ref_822_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_822_store_0_ack_0;
    array_obj_ref_822_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_822_store_0_ack_1;
    array_obj_ref_826_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_826_gather_scatter_ack_0;
    array_obj_ref_826_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_826_store_0_ack_0;
    array_obj_ref_826_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_826_store_0_ack_1;
    array_obj_ref_830_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_830_gather_scatter_ack_0;
    array_obj_ref_830_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_830_store_0_ack_0;
    array_obj_ref_830_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_830_store_0_ack_1;
    array_obj_ref_834_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_834_gather_scatter_ack_0;
    array_obj_ref_834_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_834_store_0_ack_0;
    array_obj_ref_834_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_834_store_0_ack_1;
    array_obj_ref_838_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_838_gather_scatter_ack_0;
    array_obj_ref_838_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_838_store_0_ack_0;
    array_obj_ref_838_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_838_store_0_ack_1;
    array_obj_ref_842_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_842_gather_scatter_ack_0;
    array_obj_ref_842_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_842_store_0_ack_0;
    array_obj_ref_842_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_842_store_0_ack_1;
    array_obj_ref_846_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_846_gather_scatter_ack_0;
    array_obj_ref_846_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_846_store_0_ack_0;
    array_obj_ref_846_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_846_store_0_ack_1;
    array_obj_ref_850_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_850_gather_scatter_ack_0;
    array_obj_ref_850_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_850_store_0_ack_0;
    array_obj_ref_850_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_850_store_0_ack_1;
    array_obj_ref_854_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_854_gather_scatter_ack_0;
    array_obj_ref_854_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_854_store_0_ack_0;
    array_obj_ref_854_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_854_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_798_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_798_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_802_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_802_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_806_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_806_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_810_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_810_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_814_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_814_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_818_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_822_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_822_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_826_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_826_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_830_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_830_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_834_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_834_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_838_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_838_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_842_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_842_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_846_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_846_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_850_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_850_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_854_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_854_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_799_wire_constant : std_logic_vector(7 downto 0);
    signal expr_803_wire_constant : std_logic_vector(7 downto 0);
    signal expr_807_wire_constant : std_logic_vector(7 downto 0);
    signal expr_811_wire_constant : std_logic_vector(7 downto 0);
    signal expr_815_wire_constant : std_logic_vector(7 downto 0);
    signal expr_819_wire_constant : std_logic_vector(7 downto 0);
    signal expr_823_wire_constant : std_logic_vector(7 downto 0);
    signal expr_827_wire_constant : std_logic_vector(7 downto 0);
    signal expr_831_wire_constant : std_logic_vector(7 downto 0);
    signal expr_835_wire_constant : std_logic_vector(7 downto 0);
    signal expr_839_wire_constant : std_logic_vector(7 downto 0);
    signal expr_843_wire_constant : std_logic_vector(7 downto 0);
    signal expr_847_wire_constant : std_logic_vector(7 downto 0);
    signal expr_851_wire_constant : std_logic_vector(7 downto 0);
    signal expr_855_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_798_word_address_0 <= "0000";
    array_obj_ref_802_word_address_0 <= "0001";
    array_obj_ref_806_word_address_0 <= "0010";
    array_obj_ref_810_word_address_0 <= "0011";
    array_obj_ref_814_word_address_0 <= "0100";
    array_obj_ref_818_word_address_0 <= "0101";
    array_obj_ref_822_word_address_0 <= "0110";
    array_obj_ref_826_word_address_0 <= "0111";
    array_obj_ref_830_word_address_0 <= "1000";
    array_obj_ref_834_word_address_0 <= "1001";
    array_obj_ref_838_word_address_0 <= "1010";
    array_obj_ref_842_word_address_0 <= "1011";
    array_obj_ref_846_word_address_0 <= "1100";
    array_obj_ref_850_word_address_0 <= "1101";
    array_obj_ref_854_word_address_0 <= "1110";
    expr_799_wire_constant <= "01100110";
    expr_803_wire_constant <= "01110010";
    expr_807_wire_constant <= "01100101";
    expr_811_wire_constant <= "01100101";
    expr_815_wire_constant <= "01011111";
    expr_819_wire_constant <= "01110001";
    expr_823_wire_constant <= "01110101";
    expr_827_wire_constant <= "01100101";
    expr_831_wire_constant <= "01110101";
    expr_835_wire_constant <= "01100101";
    expr_839_wire_constant <= "01011111";
    expr_843_wire_constant <= "01100001";
    expr_847_wire_constant <= "01100011";
    expr_851_wire_constant <= "01101011";
    expr_855_wire_constant <= "00000000";
    array_obj_ref_798_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_798_gather_scatter_ack_0 <= array_obj_ref_798_gather_scatter_req_0;
      aggregated_sig <= expr_799_wire_constant;
      array_obj_ref_798_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_802_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_802_gather_scatter_ack_0 <= array_obj_ref_802_gather_scatter_req_0;
      aggregated_sig <= expr_803_wire_constant;
      array_obj_ref_802_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_806_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_806_gather_scatter_ack_0 <= array_obj_ref_806_gather_scatter_req_0;
      aggregated_sig <= expr_807_wire_constant;
      array_obj_ref_806_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_810_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_810_gather_scatter_ack_0 <= array_obj_ref_810_gather_scatter_req_0;
      aggregated_sig <= expr_811_wire_constant;
      array_obj_ref_810_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_814_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_814_gather_scatter_ack_0 <= array_obj_ref_814_gather_scatter_req_0;
      aggregated_sig <= expr_815_wire_constant;
      array_obj_ref_814_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_818_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_818_gather_scatter_ack_0 <= array_obj_ref_818_gather_scatter_req_0;
      aggregated_sig <= expr_819_wire_constant;
      array_obj_ref_818_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_822_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_822_gather_scatter_ack_0 <= array_obj_ref_822_gather_scatter_req_0;
      aggregated_sig <= expr_823_wire_constant;
      array_obj_ref_822_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_826_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_826_gather_scatter_ack_0 <= array_obj_ref_826_gather_scatter_req_0;
      aggregated_sig <= expr_827_wire_constant;
      array_obj_ref_826_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_830_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_830_gather_scatter_ack_0 <= array_obj_ref_830_gather_scatter_req_0;
      aggregated_sig <= expr_831_wire_constant;
      array_obj_ref_830_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_834_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_834_gather_scatter_ack_0 <= array_obj_ref_834_gather_scatter_req_0;
      aggregated_sig <= expr_835_wire_constant;
      array_obj_ref_834_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_838_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_838_gather_scatter_ack_0 <= array_obj_ref_838_gather_scatter_req_0;
      aggregated_sig <= expr_839_wire_constant;
      array_obj_ref_838_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_842_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_842_gather_scatter_ack_0 <= array_obj_ref_842_gather_scatter_req_0;
      aggregated_sig <= expr_843_wire_constant;
      array_obj_ref_842_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_846_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_846_gather_scatter_ack_0 <= array_obj_ref_846_gather_scatter_req_0;
      aggregated_sig <= expr_847_wire_constant;
      array_obj_ref_846_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_850_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_850_gather_scatter_ack_0 <= array_obj_ref_850_gather_scatter_req_0;
      aggregated_sig <= expr_851_wire_constant;
      array_obj_ref_850_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_854_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_854_gather_scatter_ack_0 <= array_obj_ref_854_gather_scatter_req_0;
      aggregated_sig <= expr_855_wire_constant;
      array_obj_ref_854_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_826_store_0 array_obj_ref_838_store_0 array_obj_ref_830_store_0 array_obj_ref_802_store_0 array_obj_ref_850_store_0 array_obj_ref_814_store_0 array_obj_ref_842_store_0 array_obj_ref_846_store_0 array_obj_ref_834_store_0 array_obj_ref_854_store_0 array_obj_ref_822_store_0 array_obj_ref_798_store_0 array_obj_ref_810_store_0 array_obj_ref_818_store_0 array_obj_ref_806_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(59 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_826_store_0_req_0;
      reqL(13) <= array_obj_ref_838_store_0_req_0;
      reqL(12) <= array_obj_ref_830_store_0_req_0;
      reqL(11) <= array_obj_ref_802_store_0_req_0;
      reqL(10) <= array_obj_ref_850_store_0_req_0;
      reqL(9) <= array_obj_ref_814_store_0_req_0;
      reqL(8) <= array_obj_ref_842_store_0_req_0;
      reqL(7) <= array_obj_ref_846_store_0_req_0;
      reqL(6) <= array_obj_ref_834_store_0_req_0;
      reqL(5) <= array_obj_ref_854_store_0_req_0;
      reqL(4) <= array_obj_ref_822_store_0_req_0;
      reqL(3) <= array_obj_ref_798_store_0_req_0;
      reqL(2) <= array_obj_ref_810_store_0_req_0;
      reqL(1) <= array_obj_ref_818_store_0_req_0;
      reqL(0) <= array_obj_ref_806_store_0_req_0;
      array_obj_ref_826_store_0_ack_0 <= ackL(14);
      array_obj_ref_838_store_0_ack_0 <= ackL(13);
      array_obj_ref_830_store_0_ack_0 <= ackL(12);
      array_obj_ref_802_store_0_ack_0 <= ackL(11);
      array_obj_ref_850_store_0_ack_0 <= ackL(10);
      array_obj_ref_814_store_0_ack_0 <= ackL(9);
      array_obj_ref_842_store_0_ack_0 <= ackL(8);
      array_obj_ref_846_store_0_ack_0 <= ackL(7);
      array_obj_ref_834_store_0_ack_0 <= ackL(6);
      array_obj_ref_854_store_0_ack_0 <= ackL(5);
      array_obj_ref_822_store_0_ack_0 <= ackL(4);
      array_obj_ref_798_store_0_ack_0 <= ackL(3);
      array_obj_ref_810_store_0_ack_0 <= ackL(2);
      array_obj_ref_818_store_0_ack_0 <= ackL(1);
      array_obj_ref_806_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_826_store_0_req_1;
      reqR(13) <= array_obj_ref_838_store_0_req_1;
      reqR(12) <= array_obj_ref_830_store_0_req_1;
      reqR(11) <= array_obj_ref_802_store_0_req_1;
      reqR(10) <= array_obj_ref_850_store_0_req_1;
      reqR(9) <= array_obj_ref_814_store_0_req_1;
      reqR(8) <= array_obj_ref_842_store_0_req_1;
      reqR(7) <= array_obj_ref_846_store_0_req_1;
      reqR(6) <= array_obj_ref_834_store_0_req_1;
      reqR(5) <= array_obj_ref_854_store_0_req_1;
      reqR(4) <= array_obj_ref_822_store_0_req_1;
      reqR(3) <= array_obj_ref_798_store_0_req_1;
      reqR(2) <= array_obj_ref_810_store_0_req_1;
      reqR(1) <= array_obj_ref_818_store_0_req_1;
      reqR(0) <= array_obj_ref_806_store_0_req_1;
      array_obj_ref_826_store_0_ack_1 <= ackR(14);
      array_obj_ref_838_store_0_ack_1 <= ackR(13);
      array_obj_ref_830_store_0_ack_1 <= ackR(12);
      array_obj_ref_802_store_0_ack_1 <= ackR(11);
      array_obj_ref_850_store_0_ack_1 <= ackR(10);
      array_obj_ref_814_store_0_ack_1 <= ackR(9);
      array_obj_ref_842_store_0_ack_1 <= ackR(8);
      array_obj_ref_846_store_0_ack_1 <= ackR(7);
      array_obj_ref_834_store_0_ack_1 <= ackR(6);
      array_obj_ref_854_store_0_ack_1 <= ackR(5);
      array_obj_ref_822_store_0_ack_1 <= ackR(4);
      array_obj_ref_798_store_0_ack_1 <= ackR(3);
      array_obj_ref_810_store_0_ack_1 <= ackR(2);
      array_obj_ref_818_store_0_ack_1 <= ackR(1);
      array_obj_ref_806_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_826_word_address_0 & array_obj_ref_838_word_address_0 & array_obj_ref_830_word_address_0 & array_obj_ref_802_word_address_0 & array_obj_ref_850_word_address_0 & array_obj_ref_814_word_address_0 & array_obj_ref_842_word_address_0 & array_obj_ref_846_word_address_0 & array_obj_ref_834_word_address_0 & array_obj_ref_854_word_address_0 & array_obj_ref_822_word_address_0 & array_obj_ref_798_word_address_0 & array_obj_ref_810_word_address_0 & array_obj_ref_818_word_address_0 & array_obj_ref_806_word_address_0;
      data_in <= array_obj_ref_826_data_0 & array_obj_ref_838_data_0 & array_obj_ref_830_data_0 & array_obj_ref_802_data_0 & array_obj_ref_850_data_0 & array_obj_ref_814_data_0 & array_obj_ref_842_data_0 & array_obj_ref_846_data_0 & array_obj_ref_834_data_0 & array_obj_ref_854_data_0 & array_obj_ref_822_data_0 & array_obj_ref_798_data_0 & array_obj_ref_810_data_0 & array_obj_ref_818_data_0 & array_obj_ref_806_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 15,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_16_sr_req(0),
          mack => memory_space_16_sr_ack(0),
          maddr => memory_space_16_sr_addr(3 downto 0),
          mdata => memory_space_16_sr_data(7 downto 0),
          mtag => memory_space_16_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_16_sc_req(0),
          mack => memory_space_16_sc_ack(0),
          mtag => memory_space_16_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr7 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_17_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_17_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_17_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_17_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_17_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_17_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_17_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_17_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr7;
architecture Default of default_initializer_xx_xstr7 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr7_CP_3948_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_860_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_864_store_0_ack_0 : boolean;
  signal array_obj_ref_864_gather_scatter_req_0 : boolean;
  signal array_obj_ref_864_store_0_req_1 : boolean;
  signal array_obj_ref_864_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_860_gather_scatter_req_0 : boolean;
  signal array_obj_ref_860_store_0_req_1 : boolean;
  signal array_obj_ref_860_store_0_ack_0 : boolean;
  signal array_obj_ref_864_store_0_req_0 : boolean;
  signal array_obj_ref_860_store_0_req_0 : boolean;
  signal array_obj_ref_864_store_0_ack_1 : boolean;
  signal array_obj_ref_868_gather_scatter_req_0 : boolean;
  signal array_obj_ref_860_store_0_ack_1 : boolean;
  signal array_obj_ref_868_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_868_store_0_req_0 : boolean;
  signal array_obj_ref_868_store_0_ack_0 : boolean;
  signal array_obj_ref_868_store_0_req_1 : boolean;
  signal array_obj_ref_868_store_0_ack_1 : boolean;
  signal array_obj_ref_872_gather_scatter_req_0 : boolean;
  signal array_obj_ref_872_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_872_store_0_req_0 : boolean;
  signal array_obj_ref_872_store_0_ack_0 : boolean;
  signal array_obj_ref_872_store_0_req_1 : boolean;
  signal array_obj_ref_872_store_0_ack_1 : boolean;
  signal array_obj_ref_876_gather_scatter_req_0 : boolean;
  signal array_obj_ref_876_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_876_store_0_req_0 : boolean;
  signal array_obj_ref_876_store_0_ack_0 : boolean;
  signal array_obj_ref_876_store_0_req_1 : boolean;
  signal array_obj_ref_876_store_0_ack_1 : boolean;
  signal array_obj_ref_880_gather_scatter_req_0 : boolean;
  signal array_obj_ref_880_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_880_store_0_req_0 : boolean;
  signal array_obj_ref_880_store_0_ack_0 : boolean;
  signal array_obj_ref_880_store_0_req_1 : boolean;
  signal array_obj_ref_880_store_0_ack_1 : boolean;
  signal array_obj_ref_884_gather_scatter_req_0 : boolean;
  signal array_obj_ref_884_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_884_store_0_req_0 : boolean;
  signal array_obj_ref_884_store_0_ack_0 : boolean;
  signal array_obj_ref_884_store_0_req_1 : boolean;
  signal array_obj_ref_884_store_0_ack_1 : boolean;
  signal array_obj_ref_888_gather_scatter_req_0 : boolean;
  signal array_obj_ref_888_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_888_store_0_req_0 : boolean;
  signal array_obj_ref_888_store_0_ack_0 : boolean;
  signal array_obj_ref_888_store_0_req_1 : boolean;
  signal array_obj_ref_888_store_0_ack_1 : boolean;
  signal array_obj_ref_892_gather_scatter_req_0 : boolean;
  signal array_obj_ref_892_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_892_store_0_req_0 : boolean;
  signal array_obj_ref_892_store_0_ack_0 : boolean;
  signal array_obj_ref_892_store_0_req_1 : boolean;
  signal array_obj_ref_892_store_0_ack_1 : boolean;
  signal array_obj_ref_896_gather_scatter_req_0 : boolean;
  signal array_obj_ref_896_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_896_store_0_req_0 : boolean;
  signal array_obj_ref_896_store_0_ack_0 : boolean;
  signal array_obj_ref_896_store_0_req_1 : boolean;
  signal array_obj_ref_896_store_0_ack_1 : boolean;
  signal array_obj_ref_900_gather_scatter_req_0 : boolean;
  signal array_obj_ref_900_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_900_store_0_req_0 : boolean;
  signal array_obj_ref_900_store_0_ack_0 : boolean;
  signal array_obj_ref_900_store_0_req_1 : boolean;
  signal array_obj_ref_900_store_0_ack_1 : boolean;
  signal array_obj_ref_904_gather_scatter_req_0 : boolean;
  signal array_obj_ref_904_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_904_store_0_req_0 : boolean;
  signal array_obj_ref_904_store_0_ack_0 : boolean;
  signal array_obj_ref_904_store_0_req_1 : boolean;
  signal array_obj_ref_904_store_0_ack_1 : boolean;
  signal array_obj_ref_908_gather_scatter_req_0 : boolean;
  signal array_obj_ref_908_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_908_store_0_req_0 : boolean;
  signal array_obj_ref_908_store_0_ack_0 : boolean;
  signal array_obj_ref_908_store_0_req_1 : boolean;
  signal array_obj_ref_908_store_0_ack_1 : boolean;
  signal array_obj_ref_912_gather_scatter_req_0 : boolean;
  signal array_obj_ref_912_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_912_store_0_req_0 : boolean;
  signal array_obj_ref_912_store_0_ack_0 : boolean;
  signal array_obj_ref_912_store_0_req_1 : boolean;
  signal array_obj_ref_912_store_0_ack_1 : boolean;
  signal array_obj_ref_916_gather_scatter_req_0 : boolean;
  signal array_obj_ref_916_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_916_store_0_req_0 : boolean;
  signal array_obj_ref_916_store_0_ack_0 : boolean;
  signal array_obj_ref_916_store_0_req_1 : boolean;
  signal array_obj_ref_916_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 15 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr7_CP_3948: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_860_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_860_gather_scatter_ack_0;
    array_obj_ref_860_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_860_store_0_ack_0;
    array_obj_ref_860_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_860_store_0_ack_1;
    array_obj_ref_864_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_864_gather_scatter_ack_0;
    array_obj_ref_864_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_864_store_0_ack_0;
    array_obj_ref_864_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_864_store_0_ack_1;
    array_obj_ref_868_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_868_gather_scatter_ack_0;
    array_obj_ref_868_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_868_store_0_ack_0;
    array_obj_ref_868_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_868_store_0_ack_1;
    array_obj_ref_872_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_872_gather_scatter_ack_0;
    array_obj_ref_872_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_872_store_0_ack_0;
    array_obj_ref_872_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_872_store_0_ack_1;
    array_obj_ref_876_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_876_gather_scatter_ack_0;
    array_obj_ref_876_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_876_store_0_ack_0;
    array_obj_ref_876_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_876_store_0_ack_1;
    array_obj_ref_880_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_880_gather_scatter_ack_0;
    array_obj_ref_880_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_880_store_0_ack_0;
    array_obj_ref_880_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_880_store_0_ack_1;
    array_obj_ref_884_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_884_gather_scatter_ack_0;
    array_obj_ref_884_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_884_store_0_ack_0;
    array_obj_ref_884_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_884_store_0_ack_1;
    array_obj_ref_888_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_888_gather_scatter_ack_0;
    array_obj_ref_888_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_888_store_0_ack_0;
    array_obj_ref_888_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_888_store_0_ack_1;
    array_obj_ref_892_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_892_gather_scatter_ack_0;
    array_obj_ref_892_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_892_store_0_ack_0;
    array_obj_ref_892_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_892_store_0_ack_1;
    array_obj_ref_896_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_896_gather_scatter_ack_0;
    array_obj_ref_896_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_896_store_0_ack_0;
    array_obj_ref_896_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_896_store_0_ack_1;
    array_obj_ref_900_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_900_gather_scatter_ack_0;
    array_obj_ref_900_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_900_store_0_ack_0;
    array_obj_ref_900_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_900_store_0_ack_1;
    array_obj_ref_904_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_904_gather_scatter_ack_0;
    array_obj_ref_904_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_904_store_0_ack_0;
    array_obj_ref_904_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_904_store_0_ack_1;
    array_obj_ref_908_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_908_gather_scatter_ack_0;
    array_obj_ref_908_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_908_store_0_ack_0;
    array_obj_ref_908_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_908_store_0_ack_1;
    array_obj_ref_912_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_912_gather_scatter_ack_0;
    array_obj_ref_912_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_912_store_0_ack_0;
    array_obj_ref_912_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_912_store_0_ack_1;
    array_obj_ref_916_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_916_gather_scatter_ack_0;
    array_obj_ref_916_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_916_store_0_ack_0;
    array_obj_ref_916_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_916_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_860_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_860_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_864_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_864_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_868_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_868_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_872_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_872_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_876_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_876_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_880_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_880_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_884_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_884_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_888_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_888_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_892_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_892_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_896_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_896_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_900_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_900_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_904_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_904_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_908_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_908_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_912_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_912_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_916_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_916_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_861_wire_constant : std_logic_vector(7 downto 0);
    signal expr_865_wire_constant : std_logic_vector(7 downto 0);
    signal expr_869_wire_constant : std_logic_vector(7 downto 0);
    signal expr_873_wire_constant : std_logic_vector(7 downto 0);
    signal expr_877_wire_constant : std_logic_vector(7 downto 0);
    signal expr_881_wire_constant : std_logic_vector(7 downto 0);
    signal expr_885_wire_constant : std_logic_vector(7 downto 0);
    signal expr_889_wire_constant : std_logic_vector(7 downto 0);
    signal expr_893_wire_constant : std_logic_vector(7 downto 0);
    signal expr_897_wire_constant : std_logic_vector(7 downto 0);
    signal expr_901_wire_constant : std_logic_vector(7 downto 0);
    signal expr_905_wire_constant : std_logic_vector(7 downto 0);
    signal expr_909_wire_constant : std_logic_vector(7 downto 0);
    signal expr_913_wire_constant : std_logic_vector(7 downto 0);
    signal expr_917_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_860_word_address_0 <= "0000";
    array_obj_ref_864_word_address_0 <= "0001";
    array_obj_ref_868_word_address_0 <= "0010";
    array_obj_ref_872_word_address_0 <= "0011";
    array_obj_ref_876_word_address_0 <= "0100";
    array_obj_ref_880_word_address_0 <= "0101";
    array_obj_ref_884_word_address_0 <= "0110";
    array_obj_ref_888_word_address_0 <= "0111";
    array_obj_ref_892_word_address_0 <= "1000";
    array_obj_ref_896_word_address_0 <= "1001";
    array_obj_ref_900_word_address_0 <= "1010";
    array_obj_ref_904_word_address_0 <= "1011";
    array_obj_ref_908_word_address_0 <= "1100";
    array_obj_ref_912_word_address_0 <= "1101";
    array_obj_ref_916_word_address_0 <= "1110";
    expr_861_wire_constant <= "01100110";
    expr_865_wire_constant <= "01110010";
    expr_869_wire_constant <= "01100101";
    expr_873_wire_constant <= "01100101";
    expr_877_wire_constant <= "01011111";
    expr_881_wire_constant <= "01110001";
    expr_885_wire_constant <= "01110101";
    expr_889_wire_constant <= "01100101";
    expr_893_wire_constant <= "01110101";
    expr_897_wire_constant <= "01100101";
    expr_901_wire_constant <= "01011111";
    expr_905_wire_constant <= "01100111";
    expr_909_wire_constant <= "01100101";
    expr_913_wire_constant <= "01110100";
    expr_917_wire_constant <= "00000000";
    array_obj_ref_860_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_860_gather_scatter_ack_0 <= array_obj_ref_860_gather_scatter_req_0;
      aggregated_sig <= expr_861_wire_constant;
      array_obj_ref_860_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_864_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_864_gather_scatter_ack_0 <= array_obj_ref_864_gather_scatter_req_0;
      aggregated_sig <= expr_865_wire_constant;
      array_obj_ref_864_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_868_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_868_gather_scatter_ack_0 <= array_obj_ref_868_gather_scatter_req_0;
      aggregated_sig <= expr_869_wire_constant;
      array_obj_ref_868_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_872_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_872_gather_scatter_ack_0 <= array_obj_ref_872_gather_scatter_req_0;
      aggregated_sig <= expr_873_wire_constant;
      array_obj_ref_872_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_876_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_876_gather_scatter_ack_0 <= array_obj_ref_876_gather_scatter_req_0;
      aggregated_sig <= expr_877_wire_constant;
      array_obj_ref_876_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_880_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_880_gather_scatter_ack_0 <= array_obj_ref_880_gather_scatter_req_0;
      aggregated_sig <= expr_881_wire_constant;
      array_obj_ref_880_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_884_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_884_gather_scatter_ack_0 <= array_obj_ref_884_gather_scatter_req_0;
      aggregated_sig <= expr_885_wire_constant;
      array_obj_ref_884_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_888_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_888_gather_scatter_ack_0 <= array_obj_ref_888_gather_scatter_req_0;
      aggregated_sig <= expr_889_wire_constant;
      array_obj_ref_888_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_892_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_892_gather_scatter_ack_0 <= array_obj_ref_892_gather_scatter_req_0;
      aggregated_sig <= expr_893_wire_constant;
      array_obj_ref_892_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_896_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_896_gather_scatter_ack_0 <= array_obj_ref_896_gather_scatter_req_0;
      aggregated_sig <= expr_897_wire_constant;
      array_obj_ref_896_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_900_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_900_gather_scatter_ack_0 <= array_obj_ref_900_gather_scatter_req_0;
      aggregated_sig <= expr_901_wire_constant;
      array_obj_ref_900_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_904_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_904_gather_scatter_ack_0 <= array_obj_ref_904_gather_scatter_req_0;
      aggregated_sig <= expr_905_wire_constant;
      array_obj_ref_904_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_908_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_908_gather_scatter_ack_0 <= array_obj_ref_908_gather_scatter_req_0;
      aggregated_sig <= expr_909_wire_constant;
      array_obj_ref_908_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_912_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_912_gather_scatter_ack_0 <= array_obj_ref_912_gather_scatter_req_0;
      aggregated_sig <= expr_913_wire_constant;
      array_obj_ref_912_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_916_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_916_gather_scatter_ack_0 <= array_obj_ref_916_gather_scatter_req_0;
      aggregated_sig <= expr_917_wire_constant;
      array_obj_ref_916_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_860_store_0 array_obj_ref_864_store_0 array_obj_ref_868_store_0 array_obj_ref_872_store_0 array_obj_ref_876_store_0 array_obj_ref_880_store_0 array_obj_ref_884_store_0 array_obj_ref_888_store_0 array_obj_ref_892_store_0 array_obj_ref_896_store_0 array_obj_ref_900_store_0 array_obj_ref_904_store_0 array_obj_ref_908_store_0 array_obj_ref_912_store_0 array_obj_ref_916_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(59 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_860_store_0_req_0;
      reqL(13) <= array_obj_ref_864_store_0_req_0;
      reqL(12) <= array_obj_ref_868_store_0_req_0;
      reqL(11) <= array_obj_ref_872_store_0_req_0;
      reqL(10) <= array_obj_ref_876_store_0_req_0;
      reqL(9) <= array_obj_ref_880_store_0_req_0;
      reqL(8) <= array_obj_ref_884_store_0_req_0;
      reqL(7) <= array_obj_ref_888_store_0_req_0;
      reqL(6) <= array_obj_ref_892_store_0_req_0;
      reqL(5) <= array_obj_ref_896_store_0_req_0;
      reqL(4) <= array_obj_ref_900_store_0_req_0;
      reqL(3) <= array_obj_ref_904_store_0_req_0;
      reqL(2) <= array_obj_ref_908_store_0_req_0;
      reqL(1) <= array_obj_ref_912_store_0_req_0;
      reqL(0) <= array_obj_ref_916_store_0_req_0;
      array_obj_ref_860_store_0_ack_0 <= ackL(14);
      array_obj_ref_864_store_0_ack_0 <= ackL(13);
      array_obj_ref_868_store_0_ack_0 <= ackL(12);
      array_obj_ref_872_store_0_ack_0 <= ackL(11);
      array_obj_ref_876_store_0_ack_0 <= ackL(10);
      array_obj_ref_880_store_0_ack_0 <= ackL(9);
      array_obj_ref_884_store_0_ack_0 <= ackL(8);
      array_obj_ref_888_store_0_ack_0 <= ackL(7);
      array_obj_ref_892_store_0_ack_0 <= ackL(6);
      array_obj_ref_896_store_0_ack_0 <= ackL(5);
      array_obj_ref_900_store_0_ack_0 <= ackL(4);
      array_obj_ref_904_store_0_ack_0 <= ackL(3);
      array_obj_ref_908_store_0_ack_0 <= ackL(2);
      array_obj_ref_912_store_0_ack_0 <= ackL(1);
      array_obj_ref_916_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_860_store_0_req_1;
      reqR(13) <= array_obj_ref_864_store_0_req_1;
      reqR(12) <= array_obj_ref_868_store_0_req_1;
      reqR(11) <= array_obj_ref_872_store_0_req_1;
      reqR(10) <= array_obj_ref_876_store_0_req_1;
      reqR(9) <= array_obj_ref_880_store_0_req_1;
      reqR(8) <= array_obj_ref_884_store_0_req_1;
      reqR(7) <= array_obj_ref_888_store_0_req_1;
      reqR(6) <= array_obj_ref_892_store_0_req_1;
      reqR(5) <= array_obj_ref_896_store_0_req_1;
      reqR(4) <= array_obj_ref_900_store_0_req_1;
      reqR(3) <= array_obj_ref_904_store_0_req_1;
      reqR(2) <= array_obj_ref_908_store_0_req_1;
      reqR(1) <= array_obj_ref_912_store_0_req_1;
      reqR(0) <= array_obj_ref_916_store_0_req_1;
      array_obj_ref_860_store_0_ack_1 <= ackR(14);
      array_obj_ref_864_store_0_ack_1 <= ackR(13);
      array_obj_ref_868_store_0_ack_1 <= ackR(12);
      array_obj_ref_872_store_0_ack_1 <= ackR(11);
      array_obj_ref_876_store_0_ack_1 <= ackR(10);
      array_obj_ref_880_store_0_ack_1 <= ackR(9);
      array_obj_ref_884_store_0_ack_1 <= ackR(8);
      array_obj_ref_888_store_0_ack_1 <= ackR(7);
      array_obj_ref_892_store_0_ack_1 <= ackR(6);
      array_obj_ref_896_store_0_ack_1 <= ackR(5);
      array_obj_ref_900_store_0_ack_1 <= ackR(4);
      array_obj_ref_904_store_0_ack_1 <= ackR(3);
      array_obj_ref_908_store_0_ack_1 <= ackR(2);
      array_obj_ref_912_store_0_ack_1 <= ackR(1);
      array_obj_ref_916_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_860_word_address_0 & array_obj_ref_864_word_address_0 & array_obj_ref_868_word_address_0 & array_obj_ref_872_word_address_0 & array_obj_ref_876_word_address_0 & array_obj_ref_880_word_address_0 & array_obj_ref_884_word_address_0 & array_obj_ref_888_word_address_0 & array_obj_ref_892_word_address_0 & array_obj_ref_896_word_address_0 & array_obj_ref_900_word_address_0 & array_obj_ref_904_word_address_0 & array_obj_ref_908_word_address_0 & array_obj_ref_912_word_address_0 & array_obj_ref_916_word_address_0;
      data_in <= array_obj_ref_860_data_0 & array_obj_ref_864_data_0 & array_obj_ref_868_data_0 & array_obj_ref_872_data_0 & array_obj_ref_876_data_0 & array_obj_ref_880_data_0 & array_obj_ref_884_data_0 & array_obj_ref_888_data_0 & array_obj_ref_892_data_0 & array_obj_ref_896_data_0 & array_obj_ref_900_data_0 & array_obj_ref_904_data_0 & array_obj_ref_908_data_0 & array_obj_ref_912_data_0 & array_obj_ref_916_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 15,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_17_sr_req(0),
          mack => memory_space_17_sr_ack(0),
          maddr => memory_space_17_sr_addr(3 downto 0),
          mdata => memory_space_17_sr_data(7 downto 0),
          mtag => memory_space_17_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_17_sc_req(0),
          mack => memory_space_17_sc_ack(0),
          mtag => memory_space_17_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr8 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_18_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_18_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_18_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_18_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_18_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_18_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_18_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_18_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr8;
architecture Default of default_initializer_xx_xstr8 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr8_CP_4266_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_934_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_930_store_0_ack_0 : boolean;
  signal array_obj_ref_962_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_958_store_0_ack_0 : boolean;
  signal array_obj_ref_922_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_922_store_0_ack_1 : boolean;
  signal array_obj_ref_978_store_0_ack_1 : boolean;
  signal array_obj_ref_974_gather_scatter_req_0 : boolean;
  signal array_obj_ref_938_store_0_ack_1 : boolean;
  signal array_obj_ref_934_gather_scatter_req_0 : boolean;
  signal array_obj_ref_950_gather_scatter_req_0 : boolean;
  signal array_obj_ref_978_store_0_req_1 : boolean;
  signal array_obj_ref_958_store_0_req_1 : boolean;
  signal array_obj_ref_978_store_0_req_0 : boolean;
  signal array_obj_ref_962_gather_scatter_req_0 : boolean;
  signal array_obj_ref_954_gather_scatter_req_0 : boolean;
  signal array_obj_ref_958_store_0_ack_1 : boolean;
  signal array_obj_ref_922_gather_scatter_req_0 : boolean;
  signal array_obj_ref_954_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_954_store_0_req_0 : boolean;
  signal array_obj_ref_922_store_0_req_0 : boolean;
  signal array_obj_ref_922_store_0_ack_0 : boolean;
  signal array_obj_ref_922_store_0_req_1 : boolean;
  signal array_obj_ref_942_gather_scatter_req_0 : boolean;
  signal array_obj_ref_942_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_978_store_0_ack_0 : boolean;
  signal array_obj_ref_974_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_934_store_0_req_0 : boolean;
  signal array_obj_ref_954_store_0_req_1 : boolean;
  signal array_obj_ref_962_store_0_ack_0 : boolean;
  signal array_obj_ref_974_store_0_req_0 : boolean;
  signal array_obj_ref_962_store_0_req_1 : boolean;
  signal array_obj_ref_926_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_974_store_0_ack_0 : boolean;
  signal array_obj_ref_954_store_0_ack_1 : boolean;
  signal array_obj_ref_962_store_0_req_0 : boolean;
  signal array_obj_ref_954_store_0_ack_0 : boolean;
  signal array_obj_ref_926_gather_scatter_req_0 : boolean;
  signal array_obj_ref_934_store_0_ack_0 : boolean;
  signal array_obj_ref_934_store_0_req_1 : boolean;
  signal array_obj_ref_934_store_0_ack_1 : boolean;
  signal array_obj_ref_974_store_0_req_1 : boolean;
  signal array_obj_ref_970_store_0_req_1 : boolean;
  signal array_obj_ref_958_store_0_req_0 : boolean;
  signal array_obj_ref_950_store_0_ack_1 : boolean;
  signal array_obj_ref_950_store_0_req_1 : boolean;
  signal array_obj_ref_938_store_0_req_1 : boolean;
  signal array_obj_ref_938_store_0_ack_0 : boolean;
  signal array_obj_ref_950_store_0_ack_0 : boolean;
  signal array_obj_ref_950_store_0_req_0 : boolean;
  signal array_obj_ref_950_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_930_store_0_req_1 : boolean;
  signal array_obj_ref_930_store_0_ack_1 : boolean;
  signal array_obj_ref_970_store_0_ack_1 : boolean;
  signal array_obj_ref_974_store_0_ack_1 : boolean;
  signal array_obj_ref_962_store_0_ack_1 : boolean;
  signal array_obj_ref_958_gather_scatter_req_0 : boolean;
  signal array_obj_ref_926_store_0_req_0 : boolean;
  signal array_obj_ref_926_store_0_ack_0 : boolean;
  signal array_obj_ref_958_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_926_store_0_req_1 : boolean;
  signal array_obj_ref_926_store_0_ack_1 : boolean;
  signal array_obj_ref_978_gather_scatter_req_0 : boolean;
  signal array_obj_ref_978_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_938_gather_scatter_req_0 : boolean;
  signal array_obj_ref_938_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_938_store_0_req_0 : boolean;
  signal array_obj_ref_970_store_0_ack_0 : boolean;
  signal array_obj_ref_970_store_0_req_0 : boolean;
  signal array_obj_ref_946_store_0_ack_1 : boolean;
  signal array_obj_ref_946_store_0_req_1 : boolean;
  signal array_obj_ref_970_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_970_gather_scatter_req_0 : boolean;
  signal array_obj_ref_946_store_0_ack_0 : boolean;
  signal array_obj_ref_946_store_0_req_0 : boolean;
  signal array_obj_ref_946_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_946_gather_scatter_req_0 : boolean;
  signal array_obj_ref_966_store_0_ack_1 : boolean;
  signal array_obj_ref_966_store_0_req_1 : boolean;
  signal array_obj_ref_966_store_0_ack_0 : boolean;
  signal array_obj_ref_966_store_0_req_0 : boolean;
  signal array_obj_ref_942_store_0_ack_1 : boolean;
  signal array_obj_ref_966_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_942_store_0_req_1 : boolean;
  signal array_obj_ref_966_gather_scatter_req_0 : boolean;
  signal array_obj_ref_942_store_0_ack_0 : boolean;
  signal array_obj_ref_942_store_0_req_0 : boolean;
  signal array_obj_ref_930_store_0_req_0 : boolean;
  signal array_obj_ref_930_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_930_gather_scatter_req_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 15 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr8_CP_4266: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_922_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_922_gather_scatter_ack_0;
    array_obj_ref_922_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_922_store_0_ack_0;
    array_obj_ref_922_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_922_store_0_ack_1;
    array_obj_ref_926_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_926_gather_scatter_ack_0;
    array_obj_ref_926_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_926_store_0_ack_0;
    array_obj_ref_926_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_926_store_0_ack_1;
    array_obj_ref_930_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_930_gather_scatter_ack_0;
    array_obj_ref_930_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_930_store_0_ack_0;
    array_obj_ref_930_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_930_store_0_ack_1;
    array_obj_ref_934_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_934_gather_scatter_ack_0;
    array_obj_ref_934_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_934_store_0_ack_0;
    array_obj_ref_934_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_934_store_0_ack_1;
    array_obj_ref_938_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_938_gather_scatter_ack_0;
    array_obj_ref_938_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_938_store_0_ack_0;
    array_obj_ref_938_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_938_store_0_ack_1;
    array_obj_ref_942_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_942_gather_scatter_ack_0;
    array_obj_ref_942_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_942_store_0_ack_0;
    array_obj_ref_942_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_942_store_0_ack_1;
    array_obj_ref_946_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_946_gather_scatter_ack_0;
    array_obj_ref_946_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_946_store_0_ack_0;
    array_obj_ref_946_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_946_store_0_ack_1;
    array_obj_ref_950_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_950_gather_scatter_ack_0;
    array_obj_ref_950_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_950_store_0_ack_0;
    array_obj_ref_950_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_950_store_0_ack_1;
    array_obj_ref_954_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_954_gather_scatter_ack_0;
    array_obj_ref_954_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_954_store_0_ack_0;
    array_obj_ref_954_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_954_store_0_ack_1;
    array_obj_ref_958_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_958_gather_scatter_ack_0;
    array_obj_ref_958_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_958_store_0_ack_0;
    array_obj_ref_958_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_958_store_0_ack_1;
    array_obj_ref_962_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_962_gather_scatter_ack_0;
    array_obj_ref_962_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_962_store_0_ack_0;
    array_obj_ref_962_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_962_store_0_ack_1;
    array_obj_ref_966_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_966_gather_scatter_ack_0;
    array_obj_ref_966_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_966_store_0_ack_0;
    array_obj_ref_966_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_966_store_0_ack_1;
    array_obj_ref_970_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_970_gather_scatter_ack_0;
    array_obj_ref_970_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_970_store_0_ack_0;
    array_obj_ref_970_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_970_store_0_ack_1;
    array_obj_ref_974_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_974_gather_scatter_ack_0;
    array_obj_ref_974_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_974_store_0_ack_0;
    array_obj_ref_974_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_974_store_0_ack_1;
    array_obj_ref_978_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_978_gather_scatter_ack_0;
    array_obj_ref_978_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_978_store_0_ack_0;
    array_obj_ref_978_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_978_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_922_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_922_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_926_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_926_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_930_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_930_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_934_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_934_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_938_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_938_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_942_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_942_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_946_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_946_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_950_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_950_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_954_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_954_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_958_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_958_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_962_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_962_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_966_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_966_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_970_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_970_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_974_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_974_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_978_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_978_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_923_wire_constant : std_logic_vector(7 downto 0);
    signal expr_927_wire_constant : std_logic_vector(7 downto 0);
    signal expr_931_wire_constant : std_logic_vector(7 downto 0);
    signal expr_935_wire_constant : std_logic_vector(7 downto 0);
    signal expr_939_wire_constant : std_logic_vector(7 downto 0);
    signal expr_943_wire_constant : std_logic_vector(7 downto 0);
    signal expr_947_wire_constant : std_logic_vector(7 downto 0);
    signal expr_951_wire_constant : std_logic_vector(7 downto 0);
    signal expr_955_wire_constant : std_logic_vector(7 downto 0);
    signal expr_959_wire_constant : std_logic_vector(7 downto 0);
    signal expr_963_wire_constant : std_logic_vector(7 downto 0);
    signal expr_967_wire_constant : std_logic_vector(7 downto 0);
    signal expr_971_wire_constant : std_logic_vector(7 downto 0);
    signal expr_975_wire_constant : std_logic_vector(7 downto 0);
    signal expr_979_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_922_word_address_0 <= "0000";
    array_obj_ref_926_word_address_0 <= "0001";
    array_obj_ref_930_word_address_0 <= "0010";
    array_obj_ref_934_word_address_0 <= "0011";
    array_obj_ref_938_word_address_0 <= "0100";
    array_obj_ref_942_word_address_0 <= "0101";
    array_obj_ref_946_word_address_0 <= "0110";
    array_obj_ref_950_word_address_0 <= "0111";
    array_obj_ref_954_word_address_0 <= "1000";
    array_obj_ref_958_word_address_0 <= "1001";
    array_obj_ref_962_word_address_0 <= "1010";
    array_obj_ref_966_word_address_0 <= "1011";
    array_obj_ref_970_word_address_0 <= "1100";
    array_obj_ref_974_word_address_0 <= "1101";
    array_obj_ref_978_word_address_0 <= "1110";
    expr_923_wire_constant <= "01100110";
    expr_927_wire_constant <= "01110010";
    expr_931_wire_constant <= "01100101";
    expr_935_wire_constant <= "01100101";
    expr_939_wire_constant <= "01011111";
    expr_943_wire_constant <= "01110001";
    expr_947_wire_constant <= "01110101";
    expr_951_wire_constant <= "01100101";
    expr_955_wire_constant <= "01110101";
    expr_959_wire_constant <= "01100101";
    expr_963_wire_constant <= "01011111";
    expr_967_wire_constant <= "01110000";
    expr_971_wire_constant <= "01110101";
    expr_975_wire_constant <= "01110100";
    expr_979_wire_constant <= "00000000";
    array_obj_ref_922_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_922_gather_scatter_ack_0 <= array_obj_ref_922_gather_scatter_req_0;
      aggregated_sig <= expr_923_wire_constant;
      array_obj_ref_922_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_926_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_926_gather_scatter_ack_0 <= array_obj_ref_926_gather_scatter_req_0;
      aggregated_sig <= expr_927_wire_constant;
      array_obj_ref_926_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_930_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_930_gather_scatter_ack_0 <= array_obj_ref_930_gather_scatter_req_0;
      aggregated_sig <= expr_931_wire_constant;
      array_obj_ref_930_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_934_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_934_gather_scatter_ack_0 <= array_obj_ref_934_gather_scatter_req_0;
      aggregated_sig <= expr_935_wire_constant;
      array_obj_ref_934_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_938_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_938_gather_scatter_ack_0 <= array_obj_ref_938_gather_scatter_req_0;
      aggregated_sig <= expr_939_wire_constant;
      array_obj_ref_938_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_942_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_942_gather_scatter_ack_0 <= array_obj_ref_942_gather_scatter_req_0;
      aggregated_sig <= expr_943_wire_constant;
      array_obj_ref_942_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_946_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_946_gather_scatter_ack_0 <= array_obj_ref_946_gather_scatter_req_0;
      aggregated_sig <= expr_947_wire_constant;
      array_obj_ref_946_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_950_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_950_gather_scatter_ack_0 <= array_obj_ref_950_gather_scatter_req_0;
      aggregated_sig <= expr_951_wire_constant;
      array_obj_ref_950_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_954_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_954_gather_scatter_ack_0 <= array_obj_ref_954_gather_scatter_req_0;
      aggregated_sig <= expr_955_wire_constant;
      array_obj_ref_954_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_958_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_958_gather_scatter_ack_0 <= array_obj_ref_958_gather_scatter_req_0;
      aggregated_sig <= expr_959_wire_constant;
      array_obj_ref_958_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_962_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_962_gather_scatter_ack_0 <= array_obj_ref_962_gather_scatter_req_0;
      aggregated_sig <= expr_963_wire_constant;
      array_obj_ref_962_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_966_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_966_gather_scatter_ack_0 <= array_obj_ref_966_gather_scatter_req_0;
      aggregated_sig <= expr_967_wire_constant;
      array_obj_ref_966_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_970_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_970_gather_scatter_ack_0 <= array_obj_ref_970_gather_scatter_req_0;
      aggregated_sig <= expr_971_wire_constant;
      array_obj_ref_970_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_974_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_974_gather_scatter_ack_0 <= array_obj_ref_974_gather_scatter_req_0;
      aggregated_sig <= expr_975_wire_constant;
      array_obj_ref_974_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_978_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_978_gather_scatter_ack_0 <= array_obj_ref_978_gather_scatter_req_0;
      aggregated_sig <= expr_979_wire_constant;
      array_obj_ref_978_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_970_store_0 array_obj_ref_950_store_0 array_obj_ref_978_store_0 array_obj_ref_954_store_0 array_obj_ref_958_store_0 array_obj_ref_962_store_0 array_obj_ref_966_store_0 array_obj_ref_974_store_0 array_obj_ref_946_store_0 array_obj_ref_942_store_0 array_obj_ref_938_store_0 array_obj_ref_934_store_0 array_obj_ref_930_store_0 array_obj_ref_926_store_0 array_obj_ref_922_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(59 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_970_store_0_req_0;
      reqL(13) <= array_obj_ref_950_store_0_req_0;
      reqL(12) <= array_obj_ref_978_store_0_req_0;
      reqL(11) <= array_obj_ref_954_store_0_req_0;
      reqL(10) <= array_obj_ref_958_store_0_req_0;
      reqL(9) <= array_obj_ref_962_store_0_req_0;
      reqL(8) <= array_obj_ref_966_store_0_req_0;
      reqL(7) <= array_obj_ref_974_store_0_req_0;
      reqL(6) <= array_obj_ref_946_store_0_req_0;
      reqL(5) <= array_obj_ref_942_store_0_req_0;
      reqL(4) <= array_obj_ref_938_store_0_req_0;
      reqL(3) <= array_obj_ref_934_store_0_req_0;
      reqL(2) <= array_obj_ref_930_store_0_req_0;
      reqL(1) <= array_obj_ref_926_store_0_req_0;
      reqL(0) <= array_obj_ref_922_store_0_req_0;
      array_obj_ref_970_store_0_ack_0 <= ackL(14);
      array_obj_ref_950_store_0_ack_0 <= ackL(13);
      array_obj_ref_978_store_0_ack_0 <= ackL(12);
      array_obj_ref_954_store_0_ack_0 <= ackL(11);
      array_obj_ref_958_store_0_ack_0 <= ackL(10);
      array_obj_ref_962_store_0_ack_0 <= ackL(9);
      array_obj_ref_966_store_0_ack_0 <= ackL(8);
      array_obj_ref_974_store_0_ack_0 <= ackL(7);
      array_obj_ref_946_store_0_ack_0 <= ackL(6);
      array_obj_ref_942_store_0_ack_0 <= ackL(5);
      array_obj_ref_938_store_0_ack_0 <= ackL(4);
      array_obj_ref_934_store_0_ack_0 <= ackL(3);
      array_obj_ref_930_store_0_ack_0 <= ackL(2);
      array_obj_ref_926_store_0_ack_0 <= ackL(1);
      array_obj_ref_922_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_970_store_0_req_1;
      reqR(13) <= array_obj_ref_950_store_0_req_1;
      reqR(12) <= array_obj_ref_978_store_0_req_1;
      reqR(11) <= array_obj_ref_954_store_0_req_1;
      reqR(10) <= array_obj_ref_958_store_0_req_1;
      reqR(9) <= array_obj_ref_962_store_0_req_1;
      reqR(8) <= array_obj_ref_966_store_0_req_1;
      reqR(7) <= array_obj_ref_974_store_0_req_1;
      reqR(6) <= array_obj_ref_946_store_0_req_1;
      reqR(5) <= array_obj_ref_942_store_0_req_1;
      reqR(4) <= array_obj_ref_938_store_0_req_1;
      reqR(3) <= array_obj_ref_934_store_0_req_1;
      reqR(2) <= array_obj_ref_930_store_0_req_1;
      reqR(1) <= array_obj_ref_926_store_0_req_1;
      reqR(0) <= array_obj_ref_922_store_0_req_1;
      array_obj_ref_970_store_0_ack_1 <= ackR(14);
      array_obj_ref_950_store_0_ack_1 <= ackR(13);
      array_obj_ref_978_store_0_ack_1 <= ackR(12);
      array_obj_ref_954_store_0_ack_1 <= ackR(11);
      array_obj_ref_958_store_0_ack_1 <= ackR(10);
      array_obj_ref_962_store_0_ack_1 <= ackR(9);
      array_obj_ref_966_store_0_ack_1 <= ackR(8);
      array_obj_ref_974_store_0_ack_1 <= ackR(7);
      array_obj_ref_946_store_0_ack_1 <= ackR(6);
      array_obj_ref_942_store_0_ack_1 <= ackR(5);
      array_obj_ref_938_store_0_ack_1 <= ackR(4);
      array_obj_ref_934_store_0_ack_1 <= ackR(3);
      array_obj_ref_930_store_0_ack_1 <= ackR(2);
      array_obj_ref_926_store_0_ack_1 <= ackR(1);
      array_obj_ref_922_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_970_word_address_0 & array_obj_ref_950_word_address_0 & array_obj_ref_978_word_address_0 & array_obj_ref_954_word_address_0 & array_obj_ref_958_word_address_0 & array_obj_ref_962_word_address_0 & array_obj_ref_966_word_address_0 & array_obj_ref_974_word_address_0 & array_obj_ref_946_word_address_0 & array_obj_ref_942_word_address_0 & array_obj_ref_938_word_address_0 & array_obj_ref_934_word_address_0 & array_obj_ref_930_word_address_0 & array_obj_ref_926_word_address_0 & array_obj_ref_922_word_address_0;
      data_in <= array_obj_ref_970_data_0 & array_obj_ref_950_data_0 & array_obj_ref_978_data_0 & array_obj_ref_954_data_0 & array_obj_ref_958_data_0 & array_obj_ref_962_data_0 & array_obj_ref_966_data_0 & array_obj_ref_974_data_0 & array_obj_ref_946_data_0 & array_obj_ref_942_data_0 & array_obj_ref_938_data_0 & array_obj_ref_934_data_0 & array_obj_ref_930_data_0 & array_obj_ref_926_data_0 & array_obj_ref_922_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 15,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_18_sr_req(0),
          mack => memory_space_18_sr_ack(0),
          maddr => memory_space_18_sr_addr(3 downto 0),
          mdata => memory_space_18_sr_data(7 downto 0),
          mtag => memory_space_18_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_18_sc_req(0),
          mack => memory_space_18_sc_ack(0),
          mtag => memory_space_18_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr9 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_19_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_19_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_19_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_19_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_19_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_19_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_19_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_19_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr9;
architecture Default of default_initializer_xx_xstr9 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr9_CP_4584_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_984_gather_scatter_req_0 : boolean;
  signal array_obj_ref_984_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_984_store_0_req_0 : boolean;
  signal array_obj_ref_984_store_0_ack_0 : boolean;
  signal array_obj_ref_984_store_0_req_1 : boolean;
  signal array_obj_ref_984_store_0_ack_1 : boolean;
  signal array_obj_ref_988_gather_scatter_req_0 : boolean;
  signal array_obj_ref_988_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_988_store_0_req_0 : boolean;
  signal array_obj_ref_988_store_0_ack_0 : boolean;
  signal array_obj_ref_988_store_0_req_1 : boolean;
  signal array_obj_ref_988_store_0_ack_1 : boolean;
  signal array_obj_ref_992_gather_scatter_req_0 : boolean;
  signal array_obj_ref_992_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_992_store_0_req_0 : boolean;
  signal array_obj_ref_992_store_0_ack_0 : boolean;
  signal array_obj_ref_992_store_0_req_1 : boolean;
  signal array_obj_ref_992_store_0_ack_1 : boolean;
  signal array_obj_ref_996_gather_scatter_req_0 : boolean;
  signal array_obj_ref_996_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_996_store_0_req_0 : boolean;
  signal array_obj_ref_996_store_0_ack_0 : boolean;
  signal array_obj_ref_996_store_0_req_1 : boolean;
  signal array_obj_ref_996_store_0_ack_1 : boolean;
  signal array_obj_ref_1000_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1000_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1000_store_0_req_0 : boolean;
  signal array_obj_ref_1000_store_0_ack_0 : boolean;
  signal array_obj_ref_1000_store_0_req_1 : boolean;
  signal array_obj_ref_1000_store_0_ack_1 : boolean;
  signal array_obj_ref_1004_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1004_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1004_store_0_req_0 : boolean;
  signal array_obj_ref_1004_store_0_ack_0 : boolean;
  signal array_obj_ref_1004_store_0_req_1 : boolean;
  signal array_obj_ref_1004_store_0_ack_1 : boolean;
  signal array_obj_ref_1008_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1008_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1008_store_0_req_0 : boolean;
  signal array_obj_ref_1008_store_0_ack_0 : boolean;
  signal array_obj_ref_1008_store_0_req_1 : boolean;
  signal array_obj_ref_1008_store_0_ack_1 : boolean;
  signal array_obj_ref_1012_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1012_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1012_store_0_req_0 : boolean;
  signal array_obj_ref_1012_store_0_ack_0 : boolean;
  signal array_obj_ref_1012_store_0_req_1 : boolean;
  signal array_obj_ref_1012_store_0_ack_1 : boolean;
  signal array_obj_ref_1016_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1016_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1016_store_0_req_0 : boolean;
  signal array_obj_ref_1016_store_0_ack_0 : boolean;
  signal array_obj_ref_1016_store_0_req_1 : boolean;
  signal array_obj_ref_1016_store_0_ack_1 : boolean;
  signal array_obj_ref_1020_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1020_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1020_store_0_req_0 : boolean;
  signal array_obj_ref_1020_store_0_ack_0 : boolean;
  signal array_obj_ref_1020_store_0_req_1 : boolean;
  signal array_obj_ref_1020_store_0_ack_1 : boolean;
  signal array_obj_ref_1024_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1024_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1024_store_0_req_0 : boolean;
  signal array_obj_ref_1024_store_0_ack_0 : boolean;
  signal array_obj_ref_1024_store_0_req_1 : boolean;
  signal array_obj_ref_1024_store_0_ack_1 : boolean;
  signal array_obj_ref_1028_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1028_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1028_store_0_req_0 : boolean;
  signal array_obj_ref_1028_store_0_ack_0 : boolean;
  signal array_obj_ref_1028_store_0_req_1 : boolean;
  signal array_obj_ref_1028_store_0_ack_1 : boolean;
  signal array_obj_ref_1032_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1032_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1032_store_0_req_0 : boolean;
  signal array_obj_ref_1032_store_0_ack_0 : boolean;
  signal array_obj_ref_1032_store_0_req_1 : boolean;
  signal array_obj_ref_1032_store_0_ack_1 : boolean;
  signal array_obj_ref_1036_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1036_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1036_store_0_req_0 : boolean;
  signal array_obj_ref_1036_store_0_ack_0 : boolean;
  signal array_obj_ref_1036_store_0_req_1 : boolean;
  signal array_obj_ref_1036_store_0_ack_1 : boolean;
  signal array_obj_ref_1040_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1040_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1040_store_0_req_0 : boolean;
  signal array_obj_ref_1040_store_0_ack_0 : boolean;
  signal array_obj_ref_1040_store_0_req_1 : boolean;
  signal array_obj_ref_1040_store_0_ack_1 : boolean;
  signal array_obj_ref_1044_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1044_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1044_store_0_req_0 : boolean;
  signal array_obj_ref_1044_store_0_ack_0 : boolean;
  signal array_obj_ref_1044_store_0_req_1 : boolean;
  signal array_obj_ref_1044_store_0_ack_1 : boolean;
  signal array_obj_ref_1048_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1048_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1048_store_0_req_0 : boolean;
  signal array_obj_ref_1048_store_0_ack_0 : boolean;
  signal array_obj_ref_1048_store_0_req_1 : boolean;
  signal array_obj_ref_1048_store_0_ack_1 : boolean;
  signal array_obj_ref_1052_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1052_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1052_store_0_req_0 : boolean;
  signal array_obj_ref_1052_store_0_ack_0 : boolean;
  signal array_obj_ref_1052_store_0_req_1 : boolean;
  signal array_obj_ref_1052_store_0_ack_1 : boolean;
  signal array_obj_ref_1056_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1056_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1056_store_0_req_0 : boolean;
  signal array_obj_ref_1056_store_0_ack_0 : boolean;
  signal array_obj_ref_1056_store_0_req_1 : boolean;
  signal array_obj_ref_1056_store_0_ack_1 : boolean;
  signal array_obj_ref_1060_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1060_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1060_store_0_req_0 : boolean;
  signal array_obj_ref_1060_store_0_ack_0 : boolean;
  signal array_obj_ref_1060_store_0_req_1 : boolean;
  signal array_obj_ref_1060_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 20 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr9_CP_4584: Block -- control-path 
    signal cp_elements: BooleanArray(60 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(60);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(60), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_984_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_984_gather_scatter_ack_0;
    array_obj_ref_984_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_984_store_0_ack_0;
    array_obj_ref_984_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_984_store_0_ack_1;
    array_obj_ref_988_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_988_gather_scatter_ack_0;
    array_obj_ref_988_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_988_store_0_ack_0;
    array_obj_ref_988_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_988_store_0_ack_1;
    array_obj_ref_992_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_992_gather_scatter_ack_0;
    array_obj_ref_992_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_992_store_0_ack_0;
    array_obj_ref_992_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_992_store_0_ack_1;
    array_obj_ref_996_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_996_gather_scatter_ack_0;
    array_obj_ref_996_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_996_store_0_ack_0;
    array_obj_ref_996_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_996_store_0_ack_1;
    array_obj_ref_1000_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_1000_gather_scatter_ack_0;
    array_obj_ref_1000_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_1000_store_0_ack_0;
    array_obj_ref_1000_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_1000_store_0_ack_1;
    array_obj_ref_1004_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_1004_gather_scatter_ack_0;
    array_obj_ref_1004_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_1004_store_0_ack_0;
    array_obj_ref_1004_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_1004_store_0_ack_1;
    array_obj_ref_1008_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_1008_gather_scatter_ack_0;
    array_obj_ref_1008_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_1008_store_0_ack_0;
    array_obj_ref_1008_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_1008_store_0_ack_1;
    array_obj_ref_1012_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_1012_gather_scatter_ack_0;
    array_obj_ref_1012_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_1012_store_0_ack_0;
    array_obj_ref_1012_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_1012_store_0_ack_1;
    array_obj_ref_1016_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_1016_gather_scatter_ack_0;
    array_obj_ref_1016_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_1016_store_0_ack_0;
    array_obj_ref_1016_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_1016_store_0_ack_1;
    array_obj_ref_1020_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_1020_gather_scatter_ack_0;
    array_obj_ref_1020_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_1020_store_0_ack_0;
    array_obj_ref_1020_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_1020_store_0_ack_1;
    array_obj_ref_1024_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_1024_gather_scatter_ack_0;
    array_obj_ref_1024_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_1024_store_0_ack_0;
    array_obj_ref_1024_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_1024_store_0_ack_1;
    array_obj_ref_1028_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_1028_gather_scatter_ack_0;
    array_obj_ref_1028_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_1028_store_0_ack_0;
    array_obj_ref_1028_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_1028_store_0_ack_1;
    array_obj_ref_1032_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_1032_gather_scatter_ack_0;
    array_obj_ref_1032_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_1032_store_0_ack_0;
    array_obj_ref_1032_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_1032_store_0_ack_1;
    array_obj_ref_1036_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_1036_gather_scatter_ack_0;
    array_obj_ref_1036_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_1036_store_0_ack_0;
    array_obj_ref_1036_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_1036_store_0_ack_1;
    array_obj_ref_1040_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_1040_gather_scatter_ack_0;
    array_obj_ref_1040_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_1040_store_0_ack_0;
    array_obj_ref_1040_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_1040_store_0_ack_1;
    array_obj_ref_1044_gather_scatter_req_0 <= cp_elements(45);
    cp_elements(46) <= array_obj_ref_1044_gather_scatter_ack_0;
    array_obj_ref_1044_store_0_req_0 <= cp_elements(46);
    cp_elements(47) <= array_obj_ref_1044_store_0_ack_0;
    array_obj_ref_1044_store_0_req_1 <= cp_elements(47);
    cp_elements(48) <= array_obj_ref_1044_store_0_ack_1;
    array_obj_ref_1048_gather_scatter_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_1048_gather_scatter_ack_0;
    array_obj_ref_1048_store_0_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_1048_store_0_ack_0;
    array_obj_ref_1048_store_0_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_1048_store_0_ack_1;
    array_obj_ref_1052_gather_scatter_req_0 <= cp_elements(51);
    cp_elements(52) <= array_obj_ref_1052_gather_scatter_ack_0;
    array_obj_ref_1052_store_0_req_0 <= cp_elements(52);
    cp_elements(53) <= array_obj_ref_1052_store_0_ack_0;
    array_obj_ref_1052_store_0_req_1 <= cp_elements(53);
    cp_elements(54) <= array_obj_ref_1052_store_0_ack_1;
    array_obj_ref_1056_gather_scatter_req_0 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_1056_gather_scatter_ack_0;
    array_obj_ref_1056_store_0_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_1056_store_0_ack_0;
    array_obj_ref_1056_store_0_req_1 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_1056_store_0_ack_1;
    array_obj_ref_1060_gather_scatter_req_0 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_1060_gather_scatter_ack_0;
    array_obj_ref_1060_store_0_req_0 <= cp_elements(58);
    cp_elements(59) <= array_obj_ref_1060_store_0_ack_0;
    array_obj_ref_1060_store_0_req_1 <= cp_elements(59);
    cp_elements(60) <= array_obj_ref_1060_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1000_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1000_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1004_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1004_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1008_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1008_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1012_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1012_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1016_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1016_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1020_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1020_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1024_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1024_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1028_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1028_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1032_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1032_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1036_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1036_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1040_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1040_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1044_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1044_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1048_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1048_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1052_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1052_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1056_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1056_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1060_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_1060_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_984_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_984_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_988_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_988_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_992_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_992_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_996_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_996_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_1001_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1005_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1009_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1013_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1017_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1021_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1025_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1029_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1033_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1037_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1041_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1045_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1049_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1053_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1057_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1061_wire_constant : std_logic_vector(7 downto 0);
    signal expr_985_wire_constant : std_logic_vector(7 downto 0);
    signal expr_989_wire_constant : std_logic_vector(7 downto 0);
    signal expr_993_wire_constant : std_logic_vector(7 downto 0);
    signal expr_997_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1000_word_address_0 <= "00100";
    array_obj_ref_1004_word_address_0 <= "00101";
    array_obj_ref_1008_word_address_0 <= "00110";
    array_obj_ref_1012_word_address_0 <= "00111";
    array_obj_ref_1016_word_address_0 <= "01000";
    array_obj_ref_1020_word_address_0 <= "01001";
    array_obj_ref_1024_word_address_0 <= "01010";
    array_obj_ref_1028_word_address_0 <= "01011";
    array_obj_ref_1032_word_address_0 <= "01100";
    array_obj_ref_1036_word_address_0 <= "01101";
    array_obj_ref_1040_word_address_0 <= "01110";
    array_obj_ref_1044_word_address_0 <= "01111";
    array_obj_ref_1048_word_address_0 <= "10000";
    array_obj_ref_1052_word_address_0 <= "10001";
    array_obj_ref_1056_word_address_0 <= "10010";
    array_obj_ref_1060_word_address_0 <= "10011";
    array_obj_ref_984_word_address_0 <= "00000";
    array_obj_ref_988_word_address_0 <= "00001";
    array_obj_ref_992_word_address_0 <= "00010";
    array_obj_ref_996_word_address_0 <= "00011";
    expr_1001_wire_constant <= "01110100";
    expr_1005_wire_constant <= "01011111";
    expr_1009_wire_constant <= "01110111";
    expr_1013_wire_constant <= "01110010";
    expr_1017_wire_constant <= "01100001";
    expr_1021_wire_constant <= "01110000";
    expr_1025_wire_constant <= "01110000";
    expr_1029_wire_constant <= "01100101";
    expr_1033_wire_constant <= "01110010";
    expr_1037_wire_constant <= "01011111";
    expr_1041_wire_constant <= "01101001";
    expr_1045_wire_constant <= "01101110";
    expr_1049_wire_constant <= "01110000";
    expr_1053_wire_constant <= "01110101";
    expr_1057_wire_constant <= "01110100";
    expr_1061_wire_constant <= "00000000";
    expr_985_wire_constant <= "01110011";
    expr_989_wire_constant <= "01110100";
    expr_993_wire_constant <= "01100001";
    expr_997_wire_constant <= "01110010";
    array_obj_ref_1000_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1000_gather_scatter_ack_0 <= array_obj_ref_1000_gather_scatter_req_0;
      aggregated_sig <= expr_1001_wire_constant;
      array_obj_ref_1000_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1004_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1004_gather_scatter_ack_0 <= array_obj_ref_1004_gather_scatter_req_0;
      aggregated_sig <= expr_1005_wire_constant;
      array_obj_ref_1004_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1008_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1008_gather_scatter_ack_0 <= array_obj_ref_1008_gather_scatter_req_0;
      aggregated_sig <= expr_1009_wire_constant;
      array_obj_ref_1008_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1012_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1012_gather_scatter_ack_0 <= array_obj_ref_1012_gather_scatter_req_0;
      aggregated_sig <= expr_1013_wire_constant;
      array_obj_ref_1012_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1016_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1016_gather_scatter_ack_0 <= array_obj_ref_1016_gather_scatter_req_0;
      aggregated_sig <= expr_1017_wire_constant;
      array_obj_ref_1016_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1020_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1020_gather_scatter_ack_0 <= array_obj_ref_1020_gather_scatter_req_0;
      aggregated_sig <= expr_1021_wire_constant;
      array_obj_ref_1020_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1024_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1024_gather_scatter_ack_0 <= array_obj_ref_1024_gather_scatter_req_0;
      aggregated_sig <= expr_1025_wire_constant;
      array_obj_ref_1024_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1028_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1028_gather_scatter_ack_0 <= array_obj_ref_1028_gather_scatter_req_0;
      aggregated_sig <= expr_1029_wire_constant;
      array_obj_ref_1028_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1032_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1032_gather_scatter_ack_0 <= array_obj_ref_1032_gather_scatter_req_0;
      aggregated_sig <= expr_1033_wire_constant;
      array_obj_ref_1032_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1036_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1036_gather_scatter_ack_0 <= array_obj_ref_1036_gather_scatter_req_0;
      aggregated_sig <= expr_1037_wire_constant;
      array_obj_ref_1036_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1040_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1040_gather_scatter_ack_0 <= array_obj_ref_1040_gather_scatter_req_0;
      aggregated_sig <= expr_1041_wire_constant;
      array_obj_ref_1040_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1044_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1044_gather_scatter_ack_0 <= array_obj_ref_1044_gather_scatter_req_0;
      aggregated_sig <= expr_1045_wire_constant;
      array_obj_ref_1044_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1048_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1048_gather_scatter_ack_0 <= array_obj_ref_1048_gather_scatter_req_0;
      aggregated_sig <= expr_1049_wire_constant;
      array_obj_ref_1048_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1052_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1052_gather_scatter_ack_0 <= array_obj_ref_1052_gather_scatter_req_0;
      aggregated_sig <= expr_1053_wire_constant;
      array_obj_ref_1052_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1056_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1056_gather_scatter_ack_0 <= array_obj_ref_1056_gather_scatter_req_0;
      aggregated_sig <= expr_1057_wire_constant;
      array_obj_ref_1056_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_1060_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_1060_gather_scatter_ack_0 <= array_obj_ref_1060_gather_scatter_req_0;
      aggregated_sig <= expr_1061_wire_constant;
      array_obj_ref_1060_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_984_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_984_gather_scatter_ack_0 <= array_obj_ref_984_gather_scatter_req_0;
      aggregated_sig <= expr_985_wire_constant;
      array_obj_ref_984_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_988_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_988_gather_scatter_ack_0 <= array_obj_ref_988_gather_scatter_req_0;
      aggregated_sig <= expr_989_wire_constant;
      array_obj_ref_988_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_992_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_992_gather_scatter_ack_0 <= array_obj_ref_992_gather_scatter_req_0;
      aggregated_sig <= expr_993_wire_constant;
      array_obj_ref_992_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_996_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_996_gather_scatter_ack_0 <= array_obj_ref_996_gather_scatter_req_0;
      aggregated_sig <= expr_997_wire_constant;
      array_obj_ref_996_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_1052_store_0 array_obj_ref_1048_store_0 array_obj_ref_1000_store_0 array_obj_ref_1020_store_0 array_obj_ref_1044_store_0 array_obj_ref_1056_store_0 array_obj_ref_1060_store_0 array_obj_ref_1016_store_0 array_obj_ref_984_store_0 array_obj_ref_1036_store_0 array_obj_ref_1024_store_0 array_obj_ref_1012_store_0 array_obj_ref_996_store_0 array_obj_ref_1028_store_0 array_obj_ref_988_store_0 array_obj_ref_992_store_0 array_obj_ref_1040_store_0 array_obj_ref_1032_store_0 array_obj_ref_1008_store_0 array_obj_ref_1004_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(99 downto 0);
      signal data_in: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 19 downto 0);
      -- 
    begin -- 
      reqL(19) <= array_obj_ref_1052_store_0_req_0;
      reqL(18) <= array_obj_ref_1048_store_0_req_0;
      reqL(17) <= array_obj_ref_1000_store_0_req_0;
      reqL(16) <= array_obj_ref_1020_store_0_req_0;
      reqL(15) <= array_obj_ref_1044_store_0_req_0;
      reqL(14) <= array_obj_ref_1056_store_0_req_0;
      reqL(13) <= array_obj_ref_1060_store_0_req_0;
      reqL(12) <= array_obj_ref_1016_store_0_req_0;
      reqL(11) <= array_obj_ref_984_store_0_req_0;
      reqL(10) <= array_obj_ref_1036_store_0_req_0;
      reqL(9) <= array_obj_ref_1024_store_0_req_0;
      reqL(8) <= array_obj_ref_1012_store_0_req_0;
      reqL(7) <= array_obj_ref_996_store_0_req_0;
      reqL(6) <= array_obj_ref_1028_store_0_req_0;
      reqL(5) <= array_obj_ref_988_store_0_req_0;
      reqL(4) <= array_obj_ref_992_store_0_req_0;
      reqL(3) <= array_obj_ref_1040_store_0_req_0;
      reqL(2) <= array_obj_ref_1032_store_0_req_0;
      reqL(1) <= array_obj_ref_1008_store_0_req_0;
      reqL(0) <= array_obj_ref_1004_store_0_req_0;
      array_obj_ref_1052_store_0_ack_0 <= ackL(19);
      array_obj_ref_1048_store_0_ack_0 <= ackL(18);
      array_obj_ref_1000_store_0_ack_0 <= ackL(17);
      array_obj_ref_1020_store_0_ack_0 <= ackL(16);
      array_obj_ref_1044_store_0_ack_0 <= ackL(15);
      array_obj_ref_1056_store_0_ack_0 <= ackL(14);
      array_obj_ref_1060_store_0_ack_0 <= ackL(13);
      array_obj_ref_1016_store_0_ack_0 <= ackL(12);
      array_obj_ref_984_store_0_ack_0 <= ackL(11);
      array_obj_ref_1036_store_0_ack_0 <= ackL(10);
      array_obj_ref_1024_store_0_ack_0 <= ackL(9);
      array_obj_ref_1012_store_0_ack_0 <= ackL(8);
      array_obj_ref_996_store_0_ack_0 <= ackL(7);
      array_obj_ref_1028_store_0_ack_0 <= ackL(6);
      array_obj_ref_988_store_0_ack_0 <= ackL(5);
      array_obj_ref_992_store_0_ack_0 <= ackL(4);
      array_obj_ref_1040_store_0_ack_0 <= ackL(3);
      array_obj_ref_1032_store_0_ack_0 <= ackL(2);
      array_obj_ref_1008_store_0_ack_0 <= ackL(1);
      array_obj_ref_1004_store_0_ack_0 <= ackL(0);
      reqR(19) <= array_obj_ref_1052_store_0_req_1;
      reqR(18) <= array_obj_ref_1048_store_0_req_1;
      reqR(17) <= array_obj_ref_1000_store_0_req_1;
      reqR(16) <= array_obj_ref_1020_store_0_req_1;
      reqR(15) <= array_obj_ref_1044_store_0_req_1;
      reqR(14) <= array_obj_ref_1056_store_0_req_1;
      reqR(13) <= array_obj_ref_1060_store_0_req_1;
      reqR(12) <= array_obj_ref_1016_store_0_req_1;
      reqR(11) <= array_obj_ref_984_store_0_req_1;
      reqR(10) <= array_obj_ref_1036_store_0_req_1;
      reqR(9) <= array_obj_ref_1024_store_0_req_1;
      reqR(8) <= array_obj_ref_1012_store_0_req_1;
      reqR(7) <= array_obj_ref_996_store_0_req_1;
      reqR(6) <= array_obj_ref_1028_store_0_req_1;
      reqR(5) <= array_obj_ref_988_store_0_req_1;
      reqR(4) <= array_obj_ref_992_store_0_req_1;
      reqR(3) <= array_obj_ref_1040_store_0_req_1;
      reqR(2) <= array_obj_ref_1032_store_0_req_1;
      reqR(1) <= array_obj_ref_1008_store_0_req_1;
      reqR(0) <= array_obj_ref_1004_store_0_req_1;
      array_obj_ref_1052_store_0_ack_1 <= ackR(19);
      array_obj_ref_1048_store_0_ack_1 <= ackR(18);
      array_obj_ref_1000_store_0_ack_1 <= ackR(17);
      array_obj_ref_1020_store_0_ack_1 <= ackR(16);
      array_obj_ref_1044_store_0_ack_1 <= ackR(15);
      array_obj_ref_1056_store_0_ack_1 <= ackR(14);
      array_obj_ref_1060_store_0_ack_1 <= ackR(13);
      array_obj_ref_1016_store_0_ack_1 <= ackR(12);
      array_obj_ref_984_store_0_ack_1 <= ackR(11);
      array_obj_ref_1036_store_0_ack_1 <= ackR(10);
      array_obj_ref_1024_store_0_ack_1 <= ackR(9);
      array_obj_ref_1012_store_0_ack_1 <= ackR(8);
      array_obj_ref_996_store_0_ack_1 <= ackR(7);
      array_obj_ref_1028_store_0_ack_1 <= ackR(6);
      array_obj_ref_988_store_0_ack_1 <= ackR(5);
      array_obj_ref_992_store_0_ack_1 <= ackR(4);
      array_obj_ref_1040_store_0_ack_1 <= ackR(3);
      array_obj_ref_1032_store_0_ack_1 <= ackR(2);
      array_obj_ref_1008_store_0_ack_1 <= ackR(1);
      array_obj_ref_1004_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_1052_word_address_0 & array_obj_ref_1048_word_address_0 & array_obj_ref_1000_word_address_0 & array_obj_ref_1020_word_address_0 & array_obj_ref_1044_word_address_0 & array_obj_ref_1056_word_address_0 & array_obj_ref_1060_word_address_0 & array_obj_ref_1016_word_address_0 & array_obj_ref_984_word_address_0 & array_obj_ref_1036_word_address_0 & array_obj_ref_1024_word_address_0 & array_obj_ref_1012_word_address_0 & array_obj_ref_996_word_address_0 & array_obj_ref_1028_word_address_0 & array_obj_ref_988_word_address_0 & array_obj_ref_992_word_address_0 & array_obj_ref_1040_word_address_0 & array_obj_ref_1032_word_address_0 & array_obj_ref_1008_word_address_0 & array_obj_ref_1004_word_address_0;
      data_in <= array_obj_ref_1052_data_0 & array_obj_ref_1048_data_0 & array_obj_ref_1000_data_0 & array_obj_ref_1020_data_0 & array_obj_ref_1044_data_0 & array_obj_ref_1056_data_0 & array_obj_ref_1060_data_0 & array_obj_ref_1016_data_0 & array_obj_ref_984_data_0 & array_obj_ref_1036_data_0 & array_obj_ref_1024_data_0 & array_obj_ref_1012_data_0 & array_obj_ref_996_data_0 & array_obj_ref_1028_data_0 & array_obj_ref_988_data_0 & array_obj_ref_992_data_0 & array_obj_ref_1040_data_0 & array_obj_ref_1032_data_0 & array_obj_ref_1008_data_0 & array_obj_ref_1004_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 8,
        num_reqs => 20,
        tag_length => 5,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_19_sr_req(0),
          mack => memory_space_19_sr_ack(0),
          maddr => memory_space_19_sr_addr(4 downto 0),
          mdata => memory_space_19_sr_data(7 downto 0),
          mtag => memory_space_19_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 20,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_19_sc_req(0),
          mack => memory_space_19_sc_ack(0),
          mtag => memory_space_19_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_manager is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(3 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(3 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(3 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(3 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(7 downto 0);
    free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_ack_pipe_write_data : out  std_logic_vector(7 downto 0);
    free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
    start_output_port_lookup_pipe_write_req : out  std_logic_vector(0 downto 0);
    start_output_port_lookup_pipe_write_ack : in   std_logic_vector(0 downto 0);
    start_output_port_lookup_pipe_write_data : out  std_logic_vector(7 downto 0);
    start_wrapper_input_pipe_write_req : out  std_logic_vector(0 downto 0);
    start_wrapper_input_pipe_write_ack : in   std_logic_vector(0 downto 0);
    start_wrapper_input_pipe_write_data : out  std_logic_vector(7 downto 0);
    start_wrapper_output_pipe_write_req : out  std_logic_vector(0 downto 0);
    start_wrapper_output_pipe_write_ack : in   std_logic_vector(0 downto 0);
    start_wrapper_output_pipe_write_data : out  std_logic_vector(7 downto 0);
    global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity free_queue_manager;
architecture Default of free_queue_manager is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal free_queue_manager_CP_5336_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_1194_base_resize_ack_0 : boolean;
  signal type_cast_1230_inst_req_0 : boolean;
  signal binary_1178_inst_req_1 : boolean;
  signal simple_obj_ref_1150_inst_req_0 : boolean;
  signal call_stmt_1066_call_ack_0 : boolean;
  signal ptr_deref_1115_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1126_store_0_ack_0 : boolean;
  signal call_stmt_1066_call_req_1 : boolean;
  signal switch_stmt_1152_branch_default_req_0 : boolean;
  signal array_obj_ref_1225_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1233_base_resize_ack_0 : boolean;
  signal addr_of_1190_final_reg_req_0 : boolean;
  signal ptr_deref_1194_root_address_inst_req_0 : boolean;
  signal switch_stmt_1152_select_expr_0_req_1 : boolean;
  signal switch_stmt_1152_select_expr_0_req_0 : boolean;
  signal switch_stmt_1152_select_expr_1_ack_0 : boolean;
  signal simple_obj_ref_1150_inst_ack_0 : boolean;
  signal switch_stmt_1152_select_expr_0_ack_0 : boolean;
  signal addr_of_1190_final_reg_ack_0 : boolean;
  signal switch_stmt_1152_branch_0_req_0 : boolean;
  signal if_stmt_1180_branch_req_0 : boolean;
  signal ptr_deref_1104_store_0_ack_1 : boolean;
  signal ptr_deref_1137_store_0_req_1 : boolean;
  signal array_obj_ref_1225_offset_inst_req_0 : boolean;
  signal ptr_deref_1126_store_0_ack_1 : boolean;
  signal array_obj_ref_1225_index_0_resize_req_0 : boolean;
  signal binary_1178_inst_ack_1 : boolean;
  signal ptr_deref_1194_root_address_inst_ack_0 : boolean;
  signal type_cast_1230_inst_ack_0 : boolean;
  signal ptr_deref_1126_store_0_req_1 : boolean;
  signal binary_1221_inst_ack_1 : boolean;
  signal ptr_deref_1126_gather_scatter_req_0 : boolean;
  signal ptr_deref_1233_gather_scatter_req_0 : boolean;
  signal ptr_deref_1233_store_0_req_0 : boolean;
  signal array_obj_ref_1189_offset_inst_req_0 : boolean;
  signal call_stmt_1066_call_req_0 : boolean;
  signal ptr_deref_1137_store_0_req_0 : boolean;
  signal array_obj_ref_1225_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1104_store_0_req_1 : boolean;
  signal binary_1221_inst_req_1 : boolean;
  signal array_obj_ref_1189_index_0_rename_req_0 : boolean;
  signal binary_1221_inst_req_0 : boolean;
  signal ptr_deref_1194_addr_0_ack_0 : boolean;
  signal ptr_deref_1233_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1126_gather_scatter_ack_0 : boolean;
  signal switch_stmt_1152_select_expr_0_ack_1 : boolean;
  signal ptr_deref_1115_store_0_req_0 : boolean;
  signal addr_of_1226_final_reg_ack_0 : boolean;
  signal ptr_deref_1137_store_0_ack_0 : boolean;
  signal simple_obj_ref_1243_inst_req_0 : boolean;
  signal ptr_deref_1115_store_0_ack_0 : boolean;
  signal if_stmt_1180_branch_ack_1 : boolean;
  signal array_obj_ref_1189_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1189_root_address_inst_req_0 : boolean;
  signal ptr_deref_1137_store_0_ack_1 : boolean;
  signal call_stmt_1066_call_ack_1 : boolean;
  signal array_obj_ref_1225_root_address_inst_req_0 : boolean;
  signal ptr_deref_1115_gather_scatter_req_0 : boolean;
  signal switch_stmt_1152_select_expr_1_req_0 : boolean;
  signal ptr_deref_1233_root_address_inst_req_0 : boolean;
  signal if_stmt_1180_branch_ack_0 : boolean;
  signal ptr_deref_1233_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1189_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1233_base_resize_req_0 : boolean;
  signal array_obj_ref_1189_index_0_rename_ack_0 : boolean;
  signal simple_obj_ref_1277_inst_ack_0 : boolean;
  signal simple_obj_ref_1073_inst_ack_0 : boolean;
  signal binary_1178_inst_ack_0 : boolean;
  signal ptr_deref_1126_store_0_req_0 : boolean;
  signal ptr_deref_1104_store_0_ack_0 : boolean;
  signal array_obj_ref_1189_index_0_resize_req_0 : boolean;
  signal binary_1213_inst_ack_0 : boolean;
  signal binary_1213_inst_req_0 : boolean;
  signal simple_obj_ref_1277_inst_req_0 : boolean;
  signal ptr_deref_1104_store_0_req_0 : boolean;
  signal ptr_deref_1137_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1137_gather_scatter_req_0 : boolean;
  signal binary_1213_inst_ack_1 : boolean;
  signal binary_1213_inst_req_1 : boolean;
  signal ptr_deref_1104_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1104_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1225_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1225_index_0_rename_req_0 : boolean;
  signal if_stmt_1202_branch_ack_0 : boolean;
  signal ptr_deref_1233_addr_0_ack_0 : boolean;
  signal switch_stmt_1152_select_expr_1_req_1 : boolean;
  signal binary_1221_inst_ack_0 : boolean;
  signal switch_stmt_1152_select_expr_1_ack_1 : boolean;
  signal switch_stmt_1152_branch_1_req_0 : boolean;
  signal ptr_deref_1194_base_resize_req_0 : boolean;
  signal array_obj_ref_1189_offset_inst_ack_0 : boolean;
  signal switch_stmt_1152_branch_0_ack_1 : boolean;
  signal ptr_deref_1194_addr_0_req_0 : boolean;
  signal addr_of_1226_final_reg_req_0 : boolean;
  signal array_obj_ref_1225_root_address_inst_ack_0 : boolean;
  signal switch_stmt_1152_branch_1_ack_1 : boolean;
  signal switch_stmt_1152_branch_default_ack_0 : boolean;
  signal ptr_deref_1115_store_0_req_1 : boolean;
  signal ptr_deref_1115_store_0_ack_1 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal binary_1178_inst_req_0 : boolean;
  signal simple_obj_ref_1073_inst_req_0 : boolean;
  signal if_stmt_1202_branch_ack_1 : boolean;
  signal simple_obj_ref_1253_inst_ack_0 : boolean;
  signal ptr_deref_1233_addr_0_req_0 : boolean;
  signal if_stmt_1202_branch_req_0 : boolean;
  signal simple_obj_ref_1253_inst_req_0 : boolean;
  signal ptr_deref_1233_store_0_ack_1 : boolean;
  signal ptr_deref_1233_store_0_req_1 : boolean;
  signal binary_1200_inst_ack_1 : boolean;
  signal simple_obj_ref_1093_inst_ack_0 : boolean;
  signal simple_obj_ref_1093_inst_req_0 : boolean;
  signal binary_1200_inst_req_1 : boolean;
  signal binary_1200_inst_ack_0 : boolean;
  signal binary_1200_inst_req_0 : boolean;
  signal ptr_deref_1194_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1194_gather_scatter_req_0 : boolean;
  signal ptr_deref_1194_load_0_ack_1 : boolean;
  signal ptr_deref_1194_load_0_req_1 : boolean;
  signal simple_obj_ref_1264_inst_ack_0 : boolean;
  signal ptr_deref_1233_store_0_ack_0 : boolean;
  signal simple_obj_ref_1264_inst_req_0 : boolean;
  signal simple_obj_ref_1083_inst_ack_0 : boolean;
  signal ptr_deref_1194_load_0_ack_0 : boolean;
  signal simple_obj_ref_1083_inst_req_0 : boolean;
  signal ptr_deref_1194_load_0_req_0 : boolean;
  signal simple_obj_ref_1243_inst_ack_0 : boolean;
  signal binary_1283_inst_req_0 : boolean;
  signal binary_1283_inst_ack_0 : boolean;
  signal binary_1283_inst_req_1 : boolean;
  signal binary_1283_inst_ack_1 : boolean;
  signal if_stmt_1285_branch_req_0 : boolean;
  signal if_stmt_1285_branch_ack_1 : boolean;
  signal if_stmt_1285_branch_ack_0 : boolean;
  signal binary_1304_inst_req_0 : boolean;
  signal binary_1304_inst_ack_0 : boolean;
  signal binary_1304_inst_req_1 : boolean;
  signal binary_1304_inst_ack_1 : boolean;
  signal binary_1310_inst_req_0 : boolean;
  signal binary_1310_inst_ack_0 : boolean;
  signal binary_1310_inst_req_1 : boolean;
  signal binary_1310_inst_ack_1 : boolean;
  signal binary_1316_inst_req_0 : boolean;
  signal binary_1316_inst_ack_0 : boolean;
  signal binary_1316_inst_req_1 : boolean;
  signal binary_1316_inst_ack_1 : boolean;
  signal binary_1321_inst_req_0 : boolean;
  signal binary_1321_inst_ack_0 : boolean;
  signal binary_1321_inst_req_1 : boolean;
  signal binary_1321_inst_ack_1 : boolean;
  signal if_stmt_1323_branch_req_0 : boolean;
  signal if_stmt_1323_branch_ack_1 : boolean;
  signal if_stmt_1323_branch_ack_0 : boolean;
  signal type_cast_1332_inst_req_0 : boolean;
  signal type_cast_1332_inst_ack_0 : boolean;
  signal binary_1336_inst_req_0 : boolean;
  signal binary_1336_inst_ack_0 : boolean;
  signal binary_1336_inst_req_1 : boolean;
  signal binary_1336_inst_ack_1 : boolean;
  signal if_stmt_1338_branch_req_0 : boolean;
  signal if_stmt_1338_branch_ack_1 : boolean;
  signal if_stmt_1338_branch_ack_0 : boolean;
  signal array_obj_ref_1355_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1355_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1355_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1355_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1355_offset_inst_req_0 : boolean;
  signal array_obj_ref_1355_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1355_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1355_root_address_inst_ack_0 : boolean;
  signal addr_of_1356_final_reg_req_0 : boolean;
  signal addr_of_1356_final_reg_ack_0 : boolean;
  signal ptr_deref_1359_base_resize_req_0 : boolean;
  signal ptr_deref_1359_base_resize_ack_0 : boolean;
  signal ptr_deref_1359_root_address_inst_req_0 : boolean;
  signal ptr_deref_1359_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1359_addr_0_req_0 : boolean;
  signal ptr_deref_1359_addr_0_ack_0 : boolean;
  signal ptr_deref_1359_gather_scatter_req_0 : boolean;
  signal ptr_deref_1359_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1359_store_0_req_0 : boolean;
  signal ptr_deref_1359_store_0_ack_0 : boolean;
  signal ptr_deref_1359_store_0_req_1 : boolean;
  signal ptr_deref_1359_store_0_ack_1 : boolean;
  signal type_cast_1166_inst_req_0 : boolean;
  signal type_cast_1166_inst_ack_0 : boolean;
  signal phi_stmt_1163_req_0 : boolean;
  signal phi_stmt_1163_req_1 : boolean;
  signal phi_stmt_1163_ack_0 : boolean;
  signal phi_stmt_1292_req_1 : boolean;
  signal type_cast_1295_inst_req_0 : boolean;
  signal type_cast_1295_inst_ack_0 : boolean;
  signal phi_stmt_1292_req_0 : boolean;
  signal phi_stmt_1292_ack_0 : boolean;
  signal phi_stmt_1345_req_1 : boolean;
  signal type_cast_1348_inst_req_0 : boolean;
  signal type_cast_1348_inst_ack_0 : boolean;
  signal phi_stmt_1345_req_0 : boolean;
  signal phi_stmt_1345_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  free_queue_manager_CP_5336: Block -- control-path 
    signal cp_elements: BooleanArray(260 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    call_stmt_1066_call_req_0 <= cp_elements(0);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(48);
    cp_elements(3) <= OrReduce(cp_elements(238) & cp_elements(242));
    cp_elements(4) <= OrReduce(cp_elements(84) & cp_elements(244));
    cp_elements(5) <= OrReduce(cp_elements(116) & cp_elements(246));
    cp_elements(6) <= cp_elements(149);
    simple_obj_ref_1243_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= OrReduce(cp_elements(248) & cp_elements(252));
    cp_elements(8) <= cp_elements(189);
    cp_elements(9) <= OrReduce(cp_elements(198) & cp_elements(254));
    cp_elements(10) <= OrReduce(cp_elements(256) & cp_elements(260));
    cp_elements(11) <= call_stmt_1066_call_ack_0;
    call_stmt_1066_call_req_1 <= cp_elements(11);
    cp_elements(12) <= call_stmt_1066_call_ack_1;
    simple_obj_ref_1073_inst_req_0 <= cp_elements(12);
    cp_elements(13) <= simple_obj_ref_1073_inst_ack_0;
    simple_obj_ref_1083_inst_req_0 <= cp_elements(13);
    cp_elements(14) <= simple_obj_ref_1083_inst_ack_0;
    simple_obj_ref_1093_inst_req_0 <= cp_elements(14);
    cp_elements(15) <= simple_obj_ref_1093_inst_ack_0;
    cp_elements(16) <= cp_elements(15);
    cp_elements(17) <= cp_elements(16);
    cpelement_group_18 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(17) & cp_elements(20));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(18),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1104_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(16);
    cp_elements(20) <= cp_elements(16);
    cp_elements(21) <= ptr_deref_1104_gather_scatter_ack_0;
    ptr_deref_1104_store_0_req_0 <= cp_elements(21);
    cp_elements(22) <= ptr_deref_1104_store_0_ack_0;
    cp_elements(23) <= cp_elements(22);
    ptr_deref_1104_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= ptr_deref_1104_store_0_ack_1;
    cp_elements(25) <= cp_elements(16);
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(25) & cp_elements(28));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1115_gather_scatter_req_0 <= cp_elements(26);
    cp_elements(27) <= cp_elements(16);
    cp_elements(28) <= cp_elements(16);
    cp_elements(29) <= ptr_deref_1115_gather_scatter_ack_0;
    ptr_deref_1115_store_0_req_0 <= cp_elements(29);
    cp_elements(30) <= ptr_deref_1115_store_0_ack_0;
    cp_elements(31) <= cp_elements(30);
    ptr_deref_1115_store_0_req_1 <= cp_elements(31);
    cp_elements(32) <= ptr_deref_1115_store_0_ack_1;
    cp_elements(33) <= cp_elements(16);
    cpelement_group_34 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(33) & cp_elements(36));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(34),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1126_gather_scatter_req_0 <= cp_elements(34);
    cp_elements(35) <= cp_elements(16);
    cp_elements(36) <= cp_elements(16);
    cp_elements(37) <= ptr_deref_1126_gather_scatter_ack_0;
    ptr_deref_1126_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= ptr_deref_1126_store_0_ack_0;
    cp_elements(39) <= cp_elements(38);
    ptr_deref_1126_store_0_req_1 <= cp_elements(39);
    cp_elements(40) <= ptr_deref_1126_store_0_ack_1;
    cp_elements(41) <= cp_elements(16);
    cpelement_group_42 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(38) & cp_elements(41) & cp_elements(44));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(42),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1137_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= cp_elements(16);
    cp_elements(44) <= cp_elements(16);
    cp_elements(45) <= ptr_deref_1137_gather_scatter_ack_0;
    ptr_deref_1137_store_0_req_0 <= cp_elements(45);
    cp_elements(46) <= ptr_deref_1137_store_0_ack_0;
    ptr_deref_1137_store_0_req_1 <= cp_elements(46);
    cp_elements(47) <= ptr_deref_1137_store_0_ack_1;
    cpelement_group_48 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(24) & cp_elements(27) & cp_elements(32) & cp_elements(35) & cp_elements(40) & cp_elements(43) & cp_elements(47));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(48),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(49) <= simple_obj_ref_1150_inst_ack_0;
    cp_elements(50) <= cp_elements(49);
    cp_elements(51) <= false;
    cp_elements(52) <= cp_elements(51);
    cp_elements(53) <= cp_elements(49);
    cp_elements(54) <= cp_elements(53);
    cp_elements(55) <= cp_elements(54);
    switch_stmt_1152_select_expr_0_req_0 <= cp_elements(55);
    cp_elements(56) <= switch_stmt_1152_select_expr_0_ack_0;
    switch_stmt_1152_select_expr_0_req_1 <= cp_elements(56);
    cp_elements(57) <= switch_stmt_1152_select_expr_0_ack_1;
    switch_stmt_1152_branch_0_req_0 <= cp_elements(57);
    cp_elements(58) <= cp_elements(54);
    switch_stmt_1152_select_expr_1_req_0 <= cp_elements(58);
    cp_elements(59) <= switch_stmt_1152_select_expr_1_ack_0;
    switch_stmt_1152_select_expr_1_req_1 <= cp_elements(59);
    cp_elements(60) <= switch_stmt_1152_select_expr_1_ack_1;
    switch_stmt_1152_branch_1_req_0 <= cp_elements(60);
    cpelement_group_61 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(57) & cp_elements(60));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(61),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    switch_stmt_1152_branch_default_req_0 <= cp_elements(61);
    cp_elements(62) <= cp_elements(61);
    cp_elements(63) <= cp_elements(62);
    cp_elements(64) <= switch_stmt_1152_branch_0_ack_1;
    phi_stmt_1163_req_1 <= cp_elements(64);
    cp_elements(65) <= cp_elements(62);
    cp_elements(66) <= switch_stmt_1152_branch_1_ack_1;
    simple_obj_ref_1277_inst_req_0 <= cp_elements(66);
    cp_elements(67) <= cp_elements(62);
    cp_elements(68) <= switch_stmt_1152_branch_default_ack_0;
    cp_elements(69) <= cp_elements(3);
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(75));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1178_inst_req_0 <= cp_elements(70);
    cp_elements(71) <= cp_elements(69);
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(73) & cp_elements(74));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1174_inst_req_0 <= cp_elements(72);
    cp_elements(73) <= cp_elements(69);
    cp_elements(74) <= cp_elements(69);
    cp_elements(75) <= type_cast_1174_inst_ack_0;
    cp_elements(76) <= binary_1178_inst_ack_0;
    binary_1178_inst_req_1 <= cp_elements(76);
    cp_elements(77) <= binary_1178_inst_ack_1;
    cp_elements(78) <= cp_elements(77);
    cp_elements(79) <= false;
    cp_elements(80) <= cp_elements(79);
    cp_elements(81) <= cp_elements(77);
    if_stmt_1180_branch_req_0 <= cp_elements(81);
    cp_elements(82) <= cp_elements(81);
    cp_elements(83) <= cp_elements(82);
    cp_elements(84) <= if_stmt_1180_branch_ack_1;
    cp_elements(85) <= cp_elements(82);
    cp_elements(86) <= if_stmt_1180_branch_ack_0;
    simple_obj_ref_1264_inst_req_0 <= cp_elements(86);
    cp_elements(87) <= cp_elements(4);
    cpelement_group_88 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(94));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(88),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_1190_final_reg_req_0 <= cp_elements(88);
    cp_elements(89) <= cp_elements(87);
    cp_elements(90) <= cp_elements(87);
    array_obj_ref_1189_index_0_resize_req_0 <= cp_elements(90);
    cp_elements(91) <= array_obj_ref_1189_index_0_resize_ack_0;
    array_obj_ref_1189_index_0_rename_req_0 <= cp_elements(91);
    cp_elements(92) <= array_obj_ref_1189_index_0_rename_ack_0;
    array_obj_ref_1189_offset_inst_req_0 <= cp_elements(92);
    cp_elements(93) <= array_obj_ref_1189_offset_inst_ack_0;
    array_obj_ref_1189_root_address_inst_req_0 <= cp_elements(93);
    cp_elements(94) <= array_obj_ref_1189_root_address_inst_ack_0;
    cp_elements(95) <= addr_of_1190_final_reg_ack_0;
    cpelement_group_96 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(95) & cp_elements(100));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(96),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1194_load_0_req_0 <= cp_elements(96);
    cp_elements(97) <= cp_elements(95);
    ptr_deref_1194_base_resize_req_0 <= cp_elements(97);
    cp_elements(98) <= ptr_deref_1194_base_resize_ack_0;
    ptr_deref_1194_root_address_inst_req_0 <= cp_elements(98);
    cp_elements(99) <= ptr_deref_1194_root_address_inst_ack_0;
    ptr_deref_1194_addr_0_req_0 <= cp_elements(99);
    cp_elements(100) <= ptr_deref_1194_addr_0_ack_0;
    cp_elements(101) <= ptr_deref_1194_load_0_ack_0;
    ptr_deref_1194_load_0_req_1 <= cp_elements(101);
    cp_elements(102) <= ptr_deref_1194_load_0_ack_1;
    ptr_deref_1194_gather_scatter_req_0 <= cp_elements(102);
    cp_elements(103) <= ptr_deref_1194_gather_scatter_ack_0;
    cpelement_group_104 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(103) & cp_elements(105));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(104),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1200_inst_req_0 <= cp_elements(104);
    cp_elements(105) <= cp_elements(87);
    cp_elements(106) <= binary_1200_inst_ack_0;
    binary_1200_inst_req_1 <= cp_elements(106);
    cp_elements(107) <= binary_1200_inst_ack_1;
    cp_elements(108) <= cp_elements(107);
    cp_elements(109) <= false;
    cp_elements(110) <= cp_elements(109);
    cp_elements(111) <= cp_elements(107);
    if_stmt_1202_branch_req_0 <= cp_elements(111);
    cp_elements(112) <= cp_elements(111);
    cp_elements(113) <= cp_elements(112);
    cp_elements(114) <= if_stmt_1202_branch_ack_1;
    cp_elements(115) <= cp_elements(112);
    cp_elements(116) <= if_stmt_1202_branch_ack_0;
    cp_elements(117) <= cp_elements(5);
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(119) & cp_elements(120));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1213_inst_req_0 <= cp_elements(118);
    cp_elements(119) <= cp_elements(117);
    cp_elements(120) <= cp_elements(117);
    cp_elements(121) <= binary_1213_inst_ack_0;
    binary_1213_inst_req_1 <= cp_elements(121);
    cp_elements(122) <= binary_1213_inst_ack_1;
    type_cast_1166_inst_req_0 <= cp_elements(122);
    cp_elements(123) <= cp_elements(114);
    cpelement_group_124 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(126));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(124),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1221_inst_req_0 <= cp_elements(124);
    cp_elements(125) <= cp_elements(123);
    cp_elements(126) <= cp_elements(123);
    cp_elements(127) <= binary_1221_inst_ack_0;
    binary_1221_inst_req_1 <= cp_elements(127);
    cp_elements(128) <= binary_1221_inst_ack_1;
    array_obj_ref_1225_index_0_resize_req_0 <= cp_elements(128);
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(130) & cp_elements(134));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_1226_final_reg_req_0 <= cp_elements(129);
    cp_elements(130) <= cp_elements(123);
    cp_elements(131) <= array_obj_ref_1225_index_0_resize_ack_0;
    array_obj_ref_1225_index_0_rename_req_0 <= cp_elements(131);
    cp_elements(132) <= array_obj_ref_1225_index_0_rename_ack_0;
    array_obj_ref_1225_offset_inst_req_0 <= cp_elements(132);
    cp_elements(133) <= array_obj_ref_1225_offset_inst_ack_0;
    array_obj_ref_1225_root_address_inst_req_0 <= cp_elements(133);
    cp_elements(134) <= array_obj_ref_1225_root_address_inst_ack_0;
    cp_elements(135) <= addr_of_1226_final_reg_ack_0;
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(135) & cp_elements(137));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1230_inst_req_0 <= cp_elements(136);
    cp_elements(137) <= cp_elements(123);
    cp_elements(138) <= type_cast_1230_inst_ack_0;
    cp_elements(139) <= cp_elements(123);
    cpelement_group_140 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(145));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(140),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1233_gather_scatter_req_0 <= cp_elements(140);
    cp_elements(141) <= cp_elements(123);
    cp_elements(142) <= cp_elements(141);
    ptr_deref_1233_base_resize_req_0 <= cp_elements(142);
    cp_elements(143) <= ptr_deref_1233_base_resize_ack_0;
    ptr_deref_1233_root_address_inst_req_0 <= cp_elements(143);
    cp_elements(144) <= ptr_deref_1233_root_address_inst_ack_0;
    ptr_deref_1233_addr_0_req_0 <= cp_elements(144);
    cp_elements(145) <= ptr_deref_1233_addr_0_ack_0;
    cp_elements(146) <= ptr_deref_1233_gather_scatter_ack_0;
    ptr_deref_1233_store_0_req_0 <= cp_elements(146);
    cp_elements(147) <= ptr_deref_1233_store_0_ack_0;
    ptr_deref_1233_store_0_req_1 <= cp_elements(147);
    cp_elements(148) <= ptr_deref_1233_store_0_ack_1;
    cpelement_group_149 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(138) & cp_elements(148));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(149),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(150) <= simple_obj_ref_1243_inst_ack_0;
    simple_obj_ref_1253_inst_req_0 <= cp_elements(150);
    cp_elements(151) <= simple_obj_ref_1253_inst_ack_0;
    cp_elements(152) <= simple_obj_ref_1264_inst_ack_0;
    cp_elements(153) <= simple_obj_ref_1277_inst_ack_0;
    cp_elements(154) <= cp_elements(153);
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(157));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1283_inst_req_0 <= cp_elements(155);
    cp_elements(156) <= cp_elements(154);
    cp_elements(157) <= cp_elements(154);
    cp_elements(158) <= binary_1283_inst_ack_0;
    binary_1283_inst_req_1 <= cp_elements(158);
    cp_elements(159) <= binary_1283_inst_ack_1;
    cp_elements(160) <= cp_elements(159);
    cp_elements(161) <= false;
    cp_elements(162) <= cp_elements(161);
    cp_elements(163) <= cp_elements(159);
    if_stmt_1285_branch_req_0 <= cp_elements(163);
    cp_elements(164) <= cp_elements(163);
    cp_elements(165) <= cp_elements(164);
    cp_elements(166) <= if_stmt_1285_branch_ack_1;
    phi_stmt_1292_req_1 <= cp_elements(166);
    cp_elements(167) <= cp_elements(164);
    cp_elements(168) <= if_stmt_1285_branch_ack_0;
    phi_stmt_1345_req_1 <= cp_elements(168);
    cp_elements(169) <= cp_elements(7);
    cpelement_group_170 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(171) & cp_elements(172));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(170),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1304_inst_req_0 <= cp_elements(170);
    cp_elements(171) <= cp_elements(169);
    cp_elements(172) <= cp_elements(169);
    cp_elements(173) <= binary_1304_inst_ack_0;
    binary_1304_inst_req_1 <= cp_elements(173);
    cp_elements(174) <= binary_1304_inst_ack_1;
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(176) & cp_elements(177));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1310_inst_req_0 <= cp_elements(175);
    cp_elements(176) <= cp_elements(169);
    cp_elements(177) <= cp_elements(169);
    cp_elements(178) <= binary_1310_inst_ack_0;
    binary_1310_inst_req_1 <= cp_elements(178);
    cp_elements(179) <= binary_1310_inst_ack_1;
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(174) & cp_elements(181));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1316_inst_req_0 <= cp_elements(180);
    cp_elements(181) <= cp_elements(169);
    cp_elements(182) <= binary_1316_inst_ack_0;
    binary_1316_inst_req_1 <= cp_elements(182);
    cp_elements(183) <= binary_1316_inst_ack_1;
    cpelement_group_184 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(183) & cp_elements(185) & cp_elements(186));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(184),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1321_inst_req_0 <= cp_elements(184);
    cp_elements(185) <= cp_elements(169);
    cp_elements(186) <= cp_elements(169);
    cp_elements(187) <= binary_1321_inst_ack_0;
    binary_1321_inst_req_1 <= cp_elements(187);
    cp_elements(188) <= binary_1321_inst_ack_1;
    cpelement_group_189 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(188));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(189),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(190) <= cp_elements(8);
    cp_elements(191) <= false;
    cp_elements(192) <= cp_elements(191);
    cp_elements(193) <= cp_elements(8);
    if_stmt_1323_branch_req_0 <= cp_elements(193);
    cp_elements(194) <= cp_elements(193);
    cp_elements(195) <= cp_elements(194);
    cp_elements(196) <= if_stmt_1323_branch_ack_1;
    type_cast_1295_inst_req_0 <= cp_elements(196);
    cp_elements(197) <= cp_elements(194);
    cp_elements(198) <= if_stmt_1323_branch_ack_0;
    cp_elements(199) <= cp_elements(9);
    cpelement_group_200 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(201) & cp_elements(205));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1336_inst_req_0 <= cp_elements(200);
    cp_elements(201) <= cp_elements(199);
    cpelement_group_202 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(204));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(202),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1332_inst_req_0 <= cp_elements(202);
    cp_elements(203) <= cp_elements(199);
    cp_elements(204) <= cp_elements(199);
    cp_elements(205) <= type_cast_1332_inst_ack_0;
    cp_elements(206) <= binary_1336_inst_ack_0;
    binary_1336_inst_req_1 <= cp_elements(206);
    cp_elements(207) <= binary_1336_inst_ack_1;
    cp_elements(208) <= cp_elements(207);
    cp_elements(209) <= false;
    cp_elements(210) <= cp_elements(209);
    cp_elements(211) <= cp_elements(207);
    if_stmt_1338_branch_req_0 <= cp_elements(211);
    cp_elements(212) <= cp_elements(211);
    cp_elements(213) <= cp_elements(212);
    cp_elements(214) <= if_stmt_1338_branch_ack_1;
    type_cast_1348_inst_req_0 <= cp_elements(214);
    cp_elements(215) <= cp_elements(212);
    cp_elements(216) <= if_stmt_1338_branch_ack_0;
    cp_elements(217) <= cp_elements(10);
    cpelement_group_218 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(219) & cp_elements(224));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(218),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_1356_final_reg_req_0 <= cp_elements(218);
    cp_elements(219) <= cp_elements(217);
    cp_elements(220) <= cp_elements(217);
    array_obj_ref_1355_index_0_resize_req_0 <= cp_elements(220);
    cp_elements(221) <= array_obj_ref_1355_index_0_resize_ack_0;
    array_obj_ref_1355_index_0_rename_req_0 <= cp_elements(221);
    cp_elements(222) <= array_obj_ref_1355_index_0_rename_ack_0;
    array_obj_ref_1355_offset_inst_req_0 <= cp_elements(222);
    cp_elements(223) <= array_obj_ref_1355_offset_inst_ack_0;
    array_obj_ref_1355_root_address_inst_req_0 <= cp_elements(223);
    cp_elements(224) <= array_obj_ref_1355_root_address_inst_ack_0;
    cp_elements(225) <= addr_of_1356_final_reg_ack_0;
    cp_elements(226) <= cp_elements(217);
    cpelement_group_227 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(225) & cp_elements(226) & cp_elements(231));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(227),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1359_gather_scatter_req_0 <= cp_elements(227);
    cp_elements(228) <= cp_elements(225);
    ptr_deref_1359_base_resize_req_0 <= cp_elements(228);
    cp_elements(229) <= ptr_deref_1359_base_resize_ack_0;
    ptr_deref_1359_root_address_inst_req_0 <= cp_elements(229);
    cp_elements(230) <= ptr_deref_1359_root_address_inst_ack_0;
    ptr_deref_1359_addr_0_req_0 <= cp_elements(230);
    cp_elements(231) <= ptr_deref_1359_addr_0_ack_0;
    cp_elements(232) <= ptr_deref_1359_gather_scatter_ack_0;
    ptr_deref_1359_store_0_req_0 <= cp_elements(232);
    cp_elements(233) <= ptr_deref_1359_store_0_ack_0;
    ptr_deref_1359_store_0_req_1 <= cp_elements(233);
    cp_elements(234) <= ptr_deref_1359_store_0_ack_1;
    cp_elements(235) <= OrReduce(cp_elements(2) & cp_elements(68) & cp_elements(151) & cp_elements(152) & cp_elements(216) & cp_elements(234));
    cp_elements(236) <= cp_elements(235);
    simple_obj_ref_1150_inst_req_0 <= cp_elements(236);
    cp_elements(237) <= false;
    cp_elements(238) <= cp_elements(237);
    cp_elements(239) <= type_cast_1166_inst_ack_0;
    phi_stmt_1163_req_0 <= cp_elements(239);
    cp_elements(240) <= OrReduce(cp_elements(64) & cp_elements(239));
    cp_elements(241) <= cp_elements(240);
    cp_elements(242) <= phi_stmt_1163_ack_0;
    cp_elements(243) <= false;
    cp_elements(244) <= cp_elements(243);
    cp_elements(245) <= false;
    cp_elements(246) <= cp_elements(245);
    cp_elements(247) <= false;
    cp_elements(248) <= cp_elements(247);
    cp_elements(249) <= type_cast_1295_inst_ack_0;
    phi_stmt_1292_req_0 <= cp_elements(249);
    cp_elements(250) <= OrReduce(cp_elements(166) & cp_elements(249));
    cp_elements(251) <= cp_elements(250);
    cp_elements(252) <= phi_stmt_1292_ack_0;
    cp_elements(253) <= false;
    cp_elements(254) <= cp_elements(253);
    cp_elements(255) <= false;
    cp_elements(256) <= cp_elements(255);
    cp_elements(257) <= type_cast_1348_inst_ack_0;
    phi_stmt_1345_req_0 <= cp_elements(257);
    cp_elements(258) <= OrReduce(cp_elements(168) & cp_elements(257));
    cp_elements(259) <= cp_elements(258);
    cp_elements(260) <= phi_stmt_1345_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1189_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1189_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1189_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1189_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1225_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1225_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1225_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1225_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1355_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1355_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1355_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1355_root_address : std_logic_vector(2 downto 0);
    signal expr_1154_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1154_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_1157_wire_constant : std_logic_vector(7 downto 0);
    signal expr_1157_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal i3x_x044_1292 : std_logic_vector(31 downto 0);
    signal i3x_x0x_xlcssa53_1345 : std_logic_vector(31 downto 0);
    signal iNsTr_11_1124 : std_logic_vector(31 downto 0);
    signal iNsTr_13_1135 : std_logic_vector(31 downto 0);
    signal iNsTr_16_1148 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1163 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1072 : std_logic_vector(31 downto 0);
    signal iNsTr_20_1275 : std_logic_vector(31 downto 0);
    signal iNsTr_23_1263 : std_logic_vector(31 downto 0);
    signal iNsTr_26_1311 : std_logic_vector(31 downto 0);
    signal iNsTr_31_1242 : std_logic_vector(31 downto 0);
    signal iNsTr_33_1252 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1082 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1092 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1102 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1113 : std_logic_vector(31 downto 0);
    signal ptr_deref_1104_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1104_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1104_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1115_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1115_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1115_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1126_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1126_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1126_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1137_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1137_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1137_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1194_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1194_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1194_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1194_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1194_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1233_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1233_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1233_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1233_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1233_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1233_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1359_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1359_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1359_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1359_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1359_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1359_word_offset_0 : std_logic_vector(2 downto 0);
    signal simple_obj_ref_1188_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_1188_scaled : std_logic_vector(2 downto 0);
    signal simple_obj_ref_1224_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1224_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1354_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_1354_scaled : std_logic_vector(2 downto 0);
    signal tmp10_1179 : std_logic_vector(0 downto 0);
    signal tmp12_1191 : std_logic_vector(31 downto 0);
    signal tmp13_1195 : std_logic_vector(7 downto 0);
    signal tmp14_1201 : std_logic_vector(0 downto 0);
    signal tmp16_1222 : std_logic_vector(31 downto 0);
    signal tmp17_1227 : std_logic_vector(31 downto 0);
    signal tmp18_1231 : std_logic_vector(31 downto 0);
    signal tmp21_1214 : std_logic_vector(31 downto 0);
    signal tmp28_1278 : std_logic_vector(31 downto 0);
    signal tmp31_1317 : std_logic_vector(31 downto 0);
    signal tmp3243_1284 : std_logic_vector(0 downto 0);
    signal tmp32_1322 : std_logic_vector(0 downto 0);
    signal tmp36_1337 : std_logic_vector(0 downto 0);
    signal tmp38_1357 : std_logic_vector(31 downto 0);
    signal tmp50_1305 : std_logic_vector(31 downto 0);
    signal tmp6_1151 : std_logic_vector(7 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1085_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1095_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1139_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1166_wire : std_logic_vector(31 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1174_wire : std_logic_vector(31 downto 0);
    signal type_cast_1177_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1199_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1212_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1220_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1235_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1282_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1295_wire : std_logic_vector(31 downto 0);
    signal type_cast_1298_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1309_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1315_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1332_wire : std_logic_vector(31 downto 0);
    signal type_cast_1335_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1348_wire : std_logic_vector(31 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1361_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1189_offset_scale_factor_0 <= "001";
    array_obj_ref_1189_resized_base_address <= "000";
    array_obj_ref_1225_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1225_resized_base_address <= "00000000000";
    array_obj_ref_1355_offset_scale_factor_0 <= "001";
    array_obj_ref_1355_resized_base_address <= "000";
    expr_1154_wire_constant <= "00000010";
    expr_1157_wire_constant <= "00000001";
    iNsTr_11_1124 <= "00000000000000000000000000000010";
    iNsTr_13_1135 <= "00000000000000000000000000000011";
    iNsTr_16_1148 <= "00000000000000000000000000000000";
    iNsTr_1_1072 <= "00000000000000000000000000000000";
    iNsTr_20_1275 <= "00000000000000000000000000000000";
    iNsTr_23_1263 <= "00000000000000000000000000000000";
    iNsTr_31_1242 <= "00000000000000000000000000000000";
    iNsTr_33_1252 <= "00000000000000000000000000000000";
    iNsTr_3_1082 <= "00000000000000000000000000000000";
    iNsTr_5_1092 <= "00000000000000000000000000000000";
    iNsTr_7_1102 <= "00000000000000000000000000000000";
    iNsTr_9_1113 <= "00000000000000000000000000000001";
    ptr_deref_1104_word_address_0 <= "000";
    ptr_deref_1115_word_address_0 <= "001";
    ptr_deref_1126_word_address_0 <= "010";
    ptr_deref_1137_word_address_0 <= "011";
    ptr_deref_1194_word_offset_0 <= "000";
    ptr_deref_1233_word_offset_0 <= "000";
    ptr_deref_1359_word_offset_0 <= "000";
    type_cast_1075_wire_constant <= "00000001";
    type_cast_1085_wire_constant <= "00000001";
    type_cast_1095_wire_constant <= "00000001";
    type_cast_1106_wire_constant <= "00000001";
    type_cast_1117_wire_constant <= "00000001";
    type_cast_1128_wire_constant <= "00000001";
    type_cast_1139_wire_constant <= "00000001";
    type_cast_1169_wire_constant <= "00000000000000000000000000000000";
    type_cast_1177_wire_constant <= "00000000000000000000000000000100";
    type_cast_1199_wire_constant <= "00000001";
    type_cast_1212_wire_constant <= "00000000000000000000000000000001";
    type_cast_1220_wire_constant <= "00000000000000000000000000001000";
    type_cast_1235_wire_constant <= "00000000";
    type_cast_1245_wire_constant <= "00000011";
    type_cast_1266_wire_constant <= "00000100";
    type_cast_1282_wire_constant <= "00000000000000000000000100000000";
    type_cast_1298_wire_constant <= "00000000000000000000000000000000";
    type_cast_1303_wire_constant <= "00000000000000000000000000001000";
    type_cast_1309_wire_constant <= "00000000000000000000000000000001";
    type_cast_1315_wire_constant <= "00000000000000000000001000000000";
    type_cast_1335_wire_constant <= "00000000000000000000000000000100";
    type_cast_1351_wire_constant <= "00000000000000000000000000000000";
    type_cast_1361_wire_constant <= "00000001";
    phi_stmt_1163: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1166_wire & type_cast_1169_wire_constant;
      req <= phi_stmt_1163_req_0 & phi_stmt_1163_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1163_ack_0,
          idata => idata,
          odata => iNsTr_18_1163,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1163
    phi_stmt_1292: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1295_wire & type_cast_1298_wire_constant;
      req <= phi_stmt_1292_req_0 & phi_stmt_1292_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1292_ack_0,
          idata => idata,
          odata => i3x_x044_1292,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1292
    phi_stmt_1345: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1348_wire & type_cast_1351_wire_constant;
      req <= phi_stmt_1345_req_0 & phi_stmt_1345_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1345_ack_0,
          idata => idata,
          odata => i3x_x0x_xlcssa53_1345,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1345
    addr_of_1190_final_reg: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1189_root_address, dout => tmp12_1191, req => addr_of_1190_final_reg_req_0, ack => addr_of_1190_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1226_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1225_root_address, dout => tmp17_1227, req => addr_of_1226_final_reg_req_0, ack => addr_of_1226_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1356_final_reg: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1355_root_address, dout => tmp38_1357, req => addr_of_1356_final_reg_req_0, ack => addr_of_1356_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1189_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => iNsTr_18_1163, dout => simple_obj_ref_1188_resized, req => array_obj_ref_1189_index_0_resize_req_0, ack => array_obj_ref_1189_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1189_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_1188_scaled, dout => array_obj_ref_1189_final_offset, req => array_obj_ref_1189_offset_inst_req_0, ack => array_obj_ref_1189_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1225_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp16_1222, dout => simple_obj_ref_1224_resized, req => array_obj_ref_1225_index_0_resize_req_0, ack => array_obj_ref_1225_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1225_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1224_scaled, dout => array_obj_ref_1225_final_offset, req => array_obj_ref_1225_offset_inst_req_0, ack => array_obj_ref_1225_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1355_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => i3x_x0x_xlcssa53_1345, dout => simple_obj_ref_1354_resized, req => array_obj_ref_1355_index_0_resize_req_0, ack => array_obj_ref_1355_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1355_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_1354_scaled, dout => array_obj_ref_1355_final_offset, req => array_obj_ref_1355_offset_inst_req_0, ack => array_obj_ref_1355_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1194_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp12_1191, dout => ptr_deref_1194_resized_base_address, req => ptr_deref_1194_base_resize_req_0, ack => ptr_deref_1194_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1233_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp12_1191, dout => ptr_deref_1233_resized_base_address, req => ptr_deref_1233_base_resize_req_0, ack => ptr_deref_1233_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1359_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp38_1357, dout => ptr_deref_1359_resized_base_address, req => ptr_deref_1359_base_resize_req_0, ack => ptr_deref_1359_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1166_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp21_1214, dout => type_cast_1166_wire, req => type_cast_1166_inst_req_0, ack => type_cast_1166_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1174_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_18_1163, dout => type_cast_1174_wire, req => type_cast_1174_inst_req_0, ack => type_cast_1174_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1230_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_1227, dout => tmp18_1231, req => type_cast_1230_inst_req_0, ack => type_cast_1230_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1295_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_26_1311, dout => type_cast_1295_wire, req => type_cast_1295_inst_req_0, ack => type_cast_1295_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1332_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_26_1311, dout => type_cast_1332_wire, req => type_cast_1332_inst_req_0, ack => type_cast_1332_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1348_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_26_1311, dout => type_cast_1348_wire, req => type_cast_1348_inst_req_0, ack => type_cast_1348_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1189_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_1189_index_0_rename_ack_0 <= array_obj_ref_1189_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1188_resized;
      simple_obj_ref_1188_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_1189_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_1189_root_address_inst_ack_0 <= array_obj_ref_1189_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1189_final_offset;
      array_obj_ref_1189_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_1225_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1225_index_0_rename_ack_0 <= array_obj_ref_1225_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1224_resized;
      simple_obj_ref_1224_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1225_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1225_root_address_inst_ack_0 <= array_obj_ref_1225_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1225_final_offset;
      array_obj_ref_1225_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1355_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_1355_index_0_rename_ack_0 <= array_obj_ref_1355_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1354_resized;
      simple_obj_ref_1354_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_1355_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_1355_root_address_inst_ack_0 <= array_obj_ref_1355_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1355_final_offset;
      array_obj_ref_1355_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1104_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1104_gather_scatter_ack_0 <= ptr_deref_1104_gather_scatter_req_0;
      aggregated_sig <= type_cast_1106_wire_constant;
      ptr_deref_1104_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1115_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1115_gather_scatter_ack_0 <= ptr_deref_1115_gather_scatter_req_0;
      aggregated_sig <= type_cast_1117_wire_constant;
      ptr_deref_1115_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1126_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1126_gather_scatter_ack_0 <= ptr_deref_1126_gather_scatter_req_0;
      aggregated_sig <= type_cast_1128_wire_constant;
      ptr_deref_1126_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1137_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1137_gather_scatter_ack_0 <= ptr_deref_1137_gather_scatter_req_0;
      aggregated_sig <= type_cast_1139_wire_constant;
      ptr_deref_1137_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1194_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1194_addr_0_ack_0 <= ptr_deref_1194_addr_0_req_0;
      aggregated_sig <= ptr_deref_1194_root_address;
      ptr_deref_1194_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1194_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1194_gather_scatter_ack_0 <= ptr_deref_1194_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1194_data_0;
      tmp13_1195 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1194_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1194_root_address_inst_ack_0 <= ptr_deref_1194_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1194_resized_base_address;
      ptr_deref_1194_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1233_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1233_addr_0_ack_0 <= ptr_deref_1233_addr_0_req_0;
      aggregated_sig <= ptr_deref_1233_root_address;
      ptr_deref_1233_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1233_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1233_gather_scatter_ack_0 <= ptr_deref_1233_gather_scatter_req_0;
      aggregated_sig <= type_cast_1235_wire_constant;
      ptr_deref_1233_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1233_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1233_root_address_inst_ack_0 <= ptr_deref_1233_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1233_resized_base_address;
      ptr_deref_1233_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1359_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1359_addr_0_ack_0 <= ptr_deref_1359_addr_0_req_0;
      aggregated_sig <= ptr_deref_1359_root_address;
      ptr_deref_1359_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1359_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1359_gather_scatter_ack_0 <= ptr_deref_1359_gather_scatter_req_0;
      aggregated_sig <= type_cast_1361_wire_constant;
      ptr_deref_1359_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1359_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1359_root_address_inst_ack_0 <= ptr_deref_1359_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1359_resized_base_address;
      ptr_deref_1359_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    if_stmt_1180_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp10_1179;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1180_branch_req_0,
          ack0 => if_stmt_1180_branch_ack_0,
          ack1 => if_stmt_1180_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1202_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp14_1201;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1202_branch_req_0,
          ack0 => if_stmt_1202_branch_ack_0,
          ack1 => if_stmt_1202_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1285_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp3243_1284;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1285_branch_req_0,
          ack0 => if_stmt_1285_branch_ack_0,
          ack1 => if_stmt_1285_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1323_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp32_1322;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1323_branch_req_0,
          ack0 => if_stmt_1323_branch_ack_0,
          ack1 => if_stmt_1323_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1338_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp36_1337;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1338_branch_req_0,
          ack0 => if_stmt_1338_branch_ack_0,
          ack1 => if_stmt_1338_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1152_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1154_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1152_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_1152_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1152_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1157_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1152_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_1152_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1152_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_1154_wire_constant_cmp & expr_1157_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1152_branch_default_req_0,
          ack0 => switch_stmt_1152_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_1336_inst binary_1178_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1332_wire & type_cast_1174_wire;
      tmp36_1337 <= data_out(1 downto 1);
      tmp10_1179 <= data_out(0 downto 0);
      reqL(1) <= binary_1336_inst_req_0;
      reqL(0) <= binary_1178_inst_req_0;
      binary_1336_inst_ack_0 <= ackL(1);
      binary_1178_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1336_inst_req_1;
      reqR(0) <= binary_1178_inst_req_1;
      binary_1336_inst_ack_1 <= ackR(1);
      binary_1178_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_1200_inst switch_stmt_1152_select_expr_1 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_1195 & tmp6_1151;
      tmp14_1201 <= data_out(1 downto 1);
      expr_1157_wire_constant_cmp <= data_out(0 downto 0);
      reqL(1) <= binary_1200_inst_req_0;
      reqL(0) <= switch_stmt_1152_select_expr_1_req_0;
      binary_1200_inst_ack_0 <= ackL(1);
      switch_stmt_1152_select_expr_1_ack_0 <= ackL(0);
      reqR(1) <= binary_1200_inst_req_1;
      reqR(0) <= switch_stmt_1152_select_expr_1_req_1;
      binary_1200_inst_ack_1 <= ackR(1);
      switch_stmt_1152_select_expr_1_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1213_inst binary_1310_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_18_1163 & i3x_x044_1292;
      tmp21_1214 <= data_out(63 downto 32);
      iNsTr_26_1311 <= data_out(31 downto 0);
      reqL(1) <= binary_1213_inst_req_0;
      reqL(0) <= binary_1310_inst_req_0;
      binary_1213_inst_ack_0 <= ackL(1);
      binary_1310_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1213_inst_req_1;
      reqR(0) <= binary_1310_inst_req_1;
      binary_1213_inst_ack_1 <= ackR(1);
      binary_1310_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1221_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_18_1163;
      tmp16_1222 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1221_inst_req_0,
          ackL => binary_1221_inst_ack_0,
          reqR => binary_1221_inst_req_1,
          ackR => binary_1221_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_1283_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp28_1278;
      tmp3243_1284 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000100000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1283_inst_req_0,
          ackL => binary_1283_inst_ack_0,
          reqR => binary_1283_inst_req_1,
          ackR => binary_1283_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_1304_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i3x_x044_1292;
      tmp50_1305 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1304_inst_req_0,
          ackL => binary_1304_inst_ack_0,
          reqR => binary_1304_inst_req_1,
          ackR => binary_1304_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_1316_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp50_1305;
      tmp31_1317 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000001000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1316_inst_req_0,
          ackL => binary_1316_inst_ack_0,
          reqR => binary_1316_inst_req_1,
          ackR => binary_1316_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_1321_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp28_1278 & tmp31_1317;
      tmp32_1322 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1321_inst_req_0,
          ackL => binary_1321_inst_ack_0,
          reqR => binary_1321_inst_req_1,
          ackR => binary_1321_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : switch_stmt_1152_select_expr_0 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_1151;
      expr_1154_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1152_select_expr_0_req_0,
          ackL => switch_stmt_1152_select_expr_0_ack_0,
          reqR => switch_stmt_1152_select_expr_0_req_1,
          ackR => switch_stmt_1152_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared load operator group (0) : ptr_deref_1194_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1194_load_0_req_0;
      ptr_deref_1194_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1194_load_0_req_1;
      ptr_deref_1194_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1194_word_address_0;
      ptr_deref_1194_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 3,  num_reqs => 1,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(2 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1233_store_0 ptr_deref_1104_store_0 ptr_deref_1359_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(8 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1233_store_0_req_0;
      reqL(1) <= ptr_deref_1104_store_0_req_0;
      reqL(0) <= ptr_deref_1359_store_0_req_0;
      ptr_deref_1233_store_0_ack_0 <= ackL(2);
      ptr_deref_1104_store_0_ack_0 <= ackL(1);
      ptr_deref_1359_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1233_store_0_req_1;
      reqR(1) <= ptr_deref_1104_store_0_req_1;
      reqR(0) <= ptr_deref_1359_store_0_req_1;
      ptr_deref_1233_store_0_ack_1 <= ackR(2);
      ptr_deref_1104_store_0_ack_1 <= ackR(1);
      ptr_deref_1359_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1233_word_address_0 & ptr_deref_1104_word_address_0 & ptr_deref_1359_word_address_0;
      data_in <= ptr_deref_1233_data_0 & ptr_deref_1104_data_0 & ptr_deref_1359_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(3),
          mack => memory_space_2_sr_ack(3),
          maddr => memory_space_2_sr_addr(11 downto 9),
          mdata => memory_space_2_sr_data(31 downto 24),
          mtag => memory_space_2_sr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(3),
          mack => memory_space_2_sc_ack(3),
          mtag => memory_space_2_sc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1115_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1115_store_0_req_0;
      ptr_deref_1115_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1115_store_0_req_1;
      ptr_deref_1115_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1115_word_address_0;
      data_in <= ptr_deref_1115_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(2),
          mack => memory_space_2_sr_ack(2),
          maddr => memory_space_2_sr_addr(8 downto 6),
          mdata => memory_space_2_sr_data(23 downto 16),
          mtag => memory_space_2_sr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(2),
          mack => memory_space_2_sc_ack(2),
          mtag => memory_space_2_sc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_1126_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1126_store_0_req_0;
      ptr_deref_1126_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1126_store_0_req_1;
      ptr_deref_1126_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1126_word_address_0;
      data_in <= ptr_deref_1126_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(1),
          mack => memory_space_2_sr_ack(1),
          maddr => memory_space_2_sr_addr(5 downto 3),
          mdata => memory_space_2_sr_data(15 downto 8),
          mtag => memory_space_2_sr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(1),
          mack => memory_space_2_sc_ack(1),
          mtag => memory_space_2_sc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_1137_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1137_store_0_req_0;
      ptr_deref_1137_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1137_store_0_req_1;
      ptr_deref_1137_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1137_word_address_0;
      data_in <= ptr_deref_1137_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(2 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : simple_obj_ref_1150_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1150_inst_req_0;
      simple_obj_ref_1150_inst_ack_0 <= ack(0);
      tmp6_1151 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_request_pipe_read_req(0),
          oack => free_queue_request_pipe_read_ack(0),
          odata => free_queue_request_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1277_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1277_inst_req_0;
      simple_obj_ref_1277_inst_ack_0 <= ack(0);
      tmp28_1278 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_put_pipe_read_req(0),
          oack => free_queue_put_pipe_read_ack(0),
          odata => free_queue_put_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_1073_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1073_inst_req_0;
      simple_obj_ref_1073_inst_ack_0 <= ack(0);
      data_in <= type_cast_1075_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => start_wrapper_input_pipe_write_req(0),
          oack => start_wrapper_input_pipe_write_ack(0),
          odata => start_wrapper_input_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_1083_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1083_inst_req_0;
      simple_obj_ref_1083_inst_ack_0 <= ack(0);
      data_in <= type_cast_1085_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => start_wrapper_output_pipe_write_req(0),
          oack => start_wrapper_output_pipe_write_ack(0),
          odata => start_wrapper_output_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_1093_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1093_inst_req_0;
      simple_obj_ref_1093_inst_ack_0 <= ack(0);
      data_in <= type_cast_1095_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => start_output_port_lookup_pipe_write_req(0),
          oack => start_output_port_lookup_pipe_write_ack(0),
          odata => start_output_port_lookup_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : simple_obj_ref_1243_inst simple_obj_ref_1264_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_1243_inst_req_0;
      req(0) <= simple_obj_ref_1264_inst_req_0;
      simple_obj_ref_1243_inst_ack_0 <= ack(1);
      simple_obj_ref_1264_inst_ack_0 <= ack(0);
      data_in <= type_cast_1245_wire_constant & type_cast_1266_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 2,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_ack_pipe_write_req(0),
          oack => free_queue_ack_pipe_write_ack(0),
          odata => free_queue_ack_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : simple_obj_ref_1253_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1253_inst_req_0;
      simple_obj_ref_1253_inst_ack_0 <= ack(0);
      data_in <= tmp18_1231;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_get_pipe_write_req(0),
          oack => free_queue_get_pipe_write_ack(0),
          odata => free_queue_get_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1066_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1066_call_req_0;
      call_stmt_1066_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1066_call_req_1;
      call_stmt_1066_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => global_storage_initializer_x_call_reqs(0),
          ackR => global_storage_initializer_x_call_acks(0),
          tagR => global_storage_initializer_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => global_storage_initializer_x_return_acks(0), -- cross-over
          ackL => global_storage_initializer_x_return_reqs(0), -- cross-over
          tagL => global_storage_initializer_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity global_storage_initializer_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    default_initializer_foo_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_foo_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_foo_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_foo_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_foo_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_foo_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr12_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr12_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr12_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr12_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr12_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr12_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr13_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr13_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr13_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr13_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr13_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr13_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr10_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr10_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr10_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr10_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr10_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr10_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr11_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr11_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr11_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr11_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr11_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr11_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr14_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr14_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr14_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr14_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr14_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr14_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr15_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr15_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr15_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr15_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr15_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr15_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr9_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr9_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr9_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr9_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr9_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr9_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity global_storage_initializer_x;
architecture Default of global_storage_initializer_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal global_storage_initializer_x_xCP_5007_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_1369_call_req_0 : boolean;
  signal call_stmt_1368_call_req_0 : boolean;
  signal call_stmt_1371_call_req_1 : boolean;
  signal call_stmt_1368_call_ack_1 : boolean;
  signal call_stmt_1368_call_ack_0 : boolean;
  signal call_stmt_1368_call_req_1 : boolean;
  signal call_stmt_1370_call_req_0 : boolean;
  signal call_stmt_1369_call_ack_0 : boolean;
  signal call_stmt_1369_call_req_1 : boolean;
  signal call_stmt_1372_call_ack_1 : boolean;
  signal call_stmt_1372_call_req_0 : boolean;
  signal call_stmt_1375_call_req_0 : boolean;
  signal call_stmt_1375_call_ack_0 : boolean;
  signal call_stmt_1372_call_ack_0 : boolean;
  signal call_stmt_1373_call_req_1 : boolean;
  signal call_stmt_1369_call_ack_1 : boolean;
  signal call_stmt_1373_call_ack_1 : boolean;
  signal call_stmt_1374_call_req_1 : boolean;
  signal call_stmt_1374_call_ack_0 : boolean;
  signal call_stmt_1372_call_req_1 : boolean;
  signal call_stmt_1374_call_ack_1 : boolean;
  signal call_stmt_1370_call_req_1 : boolean;
  signal call_stmt_1370_call_ack_1 : boolean;
  signal call_stmt_1371_call_req_0 : boolean;
  signal call_stmt_1371_call_ack_0 : boolean;
  signal call_stmt_1370_call_ack_0 : boolean;
  signal call_stmt_1375_call_req_1 : boolean;
  signal call_stmt_1375_call_ack_1 : boolean;
  signal call_stmt_1373_call_req_0 : boolean;
  signal call_stmt_1373_call_ack_0 : boolean;
  signal call_stmt_1376_call_req_0 : boolean;
  signal call_stmt_1376_call_ack_0 : boolean;
  signal call_stmt_1377_call_req_1 : boolean;
  signal call_stmt_1377_call_ack_1 : boolean;
  signal call_stmt_1379_call_ack_0 : boolean;
  signal call_stmt_1379_call_req_1 : boolean;
  signal call_stmt_1379_call_ack_1 : boolean;
  signal call_stmt_1379_call_req_0 : boolean;
  signal call_stmt_1377_call_req_0 : boolean;
  signal call_stmt_1377_call_ack_0 : boolean;
  signal call_stmt_1378_call_ack_1 : boolean;
  signal call_stmt_1378_call_ack_0 : boolean;
  signal call_stmt_1378_call_req_1 : boolean;
  signal call_stmt_1380_call_req_0 : boolean;
  signal call_stmt_1376_call_req_1 : boolean;
  signal call_stmt_1376_call_ack_1 : boolean;
  signal call_stmt_1378_call_req_0 : boolean;
  signal call_stmt_1374_call_req_0 : boolean;
  signal call_stmt_1371_call_ack_1 : boolean;
  signal call_stmt_1380_call_ack_0 : boolean;
  signal call_stmt_1380_call_req_1 : boolean;
  signal call_stmt_1380_call_ack_1 : boolean;
  signal call_stmt_1381_call_req_0 : boolean;
  signal call_stmt_1381_call_ack_0 : boolean;
  signal call_stmt_1381_call_req_1 : boolean;
  signal call_stmt_1381_call_ack_1 : boolean;
  signal call_stmt_1382_call_req_0 : boolean;
  signal call_stmt_1382_call_ack_0 : boolean;
  signal call_stmt_1382_call_req_1 : boolean;
  signal call_stmt_1382_call_ack_1 : boolean;
  signal call_stmt_1383_call_req_0 : boolean;
  signal call_stmt_1383_call_ack_0 : boolean;
  signal call_stmt_1383_call_req_1 : boolean;
  signal call_stmt_1383_call_ack_1 : boolean;
  signal call_stmt_1384_call_req_0 : boolean;
  signal call_stmt_1384_call_ack_0 : boolean;
  signal call_stmt_1384_call_req_1 : boolean;
  signal call_stmt_1384_call_ack_1 : boolean;
  signal call_stmt_1385_call_req_0 : boolean;
  signal call_stmt_1385_call_ack_0 : boolean;
  signal call_stmt_1385_call_req_1 : boolean;
  signal call_stmt_1385_call_ack_1 : boolean;
  signal call_stmt_1386_call_req_0 : boolean;
  signal call_stmt_1386_call_ack_0 : boolean;
  signal call_stmt_1386_call_req_1 : boolean;
  signal call_stmt_1386_call_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  global_storage_initializer_x_xCP_5007: Block -- control-path 
    signal cp_elements: BooleanArray(58 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(58);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(58), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    call_stmt_1368_call_req_0 <= cp_elements(1);
    cp_elements(2) <= call_stmt_1368_call_ack_0;
    call_stmt_1368_call_req_1 <= cp_elements(2);
    cp_elements(3) <= call_stmt_1368_call_ack_1;
    cp_elements(4) <= cp_elements(0);
    call_stmt_1369_call_req_0 <= cp_elements(4);
    cp_elements(5) <= call_stmt_1369_call_ack_0;
    call_stmt_1369_call_req_1 <= cp_elements(5);
    cp_elements(6) <= call_stmt_1369_call_ack_1;
    cp_elements(7) <= cp_elements(0);
    call_stmt_1370_call_req_0 <= cp_elements(7);
    cp_elements(8) <= call_stmt_1370_call_ack_0;
    call_stmt_1370_call_req_1 <= cp_elements(8);
    cp_elements(9) <= call_stmt_1370_call_ack_1;
    cp_elements(10) <= cp_elements(0);
    call_stmt_1371_call_req_0 <= cp_elements(10);
    cp_elements(11) <= call_stmt_1371_call_ack_0;
    call_stmt_1371_call_req_1 <= cp_elements(11);
    cp_elements(12) <= call_stmt_1371_call_ack_1;
    cp_elements(13) <= cp_elements(0);
    call_stmt_1372_call_req_0 <= cp_elements(13);
    cp_elements(14) <= call_stmt_1372_call_ack_0;
    call_stmt_1372_call_req_1 <= cp_elements(14);
    cp_elements(15) <= call_stmt_1372_call_ack_1;
    cp_elements(16) <= cp_elements(0);
    call_stmt_1373_call_req_0 <= cp_elements(16);
    cp_elements(17) <= call_stmt_1373_call_ack_0;
    call_stmt_1373_call_req_1 <= cp_elements(17);
    cp_elements(18) <= call_stmt_1373_call_ack_1;
    cp_elements(19) <= cp_elements(0);
    call_stmt_1374_call_req_0 <= cp_elements(19);
    cp_elements(20) <= call_stmt_1374_call_ack_0;
    call_stmt_1374_call_req_1 <= cp_elements(20);
    cp_elements(21) <= call_stmt_1374_call_ack_1;
    cp_elements(22) <= cp_elements(0);
    call_stmt_1375_call_req_0 <= cp_elements(22);
    cp_elements(23) <= call_stmt_1375_call_ack_0;
    call_stmt_1375_call_req_1 <= cp_elements(23);
    cp_elements(24) <= call_stmt_1375_call_ack_1;
    cp_elements(25) <= cp_elements(0);
    call_stmt_1376_call_req_0 <= cp_elements(25);
    cp_elements(26) <= call_stmt_1376_call_ack_0;
    call_stmt_1376_call_req_1 <= cp_elements(26);
    cp_elements(27) <= call_stmt_1376_call_ack_1;
    cp_elements(28) <= cp_elements(0);
    call_stmt_1377_call_req_0 <= cp_elements(28);
    cp_elements(29) <= call_stmt_1377_call_ack_0;
    call_stmt_1377_call_req_1 <= cp_elements(29);
    cp_elements(30) <= call_stmt_1377_call_ack_1;
    cp_elements(31) <= cp_elements(0);
    call_stmt_1378_call_req_0 <= cp_elements(31);
    cp_elements(32) <= call_stmt_1378_call_ack_0;
    call_stmt_1378_call_req_1 <= cp_elements(32);
    cp_elements(33) <= call_stmt_1378_call_ack_1;
    cp_elements(34) <= cp_elements(0);
    call_stmt_1379_call_req_0 <= cp_elements(34);
    cp_elements(35) <= call_stmt_1379_call_ack_0;
    call_stmt_1379_call_req_1 <= cp_elements(35);
    cp_elements(36) <= call_stmt_1379_call_ack_1;
    cp_elements(37) <= cp_elements(0);
    call_stmt_1380_call_req_0 <= cp_elements(37);
    cp_elements(38) <= call_stmt_1380_call_ack_0;
    call_stmt_1380_call_req_1 <= cp_elements(38);
    cp_elements(39) <= call_stmt_1380_call_ack_1;
    cp_elements(40) <= cp_elements(0);
    call_stmt_1381_call_req_0 <= cp_elements(40);
    cp_elements(41) <= call_stmt_1381_call_ack_0;
    call_stmt_1381_call_req_1 <= cp_elements(41);
    cp_elements(42) <= call_stmt_1381_call_ack_1;
    cp_elements(43) <= cp_elements(0);
    call_stmt_1382_call_req_0 <= cp_elements(43);
    cp_elements(44) <= call_stmt_1382_call_ack_0;
    call_stmt_1382_call_req_1 <= cp_elements(44);
    cp_elements(45) <= call_stmt_1382_call_ack_1;
    cp_elements(46) <= cp_elements(0);
    call_stmt_1383_call_req_0 <= cp_elements(46);
    cp_elements(47) <= call_stmt_1383_call_ack_0;
    call_stmt_1383_call_req_1 <= cp_elements(47);
    cp_elements(48) <= call_stmt_1383_call_ack_1;
    cp_elements(49) <= cp_elements(0);
    call_stmt_1384_call_req_0 <= cp_elements(49);
    cp_elements(50) <= call_stmt_1384_call_ack_0;
    call_stmt_1384_call_req_1 <= cp_elements(50);
    cp_elements(51) <= call_stmt_1384_call_ack_1;
    cp_elements(52) <= cp_elements(0);
    call_stmt_1385_call_req_0 <= cp_elements(52);
    cp_elements(53) <= call_stmt_1385_call_ack_0;
    call_stmt_1385_call_req_1 <= cp_elements(53);
    cp_elements(54) <= call_stmt_1385_call_ack_1;
    cp_elements(55) <= cp_elements(0);
    call_stmt_1386_call_req_0 <= cp_elements(55);
    cp_elements(56) <= call_stmt_1386_call_ack_0;
    call_stmt_1386_call_req_1 <= cp_elements(56);
    cp_elements(57) <= call_stmt_1386_call_ack_1;
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(18 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(6) & cp_elements(9) & cp_elements(12) & cp_elements(15) & cp_elements(18) & cp_elements(21) & cp_elements(24) & cp_elements(27) & cp_elements(30) & cp_elements(33) & cp_elements(36) & cp_elements(39) & cp_elements(42) & cp_elements(45) & cp_elements(48) & cp_elements(51) & cp_elements(54) & cp_elements(57));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_1368_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1368_call_req_0;
      call_stmt_1368_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1368_call_req_1;
      call_stmt_1368_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr_call_reqs(0),
          ackR => default_initializer_xx_xstr_call_acks(0),
          tagR => default_initializer_xx_xstr_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1369_call 
    CallGroup1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1369_call_req_0;
      call_stmt_1369_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1369_call_req_1;
      call_stmt_1369_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr1_call_reqs(0),
          ackR => default_initializer_xx_xstr1_call_acks(0),
          tagR => default_initializer_xx_xstr1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr1_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr1_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1370_call 
    CallGroup2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1370_call_req_0;
      call_stmt_1370_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1370_call_req_1;
      call_stmt_1370_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr2_call_reqs(0),
          ackR => default_initializer_xx_xstr2_call_acks(0),
          tagR => default_initializer_xx_xstr2_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr2_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr2_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr2_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1371_call 
    CallGroup3: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1371_call_req_0;
      call_stmt_1371_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1371_call_req_1;
      call_stmt_1371_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr3_call_reqs(0),
          ackR => default_initializer_xx_xstr3_call_acks(0),
          tagR => default_initializer_xx_xstr3_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr3_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr3_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr3_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1372_call 
    CallGroup4: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1372_call_req_0;
      call_stmt_1372_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1372_call_req_1;
      call_stmt_1372_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr4_call_reqs(0),
          ackR => default_initializer_xx_xstr4_call_acks(0),
          tagR => default_initializer_xx_xstr4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr4_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr4_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1373_call 
    CallGroup5: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1373_call_req_0;
      call_stmt_1373_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1373_call_req_1;
      call_stmt_1373_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr5_call_reqs(0),
          ackR => default_initializer_xx_xstr5_call_acks(0),
          tagR => default_initializer_xx_xstr5_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr5_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr5_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr5_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1374_call 
    CallGroup6: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1374_call_req_0;
      call_stmt_1374_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1374_call_req_1;
      call_stmt_1374_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr6_call_reqs(0),
          ackR => default_initializer_xx_xstr6_call_acks(0),
          tagR => default_initializer_xx_xstr6_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr6_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr6_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr6_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1375_call 
    CallGroup7: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1375_call_req_0;
      call_stmt_1375_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1375_call_req_1;
      call_stmt_1375_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr7_call_reqs(0),
          ackR => default_initializer_xx_xstr7_call_acks(0),
          tagR => default_initializer_xx_xstr7_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr7_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr7_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr7_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_1376_call 
    CallGroup8: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1376_call_req_0;
      call_stmt_1376_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1376_call_req_1;
      call_stmt_1376_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr8_call_reqs(0),
          ackR => default_initializer_xx_xstr8_call_acks(0),
          tagR => default_initializer_xx_xstr8_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr8_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr8_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr8_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- shared call operator group (9) : call_stmt_1377_call 
    CallGroup9: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1377_call_req_0;
      call_stmt_1377_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1377_call_req_1;
      call_stmt_1377_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr9_call_reqs(0),
          ackR => default_initializer_xx_xstr9_call_acks(0),
          tagR => default_initializer_xx_xstr9_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr9_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr9_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr9_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 9
    -- shared call operator group (10) : call_stmt_1378_call 
    CallGroup10: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1378_call_req_0;
      call_stmt_1378_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1378_call_req_1;
      call_stmt_1378_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr10_call_reqs(0),
          ackR => default_initializer_xx_xstr10_call_acks(0),
          tagR => default_initializer_xx_xstr10_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr10_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr10_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr10_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 10
    -- shared call operator group (11) : call_stmt_1379_call 
    CallGroup11: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1379_call_req_0;
      call_stmt_1379_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1379_call_req_1;
      call_stmt_1379_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_free_queue_call_reqs(0),
          ackR => default_initializer_free_queue_call_acks(0),
          tagR => default_initializer_free_queue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_free_queue_return_acks(0), -- cross-over
          ackL => default_initializer_free_queue_return_reqs(0), -- cross-over
          tagL => default_initializer_free_queue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 11
    -- shared call operator group (12) : call_stmt_1380_call 
    CallGroup12: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1380_call_req_0;
      call_stmt_1380_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1380_call_req_1;
      call_stmt_1380_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_free_queue_ram_call_reqs(0),
          ackR => default_initializer_free_queue_ram_call_acks(0),
          tagR => default_initializer_free_queue_ram_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_free_queue_ram_return_acks(0), -- cross-over
          ackL => default_initializer_free_queue_ram_return_reqs(0), -- cross-over
          tagL => default_initializer_free_queue_ram_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 12
    -- shared call operator group (13) : call_stmt_1381_call 
    CallGroup13: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1381_call_req_0;
      call_stmt_1381_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1381_call_req_1;
      call_stmt_1381_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_foo_call_reqs(0),
          ackR => default_initializer_foo_call_acks(0),
          tagR => default_initializer_foo_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_foo_return_acks(0), -- cross-over
          ackL => default_initializer_foo_return_reqs(0), -- cross-over
          tagL => default_initializer_foo_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 13
    -- shared call operator group (14) : call_stmt_1382_call 
    CallGroup14: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1382_call_req_0;
      call_stmt_1382_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1382_call_req_1;
      call_stmt_1382_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr11_call_reqs(0),
          ackR => default_initializer_xx_xstr11_call_acks(0),
          tagR => default_initializer_xx_xstr11_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr11_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr11_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr11_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 14
    -- shared call operator group (15) : call_stmt_1383_call 
    CallGroup15: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1383_call_req_0;
      call_stmt_1383_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1383_call_req_1;
      call_stmt_1383_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr12_call_reqs(0),
          ackR => default_initializer_xx_xstr12_call_acks(0),
          tagR => default_initializer_xx_xstr12_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr12_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr12_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr12_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 15
    -- shared call operator group (16) : call_stmt_1384_call 
    CallGroup16: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1384_call_req_0;
      call_stmt_1384_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1384_call_req_1;
      call_stmt_1384_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr13_call_reqs(0),
          ackR => default_initializer_xx_xstr13_call_acks(0),
          tagR => default_initializer_xx_xstr13_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr13_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr13_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr13_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 16
    -- shared call operator group (17) : call_stmt_1385_call 
    CallGroup17: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1385_call_req_0;
      call_stmt_1385_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1385_call_req_1;
      call_stmt_1385_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr14_call_reqs(0),
          ackR => default_initializer_xx_xstr14_call_acks(0),
          tagR => default_initializer_xx_xstr14_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr14_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr14_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr14_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 17
    -- shared call operator group (18) : call_stmt_1386_call 
    CallGroup18: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1386_call_req_0;
      call_stmt_1386_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1386_call_req_1;
      call_stmt_1386_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr15_call_reqs(0),
          ackR => default_initializer_xx_xstr15_call_acks(0),
          tagR => default_initializer_xx_xstr15_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr15_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr15_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr15_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 18
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity output_port_lookup is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    op_lut_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    op_lut_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    op_lut_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    op_lut_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    start_output_port_lookup_pipe_read_req : out  std_logic_vector(0 downto 0);
    start_output_port_lookup_pipe_read_ack : in   std_logic_vector(0 downto 0);
    start_output_port_lookup_pipe_read_data : in   std_logic_vector(7 downto 0);
    out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity output_port_lookup;
architecture Default of output_port_lookup is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal output_port_lookup_CP_6603_start: Boolean;
  -- links between control-path and data-path
  signal binary_1459_inst_req_1 : boolean;
  signal type_cast_1464_inst_req_0 : boolean;
  signal simple_obj_ref_1409_inst_ack_0 : boolean;
  signal binary_1447_inst_req_0 : boolean;
  signal simple_obj_ref_1409_inst_req_0 : boolean;
  signal simple_obj_ref_1418_inst_req_0 : boolean;
  signal simple_obj_ref_1418_inst_ack_0 : boolean;
  signal type_cast_1441_inst_req_0 : boolean;
  signal binary_1486_inst_req_0 : boolean;
  signal binary_1447_inst_ack_0 : boolean;
  signal type_cast_1464_inst_ack_0 : boolean;
  signal binary_1459_inst_ack_0 : boolean;
  signal binary_1486_inst_ack_0 : boolean;
  signal binary_1486_inst_ack_1 : boolean;
  signal binary_1474_inst_req_0 : boolean;
  signal type_cast_1522_inst_ack_0 : boolean;
  signal binary_1513_inst_req_0 : boolean;
  signal binary_1508_inst_req_1 : boolean;
  signal binary_1513_inst_req_1 : boolean;
  signal binary_1502_inst_req_1 : boolean;
  signal simple_obj_ref_1539_inst_ack_0 : boolean;
  signal binary_1459_inst_ack_1 : boolean;
  signal binary_1474_inst_ack_0 : boolean;
  signal binary_1437_inst_req_0 : boolean;
  signal type_cast_1441_inst_ack_0 : boolean;
  signal ternary_1492_inst_ack_0 : boolean;
  signal binary_1502_inst_ack_0 : boolean;
  signal binary_1437_inst_ack_0 : boolean;
  signal binary_1468_inst_req_0 : boolean;
  signal binary_1474_inst_ack_1 : boolean;
  signal binary_1502_inst_ack_1 : boolean;
  signal binary_1437_inst_req_1 : boolean;
  signal binary_1468_inst_ack_0 : boolean;
  signal binary_1437_inst_ack_1 : boolean;
  signal binary_1474_inst_req_1 : boolean;
  signal binary_1424_inst_req_0 : boolean;
  signal binary_1468_inst_req_1 : boolean;
  signal binary_1424_inst_ack_0 : boolean;
  signal binary_1453_inst_ack_1 : boolean;
  signal binary_1453_inst_req_1 : boolean;
  signal binary_1468_inst_ack_1 : boolean;
  signal binary_1453_inst_req_0 : boolean;
  signal binary_1424_inst_req_1 : boolean;
  signal binary_1424_inst_ack_1 : boolean;
  signal binary_1513_inst_ack_0 : boolean;
  signal simple_obj_ref_1530_inst_req_0 : boolean;
  signal binary_1508_inst_req_0 : boolean;
  signal binary_1453_inst_ack_0 : boolean;
  signal type_cast_1496_inst_req_0 : boolean;
  signal type_cast_1520_inst_ack_0 : boolean;
  signal phi_stmt_1517_ack_0 : boolean;
  signal binary_1480_inst_req_0 : boolean;
  signal simple_obj_ref_1530_inst_ack_0 : boolean;
  signal binary_1447_inst_req_1 : boolean;
  signal binary_1480_inst_ack_0 : boolean;
  signal if_stmt_1426_branch_req_0 : boolean;
  signal type_cast_1522_inst_req_0 : boolean;
  signal ternary_1492_inst_req_0 : boolean;
  signal if_stmt_1426_branch_ack_1 : boolean;
  signal type_cast_1496_inst_ack_0 : boolean;
  signal binary_1447_inst_ack_1 : boolean;
  signal binary_1508_inst_ack_1 : boolean;
  signal simple_obj_ref_1539_inst_req_0 : boolean;
  signal binary_1459_inst_req_0 : boolean;
  signal if_stmt_1426_branch_ack_0 : boolean;
  signal type_cast_1520_inst_req_0 : boolean;
  signal phi_stmt_1517_req_0 : boolean;
  signal binary_1486_inst_req_1 : boolean;
  signal phi_stmt_1517_req_1 : boolean;
  signal simple_obj_ref_1398_inst_ack_0 : boolean;
  signal simple_obj_ref_1398_inst_req_0 : boolean;
  signal binary_1480_inst_ack_1 : boolean;
  signal binary_1508_inst_ack_0 : boolean;
  signal binary_1513_inst_ack_1 : boolean;
  signal binary_1502_inst_req_0 : boolean;
  signal binary_1480_inst_req_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  output_port_lookup_CP_6603: Block -- control-path 
    signal cp_elements: BooleanArray(100 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    simple_obj_ref_1398_inst_req_0 <= cp_elements(0);
    cp_elements(1) <= false; 
    cp_elements(2) <= OrReduce(cp_elements(18) & cp_elements(89));
    cp_elements(3) <= simple_obj_ref_1398_inst_ack_0;
    cp_elements(4) <= simple_obj_ref_1409_inst_ack_0;
    simple_obj_ref_1418_inst_req_0 <= cp_elements(4);
    cp_elements(5) <= simple_obj_ref_1418_inst_ack_0;
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(8) & cp_elements(9));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1424_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= cp_elements(6);
    cp_elements(9) <= cp_elements(6);
    cp_elements(10) <= binary_1424_inst_ack_0;
    binary_1424_inst_req_1 <= cp_elements(10);
    cp_elements(11) <= binary_1424_inst_ack_1;
    cp_elements(12) <= cp_elements(11);
    cp_elements(13) <= false;
    cp_elements(14) <= cp_elements(13);
    cp_elements(15) <= cp_elements(11);
    if_stmt_1426_branch_req_0 <= cp_elements(15);
    cp_elements(16) <= cp_elements(15);
    cp_elements(17) <= cp_elements(16);
    cp_elements(18) <= if_stmt_1426_branch_ack_1;
    cp_elements(19) <= cp_elements(16);
    cp_elements(20) <= if_stmt_1426_branch_ack_0;
    cp_elements(21) <= cp_elements(2);
    cpelement_group_22 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(23) & cp_elements(24));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(22),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1437_inst_req_0 <= cp_elements(22);
    cp_elements(23) <= cp_elements(21);
    cp_elements(24) <= cp_elements(21);
    cp_elements(25) <= binary_1437_inst_ack_0;
    binary_1437_inst_req_1 <= cp_elements(25);
    cp_elements(26) <= binary_1437_inst_ack_1;
    cpelement_group_27 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(28) & cp_elements(29));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(27),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1441_inst_req_0 <= cp_elements(27);
    cp_elements(28) <= cp_elements(21);
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= type_cast_1441_inst_ack_0;
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(32));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1447_inst_req_0 <= cp_elements(31);
    cp_elements(32) <= cp_elements(21);
    cp_elements(33) <= binary_1447_inst_ack_0;
    binary_1447_inst_req_1 <= cp_elements(33);
    cp_elements(34) <= binary_1447_inst_ack_1;
    cpelement_group_35 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(34) & cp_elements(36));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(35),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1453_inst_req_0 <= cp_elements(35);
    cp_elements(36) <= cp_elements(21);
    cp_elements(37) <= binary_1453_inst_ack_0;
    binary_1453_inst_req_1 <= cp_elements(37);
    cp_elements(38) <= binary_1453_inst_ack_1;
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(40) & cp_elements(41));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1459_inst_req_0 <= cp_elements(39);
    cp_elements(40) <= cp_elements(21);
    cp_elements(41) <= cp_elements(26);
    cp_elements(42) <= binary_1459_inst_ack_0;
    binary_1459_inst_req_1 <= cp_elements(42);
    cp_elements(43) <= binary_1459_inst_ack_1;
    cpelement_group_44 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(48));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(44),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1468_inst_req_0 <= cp_elements(44);
    cp_elements(45) <= cp_elements(21);
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(43) & cp_elements(47));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1464_inst_req_0 <= cp_elements(46);
    cp_elements(47) <= cp_elements(21);
    cp_elements(48) <= type_cast_1464_inst_ack_0;
    cp_elements(49) <= binary_1468_inst_ack_0;
    binary_1468_inst_req_1 <= cp_elements(49);
    cp_elements(50) <= binary_1468_inst_ack_1;
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(52) & cp_elements(53));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1474_inst_req_0 <= cp_elements(51);
    cp_elements(52) <= cp_elements(21);
    cp_elements(53) <= cp_elements(38);
    cp_elements(54) <= binary_1474_inst_ack_0;
    binary_1474_inst_req_1 <= cp_elements(54);
    cp_elements(55) <= binary_1474_inst_ack_1;
    cpelement_group_56 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(55) & cp_elements(57));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(56),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1480_inst_req_0 <= cp_elements(56);
    cp_elements(57) <= cp_elements(21);
    cp_elements(58) <= binary_1480_inst_ack_0;
    binary_1480_inst_req_1 <= cp_elements(58);
    cp_elements(59) <= binary_1480_inst_ack_1;
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1486_inst_req_0 <= cp_elements(60);
    cp_elements(61) <= cp_elements(21);
    cp_elements(62) <= cp_elements(38);
    cp_elements(63) <= binary_1486_inst_ack_0;
    binary_1486_inst_req_1 <= cp_elements(63);
    cp_elements(64) <= binary_1486_inst_ack_1;
    cp_elements(65) <= cp_elements(21);
    cpelement_group_66 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(59) & cp_elements(64) & cp_elements(65));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(66),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ternary_1492_inst_req_0 <= cp_elements(66);
    cp_elements(67) <= ternary_1492_inst_ack_0;
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(67) & cp_elements(69));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1496_inst_req_0 <= cp_elements(68);
    cp_elements(69) <= cp_elements(21);
    cp_elements(70) <= type_cast_1496_inst_ack_0;
    cpelement_group_71 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(72) & cp_elements(73));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(71),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1502_inst_req_0 <= cp_elements(71);
    cp_elements(72) <= cp_elements(21);
    cp_elements(73) <= cp_elements(21);
    cp_elements(74) <= binary_1502_inst_ack_0;
    binary_1502_inst_req_1 <= cp_elements(74);
    cp_elements(75) <= binary_1502_inst_ack_1;
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(77));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1508_inst_req_0 <= cp_elements(76);
    cp_elements(77) <= cp_elements(21);
    cp_elements(78) <= binary_1508_inst_ack_0;
    binary_1508_inst_req_1 <= cp_elements(78);
    cp_elements(79) <= binary_1508_inst_ack_1;
    cpelement_group_80 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(79) & cp_elements(81));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(80),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1513_inst_req_0 <= cp_elements(80);
    cp_elements(81) <= cp_elements(21);
    cp_elements(82) <= binary_1513_inst_ack_0;
    binary_1513_inst_req_1 <= cp_elements(82);
    cp_elements(83) <= binary_1513_inst_ack_1;
    cp_elements(84) <= simple_obj_ref_1530_inst_ack_0;
    simple_obj_ref_1539_inst_req_0 <= cp_elements(84);
    cp_elements(85) <= simple_obj_ref_1539_inst_ack_0;
    cp_elements(86) <= OrReduce(cp_elements(3) & cp_elements(85));
    cp_elements(87) <= cp_elements(86);
    simple_obj_ref_1409_inst_req_0 <= cp_elements(87);
    cp_elements(88) <= false;
    cp_elements(89) <= cp_elements(88);
    cp_elements(90) <= cp_elements(20);
    cp_elements(91) <= cp_elements(20);
    type_cast_1522_inst_req_0 <= cp_elements(91);
    cp_elements(92) <= type_cast_1522_inst_ack_0;
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(90) & cp_elements(92));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1517_req_1 <= cp_elements(93);
    cp_elements(94) <= cp_elements(83);
    type_cast_1520_inst_req_0 <= cp_elements(94);
    cp_elements(95) <= type_cast_1520_inst_ack_0;
    cp_elements(96) <= cp_elements(83);
    cpelement_group_97 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(95) & cp_elements(96));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(97),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1517_req_0 <= cp_elements(97);
    cp_elements(98) <= OrReduce(cp_elements(93) & cp_elements(97));
    cp_elements(99) <= cp_elements(98);
    cp_elements(100) <= phi_stmt_1517_ack_0;
    simple_obj_ref_1530_inst_req_0 <= cp_elements(100);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal datax_x0_1517 : std_logic_vector(63 downto 0);
    signal iNsTr_0_1396 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1407 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1416 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1529 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1538 : std_logic_vector(31 downto 0);
    signal tmp10_1460 : std_logic_vector(63 downto 0);
    signal tmp11_1469 : std_logic_vector(0 downto 0);
    signal tmp12_1475 : std_logic_vector(31 downto 0);
    signal tmp13_1481 : std_logic_vector(31 downto 0);
    signal tmp14_1487 : std_logic_vector(31 downto 0);
    signal tmp15_1493 : std_logic_vector(31 downto 0);
    signal tmp16_1497 : std_logic_vector(63 downto 0);
    signal tmp17_1503 : std_logic_vector(63 downto 0);
    signal tmp18_1509 : std_logic_vector(63 downto 0);
    signal tmp19_1514 : std_logic_vector(63 downto 0);
    signal tmp1_1399 : std_logic_vector(7 downto 0);
    signal tmp3_1410 : std_logic_vector(7 downto 0);
    signal tmp4_1419 : std_logic_vector(63 downto 0);
    signal tmp5_1425 : std_logic_vector(0 downto 0);
    signal tmp7_1438 : std_logic_vector(63 downto 0);
    signal tmp8_1448 : std_logic_vector(31 downto 0);
    signal tmp9_1454 : std_logic_vector(31 downto 0);
    signal tmp_1442 : std_logic_vector(31 downto 0);
    signal type_cast_1423_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1451_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1458_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1464_wire : std_logic_vector(63 downto 0);
    signal type_cast_1467_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1473_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1479_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1485_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1507_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1520_wire : std_logic_vector(63 downto 0);
    signal type_cast_1522_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    iNsTr_0_1396 <= "00000000000000000000000000000000";
    iNsTr_2_1407 <= "00000000000000000000000000000000";
    iNsTr_3_1416 <= "00000000000000000000000000000000";
    iNsTr_6_1529 <= "00000000000000000000000000000000";
    iNsTr_8_1538 <= "00000000000000000000000000000000";
    type_cast_1423_wire_constant <= "11111111";
    type_cast_1436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1446_wire_constant <= "00000000000000001111111111111111";
    type_cast_1451_wire_constant <= "00000000000000000000000000000001";
    type_cast_1458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1467_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1473_wire_constant <= "00000000000000000000000000000001";
    type_cast_1479_wire_constant <= "00000000000000000111111111111111";
    type_cast_1485_wire_constant <= "00000000000000000000000000000001";
    type_cast_1501_wire_constant <= "0000000000000000111111111111111111111111111111111111111111111111";
    type_cast_1507_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    phi_stmt_1517: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1520_wire & type_cast_1522_wire;
      req <= phi_stmt_1517_req_0 & phi_stmt_1517_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1517_ack_0,
          idata => idata,
          odata => datax_x0_1517,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1517
    ternary_1492_inst: SelectBase generic map(data_width => 32) -- 
      port map( x => tmp13_1481, y => tmp14_1487, sel => tmp11_1469, z => tmp15_1493, req => ternary_1492_inst_req_0, ack => ternary_1492_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1441_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_1438, dout => tmp_1442, req => type_cast_1441_inst_req_0, ack => type_cast_1441_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1464_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 64, flow_through => true ) 
      port map( din => tmp10_1460, dout => type_cast_1464_wire, req => type_cast_1464_inst_req_0, ack => type_cast_1464_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1496_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 64, flow_through => false ) 
      port map( din => tmp15_1493, dout => tmp16_1497, req => type_cast_1496_inst_req_0, ack => type_cast_1496_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1520_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 64, flow_through => true ) 
      port map( din => tmp19_1514, dout => type_cast_1520_wire, req => type_cast_1520_inst_req_0, ack => type_cast_1520_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1522_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 64, flow_through => true ) 
      port map( din => tmp4_1419, dout => type_cast_1522_wire, req => type_cast_1522_inst_req_0, ack => type_cast_1522_inst_ack_0, clk => clk, reset => reset); -- 
    if_stmt_1426_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp5_1425;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1426_branch_req_0,
          ack0 => if_stmt_1426_branch_ack_0,
          ack1 => if_stmt_1426_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_1424_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp3_1410;
      tmp5_1425 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1424_inst_req_0,
          ackL => binary_1424_inst_ack_0,
          reqR => binary_1424_inst_req_1,
          ackR => binary_1424_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_1437_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp4_1419;
      tmp7_1438 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1437_inst_req_0,
          ackL => binary_1437_inst_ack_0,
          reqR => binary_1437_inst_req_1,
          ackR => binary_1437_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1447_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1442;
      tmp8_1448 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1447_inst_req_0,
          ackL => binary_1447_inst_ack_0,
          reqR => binary_1447_inst_req_1,
          ackR => binary_1447_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1453_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1451_wire_constant & tmp8_1448;
      tmp9_1454 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1453_inst_req_0,
          ackL => binary_1453_inst_ack_0,
          reqR => binary_1453_inst_req_1,
          ackR => binary_1453_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_1459_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp7_1438;
      tmp10_1460 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1459_inst_req_0,
          ackL => binary_1459_inst_ack_0,
          reqR => binary_1459_inst_req_1,
          ackR => binary_1459_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_1468_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1464_wire;
      tmp11_1469 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1468_inst_req_0,
          ackL => binary_1468_inst_ack_0,
          reqR => binary_1468_inst_req_1,
          ackR => binary_1468_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_1474_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp9_1454;
      tmp12_1475 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1474_inst_req_0,
          ackL => binary_1474_inst_ack_0,
          reqR => binary_1474_inst_req_1,
          ackR => binary_1474_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_1480_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp12_1475;
      tmp13_1481 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1480_inst_req_0,
          ackL => binary_1480_inst_ack_0,
          reqR => binary_1480_inst_req_1,
          ackR => binary_1480_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_1486_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp9_1454;
      tmp14_1487 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1486_inst_req_0,
          ackL => binary_1486_inst_ack_0,
          reqR => binary_1486_inst_req_1,
          ackR => binary_1486_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_1502_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp4_1419;
      tmp17_1503 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000111111111111111111111111111111111111111111111111",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1502_inst_req_0,
          ackL => binary_1502_inst_ack_0,
          reqR => binary_1502_inst_req_1,
          ackR => binary_1502_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_1508_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp16_1497;
      tmp18_1509 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1508_inst_req_0,
          ackL => binary_1508_inst_ack_0,
          reqR => binary_1508_inst_req_1,
          ackR => binary_1508_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_1513_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_1509 & tmp17_1503;
      tmp19_1514 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1513_inst_req_0,
          ackL => binary_1513_inst_ack_0,
          reqR => binary_1513_inst_req_1,
          ackR => binary_1513_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared inport operator group (0) : simple_obj_ref_1398_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1398_inst_req_0;
      simple_obj_ref_1398_inst_ack_0 <= ack(0);
      tmp1_1399 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => start_output_port_lookup_pipe_read_req(0),
          oack => start_output_port_lookup_pipe_read_ack(0),
          odata => start_output_port_lookup_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1409_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1409_inst_req_0;
      simple_obj_ref_1409_inst_ack_0 <= ack(0);
      tmp3_1410 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => op_lut_ctrl_pipe_read_req(0),
          oack => op_lut_ctrl_pipe_read_ack(0),
          odata => op_lut_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_1418_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1418_inst_req_0;
      simple_obj_ref_1418_inst_ack_0 <= ack(0);
      tmp4_1419 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => op_lut_data_pipe_read_req(0),
          oack => op_lut_data_pipe_read_ack(0),
          odata => op_lut_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : simple_obj_ref_1530_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1530_inst_req_0;
      simple_obj_ref_1530_inst_ack_0 <= ack(0);
      data_in <= tmp3_1410;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_ctrl_pipe_write_req(0),
          oack => out_ctrl_pipe_write_ack(0),
          odata => out_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_1539_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1539_inst_req_0;
      simple_obj_ref_1539_inst_ack_0 <= ack(0);
      data_in <= datax_x0_1517;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_input is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(87 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(15 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(7 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(15 downto 0);
    free_queue_ack_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
    in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    start_wrapper_input_pipe_read_req : out  std_logic_vector(0 downto 0);
    start_wrapper_input_pipe_read_ack : in   std_logic_vector(0 downto 0);
    start_wrapper_input_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    midpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    midpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    midpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    last_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    last_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    last_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    pkt_length_pipe_write_req : out  std_logic_vector(0 downto 0);
    pkt_length_pipe_write_ack : in   std_logic_vector(0 downto 0);
    pkt_length_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_input;
architecture Default of wrapper_input is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_input_CP_6993_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_1719_base_resize_req_0 : boolean;
  signal ptr_deref_1747_base_resize_ack_0 : boolean;
  signal binary_1740_inst_ack_0 : boolean;
  signal type_cast_1744_inst_req_0 : boolean;
  signal array_obj_ref_1657_root_address_inst_req_0 : boolean;
  signal ptr_deref_1747_store_0_ack_0 : boolean;
  signal ptr_deref_1719_base_resize_ack_0 : boolean;
  signal ptr_deref_1747_gather_scatter_req_0 : boolean;
  signal ptr_deref_1719_addr_0_req_0 : boolean;
  signal ptr_deref_1733_root_address_inst_req_0 : boolean;
  signal ptr_deref_1747_store_0_ack_1 : boolean;
  signal array_obj_ref_1884_base_resize_ack_0 : boolean;
  signal binary_1740_inst_req_0 : boolean;
  signal binary_1740_inst_ack_1 : boolean;
  signal array_obj_ref_1657_final_reg_req_0 : boolean;
  signal array_obj_ref_1652_root_address_inst_ack_0 : boolean;
  signal binary_1673_inst_ack_1 : boolean;
  signal binary_1712_inst_req_1 : boolean;
  signal type_cast_1744_inst_ack_0 : boolean;
  signal array_obj_ref_1647_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1647_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1876_final_reg_req_0 : boolean;
  signal ptr_deref_2093_addr_0_ack_0 : boolean;
  signal ptr_deref_1761_addr_0_ack_0 : boolean;
  signal ptr_deref_1747_addr_0_req_0 : boolean;
  signal ptr_deref_1733_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1884_index_0_resize_ack_0 : boolean;
  signal binary_1712_inst_ack_1 : boolean;
  signal array_obj_ref_1647_root_address_inst_req_1 : boolean;
  signal ptr_deref_1747_base_resize_req_0 : boolean;
  signal array_obj_ref_1647_final_reg_ack_0 : boolean;
  signal type_cast_1716_inst_req_0 : boolean;
  signal array_obj_ref_1652_root_address_inst_req_1 : boolean;
  signal type_cast_1695_inst_ack_0 : boolean;
  signal switch_stmt_1697_branch_default_req_0 : boolean;
  signal array_obj_ref_1657_base_resize_ack_0 : boolean;
  signal type_cast_1695_inst_req_0 : boolean;
  signal switch_stmt_1697_branch_default_ack_0 : boolean;
  signal type_cast_1730_inst_ack_0 : boolean;
  signal simple_obj_ref_1682_inst_req_0 : boolean;
  signal ptr_deref_1733_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1901_base_resize_ack_0 : boolean;
  signal ptr_deref_1747_store_0_req_0 : boolean;
  signal switch_stmt_1697_branch_1_ack_1 : boolean;
  signal binary_1754_inst_req_1 : boolean;
  signal ptr_deref_1915_root_address_inst_req_0 : boolean;
  signal binary_1726_inst_req_0 : boolean;
  signal ptr_deref_1719_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1719_store_0_ack_0 : boolean;
  signal simple_obj_ref_1691_inst_req_0 : boolean;
  signal ptr_deref_1901_gather_scatter_ack_0 : boolean;
  signal type_cast_1730_inst_req_0 : boolean;
  signal ptr_deref_1733_store_0_ack_0 : boolean;
  signal binary_1673_inst_ack_0 : boolean;
  signal type_cast_1716_inst_ack_0 : boolean;
  signal type_cast_1758_inst_req_0 : boolean;
  signal binary_1754_inst_ack_1 : boolean;
  signal array_obj_ref_1647_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1657_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1647_final_reg_req_0 : boolean;
  signal ptr_deref_1719_addr_0_ack_0 : boolean;
  signal array_obj_ref_2042_index_0_resize_ack_0 : boolean;
  signal phi_stmt_1661_req_0 : boolean;
  signal array_obj_ref_1864_index_0_rename_req_0 : boolean;
  signal binary_1726_inst_ack_1 : boolean;
  signal binary_1712_inst_ack_0 : boolean;
  signal ptr_deref_1747_store_0_req_1 : boolean;
  signal binary_1712_inst_req_0 : boolean;
  signal ptr_deref_1719_store_0_req_0 : boolean;
  signal ptr_deref_1733_base_resize_ack_0 : boolean;
  signal ptr_deref_1733_base_resize_req_0 : boolean;
  signal binary_1726_inst_ack_0 : boolean;
  signal array_obj_ref_1647_base_resize_req_0 : boolean;
  signal binary_1740_inst_req_1 : boolean;
  signal ptr_deref_1733_store_0_req_0 : boolean;
  signal array_obj_ref_1657_base_resize_req_0 : boolean;
  signal array_obj_ref_1864_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1652_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_1682_inst_ack_0 : boolean;
  signal array_obj_ref_1647_base_resize_ack_0 : boolean;
  signal simple_obj_ref_1691_inst_ack_0 : boolean;
  signal binary_1726_inst_req_1 : boolean;
  signal array_obj_ref_1652_base_resize_req_0 : boolean;
  signal array_obj_ref_2042_offset_inst_req_0 : boolean;
  signal binary_1673_inst_req_0 : boolean;
  signal ptr_deref_2093_addr_0_req_0 : boolean;
  signal ptr_deref_1761_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1652_final_reg_req_0 : boolean;
  signal ptr_deref_1719_store_0_req_1 : boolean;
  signal ptr_deref_1719_store_0_ack_1 : boolean;
  signal ptr_deref_1761_base_resize_req_0 : boolean;
  signal array_obj_ref_1864_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2069_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1761_store_0_ack_0 : boolean;
  signal ptr_deref_1761_gather_scatter_req_0 : boolean;
  signal ptr_deref_1761_store_0_req_0 : boolean;
  signal binary_1754_inst_ack_0 : boolean;
  signal array_obj_ref_1652_final_reg_ack_0 : boolean;
  signal array_obj_ref_2042_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1868_final_reg_req_0 : boolean;
  signal ptr_deref_1761_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1872_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1901_store_0_ack_0 : boolean;
  signal type_cast_1758_inst_ack_0 : boolean;
  signal array_obj_ref_1876_final_reg_ack_0 : boolean;
  signal ptr_deref_1761_addr_0_req_0 : boolean;
  signal type_cast_1912_inst_ack_0 : boolean;
  signal ptr_deref_1761_base_resize_ack_0 : boolean;
  signal ptr_deref_1719_gather_scatter_req_0 : boolean;
  signal ptr_deref_1747_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1719_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1652_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1868_final_reg_ack_0 : boolean;
  signal ptr_deref_2093_base_resize_ack_0 : boolean;
  signal ptr_deref_1733_addr_0_req_0 : boolean;
  signal binary_1673_inst_req_1 : boolean;
  signal ptr_deref_1719_root_address_inst_req_0 : boolean;
  signal switch_stmt_1697_select_expr_0_req_1 : boolean;
  signal ptr_deref_1733_store_0_req_1 : boolean;
  signal array_obj_ref_1657_root_address_inst_req_1 : boolean;
  signal ptr_deref_1733_addr_0_ack_0 : boolean;
  signal array_obj_ref_1657_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1733_store_0_ack_1 : boolean;
  signal ptr_deref_1915_base_resize_req_0 : boolean;
  signal array_obj_ref_1652_base_resize_ack_0 : boolean;
  signal ptr_deref_1747_root_address_inst_req_0 : boolean;
  signal ptr_deref_1761_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1657_final_reg_ack_0 : boolean;
  signal switch_stmt_1697_select_expr_0_req_0 : boolean;
  signal ptr_deref_1733_gather_scatter_req_0 : boolean;
  signal binary_1754_inst_req_0 : boolean;
  signal ptr_deref_1747_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2090_final_reg_req_0 : boolean;
  signal array_obj_ref_1884_base_resize_req_0 : boolean;
  signal ptr_deref_1915_addr_0_ack_0 : boolean;
  signal ptr_deref_1747_addr_0_ack_0 : boolean;
  signal switch_stmt_1697_select_expr_0_ack_0 : boolean;
  signal switch_stmt_1697_branch_0_ack_1 : boolean;
  signal switch_stmt_1697_branch_1_req_0 : boolean;
  signal switch_stmt_1697_select_expr_1_ack_1 : boolean;
  signal switch_stmt_1697_select_expr_1_req_1 : boolean;
  signal binary_2100_inst_req_1 : boolean;
  signal switch_stmt_1697_select_expr_1_ack_0 : boolean;
  signal ptr_deref_2093_root_address_inst_req_0 : boolean;
  signal switch_stmt_1697_select_expr_1_req_0 : boolean;
  signal switch_stmt_1697_branch_0_req_0 : boolean;
  signal switch_stmt_1697_select_expr_0_ack_1 : boolean;
  signal array_obj_ref_1884_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1880_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1880_index_0_resize_ack_0 : boolean;
  signal binary_1922_inst_req_0 : boolean;
  signal array_obj_ref_1864_offset_inst_req_0 : boolean;
  signal array_obj_ref_1864_offset_inst_ack_0 : boolean;
  signal ptr_deref_1915_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1901_gather_scatter_req_0 : boolean;
  signal ptr_deref_1929_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2090_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1929_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2045_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1884_index_0_rename_req_0 : boolean;
  signal ptr_deref_1915_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1884_index_0_rename_ack_0 : boolean;
  signal ptr_deref_2093_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1864_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2066_base_resize_req_0 : boolean;
  signal ptr_deref_1915_base_resize_ack_0 : boolean;
  signal array_obj_ref_1884_offset_inst_req_0 : boolean;
  signal array_obj_ref_1880_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1864_base_resize_req_0 : boolean;
  signal array_obj_ref_1864_base_resize_ack_0 : boolean;
  signal array_obj_ref_1884_offset_inst_ack_0 : boolean;
  signal ptr_deref_1929_root_address_inst_req_0 : boolean;
  signal ptr_deref_1929_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2114_offset_inst_req_0 : boolean;
  signal ptr_deref_2045_gather_scatter_req_0 : boolean;
  signal ptr_deref_2069_root_address_inst_req_0 : boolean;
  signal ptr_deref_2069_base_resize_req_0 : boolean;
  signal ptr_deref_1915_addr_0_req_0 : boolean;
  signal array_obj_ref_1872_index_0_resize_req_0 : boolean;
  signal ptr_deref_1915_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1880_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1864_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1880_offset_inst_req_0 : boolean;
  signal array_obj_ref_1864_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2066_final_reg_req_0 : boolean;
  signal binary_1922_inst_req_1 : boolean;
  signal array_obj_ref_1880_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1864_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1872_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1880_base_resize_req_0 : boolean;
  signal array_obj_ref_1880_base_resize_ack_0 : boolean;
  signal binary_1922_inst_ack_1 : boolean;
  signal ptr_deref_1901_base_resize_req_0 : boolean;
  signal array_obj_ref_1872_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1880_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1880_root_address_inst_ack_0 : boolean;
  signal binary_1922_inst_ack_0 : boolean;
  signal array_obj_ref_2066_final_reg_ack_0 : boolean;
  signal array_obj_ref_1864_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1880_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1880_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1880_final_reg_req_0 : boolean;
  signal ptr_deref_2093_base_resize_req_0 : boolean;
  signal array_obj_ref_1864_final_reg_req_0 : boolean;
  signal array_obj_ref_2042_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1880_final_reg_ack_0 : boolean;
  signal ptr_deref_1554_gather_scatter_req_0 : boolean;
  signal ptr_deref_1554_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1554_store_0_req_0 : boolean;
  signal ptr_deref_1554_store_0_ack_0 : boolean;
  signal ptr_deref_1554_store_0_req_1 : boolean;
  signal ptr_deref_1554_store_0_ack_1 : boolean;
  signal type_cast_1912_inst_req_0 : boolean;
  signal ptr_deref_2045_store_0_ack_1 : boolean;
  signal array_obj_ref_1864_final_reg_ack_0 : boolean;
  signal simple_obj_ref_1565_inst_req_0 : boolean;
  signal simple_obj_ref_1565_inst_ack_0 : boolean;
  signal ptr_deref_2069_base_resize_ack_0 : boolean;
  signal simple_obj_ref_1575_inst_req_0 : boolean;
  signal simple_obj_ref_1575_inst_ack_0 : boolean;
  signal simple_obj_ref_1586_inst_req_0 : boolean;
  signal simple_obj_ref_1586_inst_ack_0 : boolean;
  signal binary_1592_inst_req_0 : boolean;
  signal binary_1592_inst_ack_0 : boolean;
  signal binary_1592_inst_req_1 : boolean;
  signal binary_1592_inst_ack_1 : boolean;
  signal if_stmt_1594_branch_req_0 : boolean;
  signal if_stmt_1594_branch_ack_1 : boolean;
  signal if_stmt_1594_branch_ack_0 : boolean;
  signal simple_obj_ref_1608_inst_req_0 : boolean;
  signal simple_obj_ref_1608_inst_ack_0 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal type_cast_1618_inst_req_0 : boolean;
  signal type_cast_1618_inst_ack_0 : boolean;
  signal array_obj_ref_1884_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1623_base_resize_req_0 : boolean;
  signal array_obj_ref_1623_base_resize_ack_0 : boolean;
  signal array_obj_ref_1623_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1623_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1623_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1623_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1623_final_reg_req_0 : boolean;
  signal array_obj_ref_1623_final_reg_ack_0 : boolean;
  signal array_obj_ref_1628_base_resize_req_0 : boolean;
  signal array_obj_ref_1628_base_resize_ack_0 : boolean;
  signal array_obj_ref_1628_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1628_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1628_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1628_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1628_final_reg_req_0 : boolean;
  signal array_obj_ref_1628_final_reg_ack_0 : boolean;
  signal array_obj_ref_1633_base_resize_req_0 : boolean;
  signal array_obj_ref_1633_base_resize_ack_0 : boolean;
  signal array_obj_ref_1633_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1633_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1633_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1633_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1633_final_reg_req_0 : boolean;
  signal array_obj_ref_1633_final_reg_ack_0 : boolean;
  signal array_obj_ref_1638_base_resize_req_0 : boolean;
  signal array_obj_ref_1638_base_resize_ack_0 : boolean;
  signal array_obj_ref_1638_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1638_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1638_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1638_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1638_final_reg_req_0 : boolean;
  signal array_obj_ref_1638_final_reg_ack_0 : boolean;
  signal type_cast_1642_inst_req_0 : boolean;
  signal type_cast_1642_inst_ack_0 : boolean;
  signal array_obj_ref_1876_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1761_store_0_req_1 : boolean;
  signal array_obj_ref_1876_root_address_inst_req_1 : boolean;
  signal ptr_deref_1761_store_0_ack_1 : boolean;
  signal array_obj_ref_2066_base_resize_ack_0 : boolean;
  signal ptr_deref_1929_addr_0_ack_0 : boolean;
  signal array_obj_ref_2066_root_address_inst_req_1 : boolean;
  signal binary_2062_inst_req_0 : boolean;
  signal ptr_deref_2045_store_0_req_0 : boolean;
  signal array_obj_ref_1876_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1876_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2114_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_ack_1 : boolean;
  signal binary_1768_inst_req_0 : boolean;
  signal type_cast_1898_inst_ack_0 : boolean;
  signal binary_1768_inst_ack_0 : boolean;
  signal type_cast_1898_inst_req_0 : boolean;
  signal binary_1768_inst_req_1 : boolean;
  signal binary_1768_inst_ack_1 : boolean;
  signal ptr_deref_1929_addr_0_req_0 : boolean;
  signal ptr_deref_1901_store_0_req_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1876_base_resize_ack_0 : boolean;
  signal array_obj_ref_1876_base_resize_req_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2114_index_0_rename_req_0 : boolean;
  signal ptr_deref_1901_addr_0_ack_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_req_0 : boolean;
  signal type_cast_1772_inst_req_0 : boolean;
  signal type_cast_1772_inst_ack_0 : boolean;
  signal array_obj_ref_1876_offset_inst_ack_0 : boolean;
  signal binary_1908_inst_ack_1 : boolean;
  signal ptr_deref_2069_addr_0_req_0 : boolean;
  signal ptr_deref_1901_addr_0_req_0 : boolean;
  signal binary_1894_inst_ack_1 : boolean;
  signal array_obj_ref_1876_offset_inst_req_0 : boolean;
  signal binary_1894_inst_req_1 : boolean;
  signal binary_1894_inst_ack_0 : boolean;
  signal binary_1894_inst_req_0 : boolean;
  signal array_obj_ref_1876_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1876_index_0_rename_req_0 : boolean;
  signal ptr_deref_1775_base_resize_req_0 : boolean;
  signal ptr_deref_1775_base_resize_ack_0 : boolean;
  signal ptr_deref_2117_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2069_addr_0_ack_0 : boolean;
  signal ptr_deref_1775_root_address_inst_req_0 : boolean;
  signal ptr_deref_1775_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1868_base_resize_ack_0 : boolean;
  signal ptr_deref_1775_addr_0_req_0 : boolean;
  signal ptr_deref_1775_addr_0_ack_0 : boolean;
  signal array_obj_ref_2042_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1868_base_resize_req_0 : boolean;
  signal array_obj_ref_1888_final_reg_ack_0 : boolean;
  signal ptr_deref_1775_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1888_final_reg_req_0 : boolean;
  signal ptr_deref_1775_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1915_store_0_ack_1 : boolean;
  signal ptr_deref_1775_store_0_req_0 : boolean;
  signal array_obj_ref_1876_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1775_store_0_ack_0 : boolean;
  signal ptr_deref_1915_store_0_req_1 : boolean;
  signal ptr_deref_1775_store_0_req_1 : boolean;
  signal array_obj_ref_1876_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1888_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1775_store_0_ack_1 : boolean;
  signal array_obj_ref_2066_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2090_final_reg_ack_0 : boolean;
  signal array_obj_ref_2066_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2066_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1888_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1888_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1888_root_address_inst_req_0 : boolean;
  signal ptr_deref_1901_store_0_ack_1 : boolean;
  signal binary_1908_inst_req_1 : boolean;
  signal binary_1782_inst_req_0 : boolean;
  signal binary_1782_inst_ack_0 : boolean;
  signal binary_1782_inst_req_1 : boolean;
  signal binary_1782_inst_ack_1 : boolean;
  signal simple_obj_ref_2216_inst_req_0 : boolean;
  signal array_obj_ref_1868_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1888_base_resize_ack_0 : boolean;
  signal array_obj_ref_1888_base_resize_req_0 : boolean;
  signal type_cast_1926_inst_ack_0 : boolean;
  signal array_obj_ref_1868_offset_inst_req_0 : boolean;
  signal type_cast_1786_inst_req_0 : boolean;
  signal type_cast_1786_inst_ack_0 : boolean;
  signal ptr_deref_1929_base_resize_ack_0 : boolean;
  signal array_obj_ref_1888_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2042_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2114_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1868_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1888_offset_inst_req_0 : boolean;
  signal array_obj_ref_1872_final_reg_ack_0 : boolean;
  signal array_obj_ref_1872_final_reg_req_0 : boolean;
  signal array_obj_ref_1888_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1888_index_0_rename_req_0 : boolean;
  signal ptr_deref_1789_base_resize_req_0 : boolean;
  signal ptr_deref_1789_base_resize_ack_0 : boolean;
  signal array_obj_ref_2114_root_address_inst_req_1 : boolean;
  signal ptr_deref_1901_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2045_store_0_req_1 : boolean;
  signal array_obj_ref_1868_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1888_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1789_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1888_index_0_resize_req_0 : boolean;
  signal ptr_deref_1789_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1901_root_address_inst_req_0 : boolean;
  signal ptr_deref_1789_addr_0_req_0 : boolean;
  signal ptr_deref_1789_addr_0_ack_0 : boolean;
  signal binary_1908_inst_ack_0 : boolean;
  signal ptr_deref_1789_gather_scatter_req_0 : boolean;
  signal ptr_deref_1789_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1872_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1789_store_0_req_0 : boolean;
  signal array_obj_ref_1872_root_address_inst_req_1 : boolean;
  signal ptr_deref_1789_store_0_ack_0 : boolean;
  signal ptr_deref_1915_store_0_ack_0 : boolean;
  signal ptr_deref_1789_store_0_req_1 : boolean;
  signal array_obj_ref_1872_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1789_store_0_ack_1 : boolean;
  signal array_obj_ref_2114_base_resize_req_0 : boolean;
  signal array_obj_ref_1868_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1872_root_address_inst_req_0 : boolean;
  signal type_cast_1926_inst_req_0 : boolean;
  signal array_obj_ref_1868_index_0_resize_req_0 : boolean;
  signal ptr_deref_1901_store_0_req_1 : boolean;
  signal binary_1908_inst_req_0 : boolean;
  signal ptr_deref_1915_store_0_req_0 : boolean;
  signal binary_1796_inst_req_0 : boolean;
  signal binary_1796_inst_ack_0 : boolean;
  signal binary_1796_inst_req_1 : boolean;
  signal array_obj_ref_1884_final_reg_ack_0 : boolean;
  signal binary_1796_inst_ack_1 : boolean;
  signal ptr_deref_2045_store_0_ack_0 : boolean;
  signal array_obj_ref_1884_final_reg_req_0 : boolean;
  signal array_obj_ref_1872_base_resize_ack_0 : boolean;
  signal array_obj_ref_1872_base_resize_req_0 : boolean;
  signal array_obj_ref_2114_root_address_inst_ack_0 : boolean;
  signal type_cast_1800_inst_req_0 : boolean;
  signal array_obj_ref_1884_root_address_inst_ack_1 : boolean;
  signal type_cast_1800_inst_ack_0 : boolean;
  signal ptr_deref_1929_base_resize_req_0 : boolean;
  signal array_obj_ref_1884_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1884_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1872_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1872_offset_inst_req_0 : boolean;
  signal ptr_deref_1803_base_resize_req_0 : boolean;
  signal binary_2100_inst_ack_0 : boolean;
  signal ptr_deref_1803_base_resize_ack_0 : boolean;
  signal ptr_deref_1803_root_address_inst_req_0 : boolean;
  signal ptr_deref_1803_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1803_addr_0_req_0 : boolean;
  signal ptr_deref_1803_addr_0_ack_0 : boolean;
  signal binary_2052_inst_req_0 : boolean;
  signal binary_2052_inst_ack_0 : boolean;
  signal ptr_deref_1803_gather_scatter_req_0 : boolean;
  signal ptr_deref_1803_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1803_store_0_req_0 : boolean;
  signal ptr_deref_2069_gather_scatter_req_0 : boolean;
  signal ptr_deref_1803_store_0_ack_0 : boolean;
  signal ptr_deref_2093_gather_scatter_req_0 : boolean;
  signal ptr_deref_2069_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2093_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1803_store_0_req_1 : boolean;
  signal ptr_deref_1803_store_0_ack_1 : boolean;
  signal array_obj_ref_2042_base_resize_req_0 : boolean;
  signal binary_2100_inst_ack_1 : boolean;
  signal binary_2052_inst_req_1 : boolean;
  signal binary_2052_inst_ack_1 : boolean;
  signal array_obj_ref_2042_base_resize_ack_0 : boolean;
  signal ptr_deref_2069_store_0_req_0 : boolean;
  signal type_cast_1808_inst_req_0 : boolean;
  signal type_cast_1808_inst_ack_0 : boolean;
  signal ptr_deref_2069_store_0_ack_0 : boolean;
  signal ptr_deref_2093_store_0_req_0 : boolean;
  signal ptr_deref_2093_store_0_ack_0 : boolean;
  signal array_obj_ref_2042_root_address_inst_req_0 : boolean;
  signal ptr_deref_1811_base_resize_req_0 : boolean;
  signal ptr_deref_1811_base_resize_ack_0 : boolean;
  signal type_cast_2080_inst_req_0 : boolean;
  signal ptr_deref_2069_store_0_req_1 : boolean;
  signal ptr_deref_1811_root_address_inst_req_0 : boolean;
  signal ptr_deref_1811_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2042_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2114_base_resize_ack_0 : boolean;
  signal array_obj_ref_2042_root_address_inst_req_1 : boolean;
  signal ptr_deref_1811_addr_0_req_0 : boolean;
  signal type_cast_2080_inst_ack_0 : boolean;
  signal ptr_deref_1811_addr_0_ack_0 : boolean;
  signal array_obj_ref_2042_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1811_gather_scatter_req_0 : boolean;
  signal ptr_deref_1811_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2069_store_0_ack_1 : boolean;
  signal ptr_deref_1811_store_0_req_0 : boolean;
  signal ptr_deref_1811_store_0_ack_0 : boolean;
  signal array_obj_ref_2114_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1811_store_0_req_1 : boolean;
  signal ptr_deref_1811_store_0_ack_1 : boolean;
  signal array_obj_ref_2042_final_reg_req_0 : boolean;
  signal simple_obj_ref_2216_inst_ack_0 : boolean;
  signal array_obj_ref_2114_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2042_final_reg_ack_0 : boolean;
  signal ptr_deref_2093_store_0_req_1 : boolean;
  signal type_cast_2056_inst_req_0 : boolean;
  signal type_cast_2056_inst_ack_0 : boolean;
  signal binary_1820_inst_req_0 : boolean;
  signal ptr_deref_2093_store_0_ack_1 : boolean;
  signal binary_1820_inst_ack_0 : boolean;
  signal binary_1820_inst_req_1 : boolean;
  signal binary_1820_inst_ack_1 : boolean;
  signal binary_2076_inst_req_0 : boolean;
  signal ptr_deref_2117_base_resize_req_0 : boolean;
  signal binary_2076_inst_ack_0 : boolean;
  signal binary_1826_inst_req_0 : boolean;
  signal binary_1826_inst_ack_0 : boolean;
  signal binary_1826_inst_req_1 : boolean;
  signal binary_1826_inst_ack_1 : boolean;
  signal binary_2076_inst_req_1 : boolean;
  signal binary_2076_inst_ack_1 : boolean;
  signal binary_1832_inst_req_0 : boolean;
  signal binary_1832_inst_ack_0 : boolean;
  signal binary_2100_inst_req_0 : boolean;
  signal binary_1832_inst_req_1 : boolean;
  signal binary_1832_inst_ack_1 : boolean;
  signal binary_1838_inst_req_0 : boolean;
  signal binary_1838_inst_ack_0 : boolean;
  signal binary_1838_inst_req_1 : boolean;
  signal binary_1838_inst_ack_1 : boolean;
  signal binary_1844_inst_req_0 : boolean;
  signal binary_1844_inst_ack_0 : boolean;
  signal binary_1844_inst_req_1 : boolean;
  signal binary_1844_inst_ack_1 : boolean;
  signal binary_1850_inst_req_0 : boolean;
  signal binary_1850_inst_ack_0 : boolean;
  signal binary_1850_inst_req_1 : boolean;
  signal binary_1850_inst_ack_1 : boolean;
  signal binary_1856_inst_req_0 : boolean;
  signal binary_1856_inst_ack_0 : boolean;
  signal binary_1856_inst_req_1 : boolean;
  signal binary_1856_inst_ack_1 : boolean;
  signal array_obj_ref_1860_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1860_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1860_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1860_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1860_offset_inst_req_0 : boolean;
  signal array_obj_ref_1860_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1860_base_resize_req_0 : boolean;
  signal array_obj_ref_1860_base_resize_ack_0 : boolean;
  signal array_obj_ref_1860_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1860_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1860_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1860_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1860_final_reg_req_0 : boolean;
  signal array_obj_ref_1860_final_reg_ack_0 : boolean;
  signal array_obj_ref_2090_root_address_inst_req_1 : boolean;
  signal ptr_deref_1929_store_0_req_0 : boolean;
  signal array_obj_ref_2090_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1929_store_0_ack_0 : boolean;
  signal array_obj_ref_2090_root_address_inst_req_0 : boolean;
  signal ptr_deref_1929_store_0_req_1 : boolean;
  signal ptr_deref_1929_store_0_ack_1 : boolean;
  signal ptr_deref_2117_root_address_inst_req_0 : boolean;
  signal ptr_deref_2117_base_resize_ack_0 : boolean;
  signal type_cast_2104_inst_ack_0 : boolean;
  signal ptr_deref_2045_addr_0_ack_0 : boolean;
  signal array_obj_ref_2066_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2066_offset_inst_req_0 : boolean;
  signal ptr_deref_2045_addr_0_req_0 : boolean;
  signal array_obj_ref_2090_base_resize_ack_0 : boolean;
  signal binary_1936_inst_req_0 : boolean;
  signal array_obj_ref_2090_base_resize_req_0 : boolean;
  signal binary_1936_inst_ack_0 : boolean;
  signal binary_1936_inst_req_1 : boolean;
  signal binary_1936_inst_ack_1 : boolean;
  signal type_cast_2104_inst_req_0 : boolean;
  signal array_obj_ref_2066_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2090_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2066_index_0_rename_req_0 : boolean;
  signal ptr_deref_2045_root_address_inst_ack_0 : boolean;
  signal binary_2110_inst_ack_1 : boolean;
  signal ptr_deref_2045_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2090_offset_inst_req_0 : boolean;
  signal type_cast_1940_inst_req_0 : boolean;
  signal type_cast_1940_inst_ack_0 : boolean;
  signal binary_2110_inst_req_1 : boolean;
  signal array_obj_ref_2066_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2066_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2114_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2090_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2090_index_0_rename_req_0 : boolean;
  signal ptr_deref_2045_base_resize_ack_0 : boolean;
  signal array_obj_ref_2090_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2090_index_0_resize_req_0 : boolean;
  signal ptr_deref_1943_base_resize_req_0 : boolean;
  signal ptr_deref_1943_base_resize_ack_0 : boolean;
  signal ptr_deref_2045_base_resize_req_0 : boolean;
  signal ptr_deref_1943_root_address_inst_req_0 : boolean;
  signal ptr_deref_1943_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1943_addr_0_req_0 : boolean;
  signal ptr_deref_1943_addr_0_ack_0 : boolean;
  signal array_obj_ref_2114_index_0_resize_req_0 : boolean;
  signal ptr_deref_1943_gather_scatter_req_0 : boolean;
  signal ptr_deref_1943_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2114_final_reg_ack_0 : boolean;
  signal array_obj_ref_2114_final_reg_req_0 : boolean;
  signal ptr_deref_1943_store_0_req_0 : boolean;
  signal ptr_deref_1943_store_0_ack_0 : boolean;
  signal ptr_deref_1943_store_0_req_1 : boolean;
  signal ptr_deref_1943_store_0_ack_1 : boolean;
  signal binary_2110_inst_ack_0 : boolean;
  signal binary_2110_inst_req_0 : boolean;
  signal binary_2086_inst_ack_1 : boolean;
  signal binary_2062_inst_ack_1 : boolean;
  signal binary_2062_inst_req_1 : boolean;
  signal binary_2086_inst_req_1 : boolean;
  signal binary_1950_inst_req_0 : boolean;
  signal binary_2086_inst_ack_0 : boolean;
  signal binary_1950_inst_ack_0 : boolean;
  signal binary_2062_inst_ack_0 : boolean;
  signal binary_2086_inst_req_0 : boolean;
  signal binary_1950_inst_req_1 : boolean;
  signal binary_1950_inst_ack_1 : boolean;
  signal type_cast_1954_inst_req_0 : boolean;
  signal type_cast_1954_inst_ack_0 : boolean;
  signal ptr_deref_1957_base_resize_req_0 : boolean;
  signal ptr_deref_1957_base_resize_ack_0 : boolean;
  signal ptr_deref_1957_root_address_inst_req_0 : boolean;
  signal ptr_deref_1957_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1957_addr_0_req_0 : boolean;
  signal ptr_deref_1957_addr_0_ack_0 : boolean;
  signal ptr_deref_1957_gather_scatter_req_0 : boolean;
  signal ptr_deref_1957_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1957_store_0_req_0 : boolean;
  signal ptr_deref_1957_store_0_ack_0 : boolean;
  signal ptr_deref_1957_store_0_req_1 : boolean;
  signal ptr_deref_1957_store_0_ack_1 : boolean;
  signal binary_1964_inst_req_0 : boolean;
  signal binary_1964_inst_ack_0 : boolean;
  signal binary_1964_inst_req_1 : boolean;
  signal binary_1964_inst_ack_1 : boolean;
  signal type_cast_1968_inst_req_0 : boolean;
  signal type_cast_1968_inst_ack_0 : boolean;
  signal ptr_deref_1971_base_resize_req_0 : boolean;
  signal ptr_deref_1971_base_resize_ack_0 : boolean;
  signal ptr_deref_1971_root_address_inst_req_0 : boolean;
  signal ptr_deref_1971_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1971_addr_0_req_0 : boolean;
  signal ptr_deref_1971_addr_0_ack_0 : boolean;
  signal ptr_deref_1971_gather_scatter_req_0 : boolean;
  signal ptr_deref_1971_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1971_store_0_req_0 : boolean;
  signal ptr_deref_1971_store_0_ack_0 : boolean;
  signal ptr_deref_1971_store_0_req_1 : boolean;
  signal ptr_deref_1971_store_0_ack_1 : boolean;
  signal binary_1978_inst_req_0 : boolean;
  signal binary_1978_inst_ack_0 : boolean;
  signal binary_1978_inst_req_1 : boolean;
  signal binary_1978_inst_ack_1 : boolean;
  signal type_cast_1982_inst_req_0 : boolean;
  signal type_cast_1982_inst_ack_0 : boolean;
  signal ptr_deref_1985_base_resize_req_0 : boolean;
  signal ptr_deref_1985_base_resize_ack_0 : boolean;
  signal ptr_deref_1985_root_address_inst_req_0 : boolean;
  signal ptr_deref_1985_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1985_addr_0_req_0 : boolean;
  signal ptr_deref_1985_addr_0_ack_0 : boolean;
  signal ptr_deref_1985_gather_scatter_req_0 : boolean;
  signal ptr_deref_1985_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1985_store_0_req_0 : boolean;
  signal ptr_deref_1985_store_0_ack_0 : boolean;
  signal ptr_deref_1985_store_0_req_1 : boolean;
  signal ptr_deref_1985_store_0_ack_1 : boolean;
  signal type_cast_1990_inst_req_0 : boolean;
  signal type_cast_1990_inst_ack_0 : boolean;
  signal ptr_deref_1993_base_resize_req_0 : boolean;
  signal ptr_deref_1993_base_resize_ack_0 : boolean;
  signal ptr_deref_1993_root_address_inst_req_0 : boolean;
  signal ptr_deref_1993_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1993_addr_0_req_0 : boolean;
  signal ptr_deref_1993_addr_0_ack_0 : boolean;
  signal ptr_deref_1993_gather_scatter_req_0 : boolean;
  signal ptr_deref_1993_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1993_store_0_req_0 : boolean;
  signal ptr_deref_1993_store_0_ack_0 : boolean;
  signal ptr_deref_1993_store_0_req_1 : boolean;
  signal ptr_deref_1993_store_0_ack_1 : boolean;
  signal binary_2002_inst_req_0 : boolean;
  signal binary_2002_inst_ack_0 : boolean;
  signal binary_2002_inst_req_1 : boolean;
  signal binary_2002_inst_ack_1 : boolean;
  signal binary_2010_inst_req_0 : boolean;
  signal binary_2010_inst_ack_0 : boolean;
  signal binary_2010_inst_req_1 : boolean;
  signal binary_2010_inst_ack_1 : boolean;
  signal type_cast_2014_inst_req_0 : boolean;
  signal type_cast_2014_inst_ack_0 : boolean;
  signal array_obj_ref_2018_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2018_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2018_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2018_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2018_offset_inst_req_0 : boolean;
  signal array_obj_ref_2018_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2018_base_resize_req_0 : boolean;
  signal array_obj_ref_2018_base_resize_ack_0 : boolean;
  signal array_obj_ref_2018_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2018_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2018_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2018_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2018_final_reg_req_0 : boolean;
  signal array_obj_ref_2018_final_reg_ack_0 : boolean;
  signal ptr_deref_2021_base_resize_req_0 : boolean;
  signal ptr_deref_2021_base_resize_ack_0 : boolean;
  signal ptr_deref_2021_root_address_inst_req_0 : boolean;
  signal ptr_deref_2021_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2021_addr_0_req_0 : boolean;
  signal ptr_deref_2021_addr_0_ack_0 : boolean;
  signal ptr_deref_2021_gather_scatter_req_0 : boolean;
  signal ptr_deref_2021_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2021_store_0_req_0 : boolean;
  signal ptr_deref_2021_store_0_ack_0 : boolean;
  signal ptr_deref_2021_store_0_req_1 : boolean;
  signal ptr_deref_2021_store_0_ack_1 : boolean;
  signal binary_2028_inst_req_0 : boolean;
  signal binary_2028_inst_ack_0 : boolean;
  signal binary_2028_inst_req_1 : boolean;
  signal binary_2028_inst_ack_1 : boolean;
  signal type_cast_2032_inst_req_0 : boolean;
  signal type_cast_2032_inst_ack_0 : boolean;
  signal binary_2038_inst_req_0 : boolean;
  signal binary_2038_inst_ack_0 : boolean;
  signal binary_2038_inst_req_1 : boolean;
  signal binary_2038_inst_ack_1 : boolean;
  signal ptr_deref_2117_addr_0_req_0 : boolean;
  signal ptr_deref_2117_addr_0_ack_0 : boolean;
  signal ptr_deref_2117_gather_scatter_req_0 : boolean;
  signal ptr_deref_2117_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2117_store_0_req_0 : boolean;
  signal ptr_deref_2117_store_0_ack_0 : boolean;
  signal ptr_deref_2117_store_0_req_1 : boolean;
  signal ptr_deref_2117_store_0_ack_1 : boolean;
  signal binary_2124_inst_req_0 : boolean;
  signal binary_2124_inst_ack_0 : boolean;
  signal binary_2124_inst_req_1 : boolean;
  signal binary_2124_inst_ack_1 : boolean;
  signal type_cast_2128_inst_req_0 : boolean;
  signal type_cast_2128_inst_ack_0 : boolean;
  signal binary_2134_inst_req_0 : boolean;
  signal binary_2134_inst_ack_0 : boolean;
  signal binary_2134_inst_req_1 : boolean;
  signal binary_2134_inst_ack_1 : boolean;
  signal array_obj_ref_2138_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2138_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2138_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2138_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2138_offset_inst_req_0 : boolean;
  signal array_obj_ref_2138_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2138_base_resize_req_0 : boolean;
  signal array_obj_ref_2138_base_resize_ack_0 : boolean;
  signal array_obj_ref_2138_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2138_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2138_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2138_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2138_final_reg_req_0 : boolean;
  signal array_obj_ref_2138_final_reg_ack_0 : boolean;
  signal phi_stmt_1661_ack_0 : boolean;
  signal ptr_deref_2141_base_resize_req_0 : boolean;
  signal ptr_deref_2141_base_resize_ack_0 : boolean;
  signal ptr_deref_2141_root_address_inst_req_0 : boolean;
  signal ptr_deref_2141_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2141_addr_0_req_0 : boolean;
  signal ptr_deref_2141_addr_0_ack_0 : boolean;
  signal phi_stmt_1661_req_1 : boolean;
  signal ptr_deref_2141_gather_scatter_req_0 : boolean;
  signal ptr_deref_2141_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2141_store_0_req_0 : boolean;
  signal ptr_deref_2141_store_0_ack_0 : boolean;
  signal ptr_deref_2141_store_0_req_1 : boolean;
  signal ptr_deref_2141_store_0_ack_1 : boolean;
  signal type_cast_1667_inst_ack_0 : boolean;
  signal type_cast_1667_inst_req_0 : boolean;
  signal binary_2148_inst_req_0 : boolean;
  signal binary_2148_inst_ack_0 : boolean;
  signal binary_2148_inst_req_1 : boolean;
  signal binary_2148_inst_ack_1 : boolean;
  signal type_cast_2152_inst_req_0 : boolean;
  signal type_cast_2152_inst_ack_0 : boolean;
  signal binary_2158_inst_req_0 : boolean;
  signal binary_2158_inst_ack_0 : boolean;
  signal binary_2158_inst_req_1 : boolean;
  signal binary_2158_inst_ack_1 : boolean;
  signal array_obj_ref_2162_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2162_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2162_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2162_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2162_offset_inst_req_0 : boolean;
  signal array_obj_ref_2162_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2162_base_resize_req_0 : boolean;
  signal array_obj_ref_2162_base_resize_ack_0 : boolean;
  signal array_obj_ref_2162_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2162_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2162_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2162_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2162_final_reg_req_0 : boolean;
  signal array_obj_ref_2162_final_reg_ack_0 : boolean;
  signal ptr_deref_2165_base_resize_req_0 : boolean;
  signal ptr_deref_2165_base_resize_ack_0 : boolean;
  signal ptr_deref_2165_root_address_inst_req_0 : boolean;
  signal ptr_deref_2165_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2165_addr_0_req_0 : boolean;
  signal ptr_deref_2165_addr_0_ack_0 : boolean;
  signal ptr_deref_2165_gather_scatter_req_0 : boolean;
  signal ptr_deref_2165_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2165_store_0_req_0 : boolean;
  signal ptr_deref_2165_store_0_ack_0 : boolean;
  signal ptr_deref_2165_store_0_req_1 : boolean;
  signal ptr_deref_2165_store_0_ack_1 : boolean;
  signal type_cast_2170_inst_req_0 : boolean;
  signal type_cast_2170_inst_ack_0 : boolean;
  signal binary_2176_inst_req_0 : boolean;
  signal binary_2176_inst_ack_0 : boolean;
  signal binary_2176_inst_req_1 : boolean;
  signal binary_2176_inst_ack_1 : boolean;
  signal array_obj_ref_2180_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2180_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2180_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2180_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2180_offset_inst_req_0 : boolean;
  signal array_obj_ref_2180_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2180_base_resize_req_0 : boolean;
  signal array_obj_ref_2180_base_resize_ack_0 : boolean;
  signal array_obj_ref_2180_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2180_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2180_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2180_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2180_final_reg_req_0 : boolean;
  signal array_obj_ref_2180_final_reg_ack_0 : boolean;
  signal ptr_deref_2183_base_resize_req_0 : boolean;
  signal ptr_deref_2183_base_resize_ack_0 : boolean;
  signal ptr_deref_2183_root_address_inst_req_0 : boolean;
  signal ptr_deref_2183_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2183_addr_0_req_0 : boolean;
  signal ptr_deref_2183_addr_0_ack_0 : boolean;
  signal ptr_deref_2183_gather_scatter_req_0 : boolean;
  signal ptr_deref_2183_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2183_store_0_req_0 : boolean;
  signal ptr_deref_2183_store_0_ack_0 : boolean;
  signal ptr_deref_2183_store_0_req_1 : boolean;
  signal ptr_deref_2183_store_0_ack_1 : boolean;
  signal binary_2190_inst_req_0 : boolean;
  signal binary_2190_inst_ack_0 : boolean;
  signal binary_2190_inst_req_1 : boolean;
  signal binary_2190_inst_ack_1 : boolean;
  signal simple_obj_ref_2198_inst_req_0 : boolean;
  signal simple_obj_ref_2198_inst_ack_0 : boolean;
  signal simple_obj_ref_2207_inst_req_0 : boolean;
  signal simple_obj_ref_2207_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_input_CP_6993: Block -- control-path 
    signal cp_elements: BooleanArray(810 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(17);
    simple_obj_ref_1565_inst_req_0 <= cp_elements(2);
    cp_elements(3) <= OrReduce(cp_elements(33) & cp_elements(802));
    simple_obj_ref_1608_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= cp_elements(97);
    phi_stmt_1661_req_0 <= cp_elements(4);
    cp_elements(5) <= OrReduce(cp_elements(125) & cp_elements(808));
    cp_elements(6) <= cp_elements(270);
    cp_elements(7) <= cp_elements(527);
    cp_elements(8) <= cp_elements(795);
    simple_obj_ref_2198_inst_req_0 <= cp_elements(8);
    cp_elements(9) <= cp_elements(0);
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(10) & cp_elements(13));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1554_gather_scatter_req_0 <= cp_elements(11);
    cp_elements(12) <= cp_elements(9);
    cp_elements(13) <= cp_elements(9);
    cp_elements(14) <= ptr_deref_1554_gather_scatter_ack_0;
    ptr_deref_1554_store_0_req_0 <= cp_elements(14);
    cp_elements(15) <= ptr_deref_1554_store_0_ack_0;
    ptr_deref_1554_store_0_req_1 <= cp_elements(15);
    cp_elements(16) <= ptr_deref_1554_store_0_ack_1;
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(16));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(18) <= simple_obj_ref_1565_inst_ack_0;
    cp_elements(19) <= simple_obj_ref_1575_inst_ack_0;
    simple_obj_ref_1586_inst_req_0 <= cp_elements(19);
    cp_elements(20) <= simple_obj_ref_1586_inst_ack_0;
    cp_elements(21) <= cp_elements(20);
    cpelement_group_22 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(23) & cp_elements(24));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(22),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1592_inst_req_0 <= cp_elements(22);
    cp_elements(23) <= cp_elements(21);
    cp_elements(24) <= cp_elements(21);
    cp_elements(25) <= binary_1592_inst_ack_0;
    binary_1592_inst_req_1 <= cp_elements(25);
    cp_elements(26) <= binary_1592_inst_ack_1;
    cp_elements(27) <= cp_elements(26);
    cp_elements(28) <= false;
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= cp_elements(26);
    if_stmt_1594_branch_req_0 <= cp_elements(30);
    cp_elements(31) <= cp_elements(30);
    cp_elements(32) <= cp_elements(31);
    cp_elements(33) <= if_stmt_1594_branch_ack_1;
    cp_elements(34) <= cp_elements(31);
    cp_elements(35) <= if_stmt_1594_branch_ack_0;
    cp_elements(36) <= simple_obj_ref_1608_inst_ack_0;
    cp_elements(37) <= cp_elements(36);
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(39) & cp_elements(40));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1613_inst_req_0 <= cp_elements(38);
    cp_elements(39) <= cp_elements(37);
    cp_elements(40) <= cp_elements(37);
    cp_elements(41) <= type_cast_1613_inst_ack_0;
    array_obj_ref_1638_base_resize_req_0 <= cp_elements(41);
    cpelement_group_42 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(43) & cp_elements(44));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(42),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1618_inst_req_0 <= cp_elements(42);
    cp_elements(43) <= cp_elements(37);
    cp_elements(44) <= cp_elements(37);
    cp_elements(45) <= type_cast_1618_inst_ack_0;
    cp_elements(46) <= cp_elements(37);
    cpelement_group_47 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(46) & cp_elements(51));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(47),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1623_final_reg_req_0 <= cp_elements(47);
    cp_elements(48) <= cp_elements(45);
    array_obj_ref_1623_base_resize_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_1623_base_resize_ack_0;
    array_obj_ref_1623_root_address_inst_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_1623_root_address_inst_ack_0;
    array_obj_ref_1623_root_address_inst_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_1623_root_address_inst_ack_1;
    cp_elements(52) <= array_obj_ref_1623_final_reg_ack_0;
    cp_elements(53) <= cp_elements(37);
    cpelement_group_54 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(58));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(54),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1628_final_reg_req_0 <= cp_elements(54);
    cp_elements(55) <= cp_elements(45);
    array_obj_ref_1628_base_resize_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_1628_base_resize_ack_0;
    array_obj_ref_1628_root_address_inst_req_0 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_1628_root_address_inst_ack_0;
    array_obj_ref_1628_root_address_inst_req_1 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_1628_root_address_inst_ack_1;
    cp_elements(59) <= array_obj_ref_1628_final_reg_ack_0;
    cp_elements(60) <= cp_elements(37);
    cpelement_group_61 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(65));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(61),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1633_final_reg_req_0 <= cp_elements(61);
    cp_elements(62) <= cp_elements(45);
    array_obj_ref_1633_base_resize_req_0 <= cp_elements(62);
    cp_elements(63) <= array_obj_ref_1633_base_resize_ack_0;
    array_obj_ref_1633_root_address_inst_req_0 <= cp_elements(63);
    cp_elements(64) <= array_obj_ref_1633_root_address_inst_ack_0;
    array_obj_ref_1633_root_address_inst_req_1 <= cp_elements(64);
    cp_elements(65) <= array_obj_ref_1633_root_address_inst_ack_1;
    cp_elements(66) <= array_obj_ref_1633_final_reg_ack_0;
    cp_elements(67) <= cp_elements(37);
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(67) & cp_elements(71));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1638_final_reg_req_0 <= cp_elements(68);
    cp_elements(69) <= array_obj_ref_1638_base_resize_ack_0;
    array_obj_ref_1638_root_address_inst_req_0 <= cp_elements(69);
    cp_elements(70) <= array_obj_ref_1638_root_address_inst_ack_0;
    array_obj_ref_1638_root_address_inst_req_1 <= cp_elements(70);
    cp_elements(71) <= array_obj_ref_1638_root_address_inst_ack_1;
    cp_elements(72) <= array_obj_ref_1638_final_reg_ack_0;
    cpelement_group_73 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(72) & cp_elements(74));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(73),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1642_inst_req_0 <= cp_elements(73);
    cp_elements(74) <= cp_elements(37);
    cp_elements(75) <= type_cast_1642_inst_ack_0;
    cp_elements(76) <= cp_elements(37);
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(81));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1647_final_reg_req_0 <= cp_elements(77);
    cp_elements(78) <= cp_elements(45);
    array_obj_ref_1647_base_resize_req_0 <= cp_elements(78);
    cp_elements(79) <= array_obj_ref_1647_base_resize_ack_0;
    array_obj_ref_1647_root_address_inst_req_0 <= cp_elements(79);
    cp_elements(80) <= array_obj_ref_1647_root_address_inst_ack_0;
    array_obj_ref_1647_root_address_inst_req_1 <= cp_elements(80);
    cp_elements(81) <= array_obj_ref_1647_root_address_inst_ack_1;
    cp_elements(82) <= array_obj_ref_1647_final_reg_ack_0;
    cp_elements(83) <= cp_elements(37);
    cpelement_group_84 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(88));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(84),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1652_final_reg_req_0 <= cp_elements(84);
    cp_elements(85) <= cp_elements(45);
    array_obj_ref_1652_base_resize_req_0 <= cp_elements(85);
    cp_elements(86) <= array_obj_ref_1652_base_resize_ack_0;
    array_obj_ref_1652_root_address_inst_req_0 <= cp_elements(86);
    cp_elements(87) <= array_obj_ref_1652_root_address_inst_ack_0;
    array_obj_ref_1652_root_address_inst_req_1 <= cp_elements(87);
    cp_elements(88) <= array_obj_ref_1652_root_address_inst_ack_1;
    cp_elements(89) <= array_obj_ref_1652_final_reg_ack_0;
    cp_elements(90) <= cp_elements(37);
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(90) & cp_elements(95));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1657_final_reg_req_0 <= cp_elements(91);
    cp_elements(92) <= cp_elements(45);
    array_obj_ref_1657_base_resize_req_0 <= cp_elements(92);
    cp_elements(93) <= array_obj_ref_1657_base_resize_ack_0;
    array_obj_ref_1657_root_address_inst_req_0 <= cp_elements(93);
    cp_elements(94) <= array_obj_ref_1657_root_address_inst_ack_0;
    array_obj_ref_1657_root_address_inst_req_1 <= cp_elements(94);
    cp_elements(95) <= array_obj_ref_1657_root_address_inst_ack_1;
    cp_elements(96) <= array_obj_ref_1657_final_reg_ack_0;
    cpelement_group_97 : Block -- 
      signal predecessors: BooleanArray(6 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(52) & cp_elements(59) & cp_elements(66) & cp_elements(75) & cp_elements(82) & cp_elements(89) & cp_elements(96));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(97),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(98) <= cp_elements(806);
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(100) & cp_elements(101));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1673_inst_req_0 <= cp_elements(99);
    cp_elements(100) <= cp_elements(98);
    cp_elements(101) <= cp_elements(98);
    cp_elements(102) <= binary_1673_inst_ack_0;
    binary_1673_inst_req_1 <= cp_elements(102);
    cp_elements(103) <= binary_1673_inst_ack_1;
    simple_obj_ref_1682_inst_req_0 <= cp_elements(103);
    cp_elements(104) <= simple_obj_ref_1682_inst_ack_0;
    simple_obj_ref_1691_inst_req_0 <= cp_elements(104);
    cp_elements(105) <= simple_obj_ref_1691_inst_ack_0;
    cp_elements(106) <= cp_elements(105);
    cpelement_group_107 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(108) & cp_elements(109));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1695_inst_req_0 <= cp_elements(107);
    cp_elements(108) <= cp_elements(106);
    cp_elements(109) <= cp_elements(106);
    cp_elements(110) <= type_cast_1695_inst_ack_0;
    cp_elements(111) <= cp_elements(110);
    cp_elements(112) <= false;
    cp_elements(113) <= cp_elements(112);
    cp_elements(114) <= cp_elements(110);
    cp_elements(115) <= cp_elements(114);
    cp_elements(116) <= cp_elements(115);
    switch_stmt_1697_select_expr_0_req_0 <= cp_elements(116);
    cp_elements(117) <= switch_stmt_1697_select_expr_0_ack_0;
    switch_stmt_1697_select_expr_0_req_1 <= cp_elements(117);
    cp_elements(118) <= switch_stmt_1697_select_expr_0_ack_1;
    switch_stmt_1697_branch_0_req_0 <= cp_elements(118);
    cp_elements(119) <= cp_elements(115);
    switch_stmt_1697_select_expr_1_req_0 <= cp_elements(119);
    cp_elements(120) <= switch_stmt_1697_select_expr_1_ack_0;
    switch_stmt_1697_select_expr_1_req_1 <= cp_elements(120);
    cp_elements(121) <= switch_stmt_1697_select_expr_1_ack_1;
    switch_stmt_1697_branch_1_req_0 <= cp_elements(121);
    cpelement_group_122 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(121));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(122),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    switch_stmt_1697_branch_default_req_0 <= cp_elements(122);
    cp_elements(123) <= cp_elements(122);
    cp_elements(124) <= cp_elements(123);
    cp_elements(125) <= switch_stmt_1697_branch_0_ack_1;
    cp_elements(126) <= cp_elements(123);
    cp_elements(127) <= switch_stmt_1697_branch_1_ack_1;
    cp_elements(128) <= cp_elements(123);
    cp_elements(129) <= switch_stmt_1697_branch_default_ack_0;
    cp_elements(130) <= cp_elements(5);
    cpelement_group_131 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(132) & cp_elements(133));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(131),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1712_inst_req_0 <= cp_elements(131);
    cp_elements(132) <= cp_elements(130);
    cp_elements(133) <= cp_elements(130);
    cp_elements(134) <= binary_1712_inst_ack_0;
    binary_1712_inst_req_1 <= cp_elements(134);
    cp_elements(135) <= binary_1712_inst_ack_1;
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(135) & cp_elements(137));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1716_inst_req_0 <= cp_elements(136);
    cp_elements(137) <= cp_elements(130);
    cp_elements(138) <= type_cast_1716_inst_ack_0;
    cpelement_group_139 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(138) & cp_elements(140) & cp_elements(144));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(139),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1719_gather_scatter_req_0 <= cp_elements(139);
    cp_elements(140) <= cp_elements(130);
    cp_elements(141) <= cp_elements(140);
    ptr_deref_1719_base_resize_req_0 <= cp_elements(141);
    cp_elements(142) <= ptr_deref_1719_base_resize_ack_0;
    ptr_deref_1719_root_address_inst_req_0 <= cp_elements(142);
    cp_elements(143) <= ptr_deref_1719_root_address_inst_ack_0;
    ptr_deref_1719_addr_0_req_0 <= cp_elements(143);
    cp_elements(144) <= ptr_deref_1719_addr_0_ack_0;
    cp_elements(145) <= ptr_deref_1719_gather_scatter_ack_0;
    ptr_deref_1719_store_0_req_0 <= cp_elements(145);
    cp_elements(146) <= ptr_deref_1719_store_0_ack_0;
    cp_elements(147) <= cp_elements(146);
    ptr_deref_1719_store_0_req_1 <= cp_elements(147);
    cp_elements(148) <= ptr_deref_1719_store_0_ack_1;
    cpelement_group_149 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(150) & cp_elements(151));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(149),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1726_inst_req_0 <= cp_elements(149);
    cp_elements(150) <= cp_elements(130);
    cp_elements(151) <= cp_elements(130);
    cp_elements(152) <= binary_1726_inst_ack_0;
    binary_1726_inst_req_1 <= cp_elements(152);
    cp_elements(153) <= binary_1726_inst_ack_1;
    cpelement_group_154 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(153) & cp_elements(155));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(154),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1730_inst_req_0 <= cp_elements(154);
    cp_elements(155) <= cp_elements(130);
    cp_elements(156) <= type_cast_1730_inst_ack_0;
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(146) & cp_elements(156) & cp_elements(158) & cp_elements(162));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1733_gather_scatter_req_0 <= cp_elements(157);
    cp_elements(158) <= cp_elements(130);
    cp_elements(159) <= cp_elements(158);
    ptr_deref_1733_base_resize_req_0 <= cp_elements(159);
    cp_elements(160) <= ptr_deref_1733_base_resize_ack_0;
    ptr_deref_1733_root_address_inst_req_0 <= cp_elements(160);
    cp_elements(161) <= ptr_deref_1733_root_address_inst_ack_0;
    ptr_deref_1733_addr_0_req_0 <= cp_elements(161);
    cp_elements(162) <= ptr_deref_1733_addr_0_ack_0;
    cp_elements(163) <= ptr_deref_1733_gather_scatter_ack_0;
    ptr_deref_1733_store_0_req_0 <= cp_elements(163);
    cp_elements(164) <= ptr_deref_1733_store_0_ack_0;
    cp_elements(165) <= cp_elements(164);
    ptr_deref_1733_store_0_req_1 <= cp_elements(165);
    cp_elements(166) <= ptr_deref_1733_store_0_ack_1;
    cpelement_group_167 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(168) & cp_elements(169));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(167),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1740_inst_req_0 <= cp_elements(167);
    cp_elements(168) <= cp_elements(130);
    cp_elements(169) <= cp_elements(130);
    cp_elements(170) <= binary_1740_inst_ack_0;
    binary_1740_inst_req_1 <= cp_elements(170);
    cp_elements(171) <= binary_1740_inst_ack_1;
    cpelement_group_172 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(171) & cp_elements(173));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(172),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1744_inst_req_0 <= cp_elements(172);
    cp_elements(173) <= cp_elements(130);
    cp_elements(174) <= type_cast_1744_inst_ack_0;
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(164) & cp_elements(174) & cp_elements(176) & cp_elements(180));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1747_gather_scatter_req_0 <= cp_elements(175);
    cp_elements(176) <= cp_elements(130);
    cp_elements(177) <= cp_elements(176);
    ptr_deref_1747_base_resize_req_0 <= cp_elements(177);
    cp_elements(178) <= ptr_deref_1747_base_resize_ack_0;
    ptr_deref_1747_root_address_inst_req_0 <= cp_elements(178);
    cp_elements(179) <= ptr_deref_1747_root_address_inst_ack_0;
    ptr_deref_1747_addr_0_req_0 <= cp_elements(179);
    cp_elements(180) <= ptr_deref_1747_addr_0_ack_0;
    cp_elements(181) <= ptr_deref_1747_gather_scatter_ack_0;
    ptr_deref_1747_store_0_req_0 <= cp_elements(181);
    cp_elements(182) <= ptr_deref_1747_store_0_ack_0;
    cp_elements(183) <= cp_elements(182);
    ptr_deref_1747_store_0_req_1 <= cp_elements(183);
    cp_elements(184) <= ptr_deref_1747_store_0_ack_1;
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(187));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1754_inst_req_0 <= cp_elements(185);
    cp_elements(186) <= cp_elements(130);
    cp_elements(187) <= cp_elements(130);
    cp_elements(188) <= binary_1754_inst_ack_0;
    binary_1754_inst_req_1 <= cp_elements(188);
    cp_elements(189) <= binary_1754_inst_ack_1;
    cpelement_group_190 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(189) & cp_elements(191));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(190),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1758_inst_req_0 <= cp_elements(190);
    cp_elements(191) <= cp_elements(130);
    cp_elements(192) <= type_cast_1758_inst_ack_0;
    cpelement_group_193 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(182) & cp_elements(192) & cp_elements(194) & cp_elements(198));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(193),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1761_gather_scatter_req_0 <= cp_elements(193);
    cp_elements(194) <= cp_elements(130);
    cp_elements(195) <= cp_elements(194);
    ptr_deref_1761_base_resize_req_0 <= cp_elements(195);
    cp_elements(196) <= ptr_deref_1761_base_resize_ack_0;
    ptr_deref_1761_root_address_inst_req_0 <= cp_elements(196);
    cp_elements(197) <= ptr_deref_1761_root_address_inst_ack_0;
    ptr_deref_1761_addr_0_req_0 <= cp_elements(197);
    cp_elements(198) <= ptr_deref_1761_addr_0_ack_0;
    cp_elements(199) <= ptr_deref_1761_gather_scatter_ack_0;
    ptr_deref_1761_store_0_req_0 <= cp_elements(199);
    cp_elements(200) <= ptr_deref_1761_store_0_ack_0;
    cp_elements(201) <= cp_elements(200);
    ptr_deref_1761_store_0_req_1 <= cp_elements(201);
    cp_elements(202) <= ptr_deref_1761_store_0_ack_1;
    cpelement_group_203 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(204) & cp_elements(205));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(203),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1768_inst_req_0 <= cp_elements(203);
    cp_elements(204) <= cp_elements(130);
    cp_elements(205) <= cp_elements(130);
    cp_elements(206) <= binary_1768_inst_ack_0;
    binary_1768_inst_req_1 <= cp_elements(206);
    cp_elements(207) <= binary_1768_inst_ack_1;
    cpelement_group_208 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(207) & cp_elements(209));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(208),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1772_inst_req_0 <= cp_elements(208);
    cp_elements(209) <= cp_elements(130);
    cp_elements(210) <= type_cast_1772_inst_ack_0;
    cpelement_group_211 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(200) & cp_elements(210) & cp_elements(212) & cp_elements(216));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1775_gather_scatter_req_0 <= cp_elements(211);
    cp_elements(212) <= cp_elements(130);
    cp_elements(213) <= cp_elements(212);
    ptr_deref_1775_base_resize_req_0 <= cp_elements(213);
    cp_elements(214) <= ptr_deref_1775_base_resize_ack_0;
    ptr_deref_1775_root_address_inst_req_0 <= cp_elements(214);
    cp_elements(215) <= ptr_deref_1775_root_address_inst_ack_0;
    ptr_deref_1775_addr_0_req_0 <= cp_elements(215);
    cp_elements(216) <= ptr_deref_1775_addr_0_ack_0;
    cp_elements(217) <= ptr_deref_1775_gather_scatter_ack_0;
    ptr_deref_1775_store_0_req_0 <= cp_elements(217);
    cp_elements(218) <= ptr_deref_1775_store_0_ack_0;
    cp_elements(219) <= cp_elements(218);
    ptr_deref_1775_store_0_req_1 <= cp_elements(219);
    cp_elements(220) <= ptr_deref_1775_store_0_ack_1;
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(222) & cp_elements(223));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1782_inst_req_0 <= cp_elements(221);
    cp_elements(222) <= cp_elements(130);
    cp_elements(223) <= cp_elements(130);
    cp_elements(224) <= binary_1782_inst_ack_0;
    binary_1782_inst_req_1 <= cp_elements(224);
    cp_elements(225) <= binary_1782_inst_ack_1;
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(225) & cp_elements(227));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1786_inst_req_0 <= cp_elements(226);
    cp_elements(227) <= cp_elements(130);
    cp_elements(228) <= type_cast_1786_inst_ack_0;
    cpelement_group_229 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(228) & cp_elements(230) & cp_elements(234));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(229),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1789_gather_scatter_req_0 <= cp_elements(229);
    cp_elements(230) <= cp_elements(130);
    cp_elements(231) <= cp_elements(230);
    ptr_deref_1789_base_resize_req_0 <= cp_elements(231);
    cp_elements(232) <= ptr_deref_1789_base_resize_ack_0;
    ptr_deref_1789_root_address_inst_req_0 <= cp_elements(232);
    cp_elements(233) <= ptr_deref_1789_root_address_inst_ack_0;
    ptr_deref_1789_addr_0_req_0 <= cp_elements(233);
    cp_elements(234) <= ptr_deref_1789_addr_0_ack_0;
    cp_elements(235) <= ptr_deref_1789_gather_scatter_ack_0;
    ptr_deref_1789_store_0_req_0 <= cp_elements(235);
    cp_elements(236) <= ptr_deref_1789_store_0_ack_0;
    cp_elements(237) <= cp_elements(236);
    ptr_deref_1789_store_0_req_1 <= cp_elements(237);
    cp_elements(238) <= ptr_deref_1789_store_0_ack_1;
    cpelement_group_239 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(240) & cp_elements(241));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(239),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1796_inst_req_0 <= cp_elements(239);
    cp_elements(240) <= cp_elements(130);
    cp_elements(241) <= cp_elements(130);
    cp_elements(242) <= binary_1796_inst_ack_0;
    binary_1796_inst_req_1 <= cp_elements(242);
    cp_elements(243) <= binary_1796_inst_ack_1;
    cpelement_group_244 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(243) & cp_elements(245));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(244),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1800_inst_req_0 <= cp_elements(244);
    cp_elements(245) <= cp_elements(130);
    cp_elements(246) <= type_cast_1800_inst_ack_0;
    cpelement_group_247 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(236) & cp_elements(246) & cp_elements(248) & cp_elements(252));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(247),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1803_gather_scatter_req_0 <= cp_elements(247);
    cp_elements(248) <= cp_elements(130);
    cp_elements(249) <= cp_elements(248);
    ptr_deref_1803_base_resize_req_0 <= cp_elements(249);
    cp_elements(250) <= ptr_deref_1803_base_resize_ack_0;
    ptr_deref_1803_root_address_inst_req_0 <= cp_elements(250);
    cp_elements(251) <= ptr_deref_1803_root_address_inst_ack_0;
    ptr_deref_1803_addr_0_req_0 <= cp_elements(251);
    cp_elements(252) <= ptr_deref_1803_addr_0_ack_0;
    cp_elements(253) <= ptr_deref_1803_gather_scatter_ack_0;
    ptr_deref_1803_store_0_req_0 <= cp_elements(253);
    cp_elements(254) <= ptr_deref_1803_store_0_ack_0;
    cp_elements(255) <= cp_elements(254);
    ptr_deref_1803_store_0_req_1 <= cp_elements(255);
    cp_elements(256) <= ptr_deref_1803_store_0_ack_1;
    cpelement_group_257 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(258) & cp_elements(259));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(257),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1808_inst_req_0 <= cp_elements(257);
    cp_elements(258) <= cp_elements(130);
    cp_elements(259) <= cp_elements(130);
    cp_elements(260) <= type_cast_1808_inst_ack_0;
    cpelement_group_261 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(260) & cp_elements(262) & cp_elements(266));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(261),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1811_gather_scatter_req_0 <= cp_elements(261);
    cp_elements(262) <= cp_elements(130);
    cp_elements(263) <= cp_elements(262);
    ptr_deref_1811_base_resize_req_0 <= cp_elements(263);
    cp_elements(264) <= ptr_deref_1811_base_resize_ack_0;
    ptr_deref_1811_root_address_inst_req_0 <= cp_elements(264);
    cp_elements(265) <= ptr_deref_1811_root_address_inst_ack_0;
    ptr_deref_1811_addr_0_req_0 <= cp_elements(265);
    cp_elements(266) <= ptr_deref_1811_addr_0_ack_0;
    cp_elements(267) <= ptr_deref_1811_gather_scatter_ack_0;
    ptr_deref_1811_store_0_req_0 <= cp_elements(267);
    cp_elements(268) <= ptr_deref_1811_store_0_ack_0;
    ptr_deref_1811_store_0_req_1 <= cp_elements(268);
    cp_elements(269) <= ptr_deref_1811_store_0_ack_1;
    cpelement_group_270 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(166) & cp_elements(184) & cp_elements(202) & cp_elements(220) & cp_elements(238) & cp_elements(256) & cp_elements(269));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(270),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(271) <= cp_elements(127);
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(273) & cp_elements(274));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1820_inst_req_0 <= cp_elements(272);
    cp_elements(273) <= cp_elements(271);
    cp_elements(274) <= cp_elements(271);
    cp_elements(275) <= binary_1820_inst_ack_0;
    binary_1820_inst_req_1 <= cp_elements(275);
    cp_elements(276) <= binary_1820_inst_ack_1;
    array_obj_ref_1864_index_0_resize_req_0 <= cp_elements(276);
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(278) & cp_elements(279));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1826_inst_req_0 <= cp_elements(277);
    cp_elements(278) <= cp_elements(271);
    cp_elements(279) <= cp_elements(271);
    cp_elements(280) <= binary_1826_inst_ack_0;
    binary_1826_inst_req_1 <= cp_elements(280);
    cp_elements(281) <= binary_1826_inst_ack_1;
    array_obj_ref_1868_index_0_resize_req_0 <= cp_elements(281);
    cpelement_group_282 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(284));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(282),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1832_inst_req_0 <= cp_elements(282);
    cp_elements(283) <= cp_elements(271);
    cp_elements(284) <= cp_elements(271);
    cp_elements(285) <= binary_1832_inst_ack_0;
    binary_1832_inst_req_1 <= cp_elements(285);
    cp_elements(286) <= binary_1832_inst_ack_1;
    array_obj_ref_1872_index_0_resize_req_0 <= cp_elements(286);
    cpelement_group_287 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(288) & cp_elements(289));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(287),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1838_inst_req_0 <= cp_elements(287);
    cp_elements(288) <= cp_elements(271);
    cp_elements(289) <= cp_elements(271);
    cp_elements(290) <= binary_1838_inst_ack_0;
    binary_1838_inst_req_1 <= cp_elements(290);
    cp_elements(291) <= binary_1838_inst_ack_1;
    array_obj_ref_1876_index_0_resize_req_0 <= cp_elements(291);
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(293) & cp_elements(294));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1844_inst_req_0 <= cp_elements(292);
    cp_elements(293) <= cp_elements(271);
    cp_elements(294) <= cp_elements(271);
    cp_elements(295) <= binary_1844_inst_ack_0;
    binary_1844_inst_req_1 <= cp_elements(295);
    cp_elements(296) <= binary_1844_inst_ack_1;
    array_obj_ref_1880_index_0_resize_req_0 <= cp_elements(296);
    cpelement_group_297 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(298) & cp_elements(299));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(297),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1850_inst_req_0 <= cp_elements(297);
    cp_elements(298) <= cp_elements(271);
    cp_elements(299) <= cp_elements(271);
    cp_elements(300) <= binary_1850_inst_ack_0;
    binary_1850_inst_req_1 <= cp_elements(300);
    cp_elements(301) <= binary_1850_inst_ack_1;
    array_obj_ref_1884_index_0_resize_req_0 <= cp_elements(301);
    cpelement_group_302 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(303) & cp_elements(304));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(302),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1856_inst_req_0 <= cp_elements(302);
    cp_elements(303) <= cp_elements(271);
    cp_elements(304) <= cp_elements(271);
    cp_elements(305) <= binary_1856_inst_ack_0;
    binary_1856_inst_req_1 <= cp_elements(305);
    cp_elements(306) <= binary_1856_inst_ack_1;
    array_obj_ref_1888_index_0_resize_req_0 <= cp_elements(306);
    cp_elements(307) <= cp_elements(271);
    cpelement_group_308 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(307) & cp_elements(317));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1860_final_reg_req_0 <= cp_elements(308);
    cp_elements(309) <= cp_elements(271);
    array_obj_ref_1860_base_resize_req_0 <= cp_elements(309);
    cp_elements(310) <= cp_elements(271);
    array_obj_ref_1860_index_0_resize_req_0 <= cp_elements(310);
    cp_elements(311) <= array_obj_ref_1860_index_0_resize_ack_0;
    array_obj_ref_1860_index_0_rename_req_0 <= cp_elements(311);
    cp_elements(312) <= array_obj_ref_1860_index_0_rename_ack_0;
    array_obj_ref_1860_offset_inst_req_0 <= cp_elements(312);
    cp_elements(313) <= array_obj_ref_1860_offset_inst_ack_0;
    cp_elements(314) <= array_obj_ref_1860_base_resize_ack_0;
    cpelement_group_315 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(314));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(315),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1860_root_address_inst_req_0 <= cp_elements(315);
    cp_elements(316) <= array_obj_ref_1860_root_address_inst_ack_0;
    array_obj_ref_1860_root_address_inst_req_1 <= cp_elements(316);
    cp_elements(317) <= array_obj_ref_1860_root_address_inst_ack_1;
    cp_elements(318) <= array_obj_ref_1860_final_reg_ack_0;
    cp_elements(319) <= cp_elements(271);
    cpelement_group_320 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(319) & cp_elements(328));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(320),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1864_final_reg_req_0 <= cp_elements(320);
    cp_elements(321) <= cp_elements(271);
    array_obj_ref_1864_base_resize_req_0 <= cp_elements(321);
    cp_elements(322) <= array_obj_ref_1864_index_0_resize_ack_0;
    array_obj_ref_1864_index_0_rename_req_0 <= cp_elements(322);
    cp_elements(323) <= array_obj_ref_1864_index_0_rename_ack_0;
    array_obj_ref_1864_offset_inst_req_0 <= cp_elements(323);
    cp_elements(324) <= array_obj_ref_1864_offset_inst_ack_0;
    cp_elements(325) <= array_obj_ref_1864_base_resize_ack_0;
    cpelement_group_326 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(324) & cp_elements(325));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(326),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1864_root_address_inst_req_0 <= cp_elements(326);
    cp_elements(327) <= array_obj_ref_1864_root_address_inst_ack_0;
    array_obj_ref_1864_root_address_inst_req_1 <= cp_elements(327);
    cp_elements(328) <= array_obj_ref_1864_root_address_inst_ack_1;
    cp_elements(329) <= array_obj_ref_1864_final_reg_ack_0;
    cp_elements(330) <= cp_elements(271);
    cpelement_group_331 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(330) & cp_elements(339));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(331),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1868_final_reg_req_0 <= cp_elements(331);
    cp_elements(332) <= cp_elements(271);
    array_obj_ref_1868_base_resize_req_0 <= cp_elements(332);
    cp_elements(333) <= array_obj_ref_1868_index_0_resize_ack_0;
    array_obj_ref_1868_index_0_rename_req_0 <= cp_elements(333);
    cp_elements(334) <= array_obj_ref_1868_index_0_rename_ack_0;
    array_obj_ref_1868_offset_inst_req_0 <= cp_elements(334);
    cp_elements(335) <= array_obj_ref_1868_offset_inst_ack_0;
    cp_elements(336) <= array_obj_ref_1868_base_resize_ack_0;
    cpelement_group_337 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(335) & cp_elements(336));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(337),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1868_root_address_inst_req_0 <= cp_elements(337);
    cp_elements(338) <= array_obj_ref_1868_root_address_inst_ack_0;
    array_obj_ref_1868_root_address_inst_req_1 <= cp_elements(338);
    cp_elements(339) <= array_obj_ref_1868_root_address_inst_ack_1;
    cp_elements(340) <= array_obj_ref_1868_final_reg_ack_0;
    cp_elements(341) <= cp_elements(271);
    cpelement_group_342 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(341) & cp_elements(350));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(342),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1872_final_reg_req_0 <= cp_elements(342);
    cp_elements(343) <= cp_elements(271);
    array_obj_ref_1872_base_resize_req_0 <= cp_elements(343);
    cp_elements(344) <= array_obj_ref_1872_index_0_resize_ack_0;
    array_obj_ref_1872_index_0_rename_req_0 <= cp_elements(344);
    cp_elements(345) <= array_obj_ref_1872_index_0_rename_ack_0;
    array_obj_ref_1872_offset_inst_req_0 <= cp_elements(345);
    cp_elements(346) <= array_obj_ref_1872_offset_inst_ack_0;
    cp_elements(347) <= array_obj_ref_1872_base_resize_ack_0;
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(346) & cp_elements(347));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1872_root_address_inst_req_0 <= cp_elements(348);
    cp_elements(349) <= array_obj_ref_1872_root_address_inst_ack_0;
    array_obj_ref_1872_root_address_inst_req_1 <= cp_elements(349);
    cp_elements(350) <= array_obj_ref_1872_root_address_inst_ack_1;
    cp_elements(351) <= array_obj_ref_1872_final_reg_ack_0;
    cp_elements(352) <= cp_elements(271);
    cpelement_group_353 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(352) & cp_elements(361));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(353),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1876_final_reg_req_0 <= cp_elements(353);
    cp_elements(354) <= cp_elements(271);
    array_obj_ref_1876_base_resize_req_0 <= cp_elements(354);
    cp_elements(355) <= array_obj_ref_1876_index_0_resize_ack_0;
    array_obj_ref_1876_index_0_rename_req_0 <= cp_elements(355);
    cp_elements(356) <= array_obj_ref_1876_index_0_rename_ack_0;
    array_obj_ref_1876_offset_inst_req_0 <= cp_elements(356);
    cp_elements(357) <= array_obj_ref_1876_offset_inst_ack_0;
    cp_elements(358) <= array_obj_ref_1876_base_resize_ack_0;
    cpelement_group_359 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(357) & cp_elements(358));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(359),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1876_root_address_inst_req_0 <= cp_elements(359);
    cp_elements(360) <= array_obj_ref_1876_root_address_inst_ack_0;
    array_obj_ref_1876_root_address_inst_req_1 <= cp_elements(360);
    cp_elements(361) <= array_obj_ref_1876_root_address_inst_ack_1;
    cp_elements(362) <= array_obj_ref_1876_final_reg_ack_0;
    cp_elements(363) <= cp_elements(271);
    cpelement_group_364 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(363) & cp_elements(372));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1880_final_reg_req_0 <= cp_elements(364);
    cp_elements(365) <= cp_elements(271);
    array_obj_ref_1880_base_resize_req_0 <= cp_elements(365);
    cp_elements(366) <= array_obj_ref_1880_index_0_resize_ack_0;
    array_obj_ref_1880_index_0_rename_req_0 <= cp_elements(366);
    cp_elements(367) <= array_obj_ref_1880_index_0_rename_ack_0;
    array_obj_ref_1880_offset_inst_req_0 <= cp_elements(367);
    cp_elements(368) <= array_obj_ref_1880_offset_inst_ack_0;
    cp_elements(369) <= array_obj_ref_1880_base_resize_ack_0;
    cpelement_group_370 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(368) & cp_elements(369));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(370),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1880_root_address_inst_req_0 <= cp_elements(370);
    cp_elements(371) <= array_obj_ref_1880_root_address_inst_ack_0;
    array_obj_ref_1880_root_address_inst_req_1 <= cp_elements(371);
    cp_elements(372) <= array_obj_ref_1880_root_address_inst_ack_1;
    cp_elements(373) <= array_obj_ref_1880_final_reg_ack_0;
    cp_elements(374) <= cp_elements(271);
    cpelement_group_375 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(374) & cp_elements(383));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(375),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1884_final_reg_req_0 <= cp_elements(375);
    cp_elements(376) <= cp_elements(271);
    array_obj_ref_1884_base_resize_req_0 <= cp_elements(376);
    cp_elements(377) <= array_obj_ref_1884_index_0_resize_ack_0;
    array_obj_ref_1884_index_0_rename_req_0 <= cp_elements(377);
    cp_elements(378) <= array_obj_ref_1884_index_0_rename_ack_0;
    array_obj_ref_1884_offset_inst_req_0 <= cp_elements(378);
    cp_elements(379) <= array_obj_ref_1884_offset_inst_ack_0;
    cp_elements(380) <= array_obj_ref_1884_base_resize_ack_0;
    cpelement_group_381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(379) & cp_elements(380));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1884_root_address_inst_req_0 <= cp_elements(381);
    cp_elements(382) <= array_obj_ref_1884_root_address_inst_ack_0;
    array_obj_ref_1884_root_address_inst_req_1 <= cp_elements(382);
    cp_elements(383) <= array_obj_ref_1884_root_address_inst_ack_1;
    cp_elements(384) <= array_obj_ref_1884_final_reg_ack_0;
    cp_elements(385) <= cp_elements(271);
    cpelement_group_386 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(385) & cp_elements(394));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1888_final_reg_req_0 <= cp_elements(386);
    cp_elements(387) <= cp_elements(271);
    array_obj_ref_1888_base_resize_req_0 <= cp_elements(387);
    cp_elements(388) <= array_obj_ref_1888_index_0_resize_ack_0;
    array_obj_ref_1888_index_0_rename_req_0 <= cp_elements(388);
    cp_elements(389) <= array_obj_ref_1888_index_0_rename_ack_0;
    array_obj_ref_1888_offset_inst_req_0 <= cp_elements(389);
    cp_elements(390) <= array_obj_ref_1888_offset_inst_ack_0;
    cp_elements(391) <= array_obj_ref_1888_base_resize_ack_0;
    cpelement_group_392 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(390) & cp_elements(391));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(392),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1888_root_address_inst_req_0 <= cp_elements(392);
    cp_elements(393) <= array_obj_ref_1888_root_address_inst_ack_0;
    array_obj_ref_1888_root_address_inst_req_1 <= cp_elements(393);
    cp_elements(394) <= array_obj_ref_1888_root_address_inst_ack_1;
    cp_elements(395) <= array_obj_ref_1888_final_reg_ack_0;
    cpelement_group_396 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(397) & cp_elements(398));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(396),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1894_inst_req_0 <= cp_elements(396);
    cp_elements(397) <= cp_elements(271);
    cp_elements(398) <= cp_elements(271);
    cp_elements(399) <= binary_1894_inst_ack_0;
    binary_1894_inst_req_1 <= cp_elements(399);
    cp_elements(400) <= binary_1894_inst_ack_1;
    cpelement_group_401 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(400) & cp_elements(402));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(401),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1898_inst_req_0 <= cp_elements(401);
    cp_elements(402) <= cp_elements(271);
    cp_elements(403) <= type_cast_1898_inst_ack_0;
    cpelement_group_404 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(318) & cp_elements(403) & cp_elements(408));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(404),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1901_gather_scatter_req_0 <= cp_elements(404);
    cp_elements(405) <= cp_elements(318);
    ptr_deref_1901_base_resize_req_0 <= cp_elements(405);
    cp_elements(406) <= ptr_deref_1901_base_resize_ack_0;
    ptr_deref_1901_root_address_inst_req_0 <= cp_elements(406);
    cp_elements(407) <= ptr_deref_1901_root_address_inst_ack_0;
    ptr_deref_1901_addr_0_req_0 <= cp_elements(407);
    cp_elements(408) <= ptr_deref_1901_addr_0_ack_0;
    cp_elements(409) <= ptr_deref_1901_gather_scatter_ack_0;
    ptr_deref_1901_store_0_req_0 <= cp_elements(409);
    cp_elements(410) <= ptr_deref_1901_store_0_ack_0;
    cp_elements(411) <= cp_elements(410);
    ptr_deref_1901_store_0_req_1 <= cp_elements(411);
    cp_elements(412) <= ptr_deref_1901_store_0_ack_1;
    cpelement_group_413 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(414) & cp_elements(415));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(413),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1908_inst_req_0 <= cp_elements(413);
    cp_elements(414) <= cp_elements(271);
    cp_elements(415) <= cp_elements(271);
    cp_elements(416) <= binary_1908_inst_ack_0;
    binary_1908_inst_req_1 <= cp_elements(416);
    cp_elements(417) <= binary_1908_inst_ack_1;
    cpelement_group_418 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(417) & cp_elements(419));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(418),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1912_inst_req_0 <= cp_elements(418);
    cp_elements(419) <= cp_elements(271);
    cp_elements(420) <= type_cast_1912_inst_ack_0;
    cpelement_group_421 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(329) & cp_elements(410) & cp_elements(420) & cp_elements(425));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(421),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1915_gather_scatter_req_0 <= cp_elements(421);
    cp_elements(422) <= cp_elements(329);
    ptr_deref_1915_base_resize_req_0 <= cp_elements(422);
    cp_elements(423) <= ptr_deref_1915_base_resize_ack_0;
    ptr_deref_1915_root_address_inst_req_0 <= cp_elements(423);
    cp_elements(424) <= ptr_deref_1915_root_address_inst_ack_0;
    ptr_deref_1915_addr_0_req_0 <= cp_elements(424);
    cp_elements(425) <= ptr_deref_1915_addr_0_ack_0;
    cp_elements(426) <= ptr_deref_1915_gather_scatter_ack_0;
    ptr_deref_1915_store_0_req_0 <= cp_elements(426);
    cp_elements(427) <= ptr_deref_1915_store_0_ack_0;
    cp_elements(428) <= cp_elements(427);
    ptr_deref_1915_store_0_req_1 <= cp_elements(428);
    cp_elements(429) <= ptr_deref_1915_store_0_ack_1;
    cpelement_group_430 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(431) & cp_elements(432));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(430),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1922_inst_req_0 <= cp_elements(430);
    cp_elements(431) <= cp_elements(271);
    cp_elements(432) <= cp_elements(271);
    cp_elements(433) <= binary_1922_inst_ack_0;
    binary_1922_inst_req_1 <= cp_elements(433);
    cp_elements(434) <= binary_1922_inst_ack_1;
    cpelement_group_435 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(434) & cp_elements(436));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(435),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1926_inst_req_0 <= cp_elements(435);
    cp_elements(436) <= cp_elements(271);
    cp_elements(437) <= type_cast_1926_inst_ack_0;
    cpelement_group_438 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(340) & cp_elements(427) & cp_elements(437) & cp_elements(442));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(438),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1929_gather_scatter_req_0 <= cp_elements(438);
    cp_elements(439) <= cp_elements(340);
    ptr_deref_1929_base_resize_req_0 <= cp_elements(439);
    cp_elements(440) <= ptr_deref_1929_base_resize_ack_0;
    ptr_deref_1929_root_address_inst_req_0 <= cp_elements(440);
    cp_elements(441) <= ptr_deref_1929_root_address_inst_ack_0;
    ptr_deref_1929_addr_0_req_0 <= cp_elements(441);
    cp_elements(442) <= ptr_deref_1929_addr_0_ack_0;
    cp_elements(443) <= ptr_deref_1929_gather_scatter_ack_0;
    ptr_deref_1929_store_0_req_0 <= cp_elements(443);
    cp_elements(444) <= ptr_deref_1929_store_0_ack_0;
    cp_elements(445) <= cp_elements(444);
    ptr_deref_1929_store_0_req_1 <= cp_elements(445);
    cp_elements(446) <= ptr_deref_1929_store_0_ack_1;
    cpelement_group_447 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(448) & cp_elements(449));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(447),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1936_inst_req_0 <= cp_elements(447);
    cp_elements(448) <= cp_elements(271);
    cp_elements(449) <= cp_elements(271);
    cp_elements(450) <= binary_1936_inst_ack_0;
    binary_1936_inst_req_1 <= cp_elements(450);
    cp_elements(451) <= binary_1936_inst_ack_1;
    cpelement_group_452 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(451) & cp_elements(453));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(452),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1940_inst_req_0 <= cp_elements(452);
    cp_elements(453) <= cp_elements(271);
    cp_elements(454) <= type_cast_1940_inst_ack_0;
    cpelement_group_455 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(351) & cp_elements(444) & cp_elements(454) & cp_elements(459));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(455),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1943_gather_scatter_req_0 <= cp_elements(455);
    cp_elements(456) <= cp_elements(351);
    ptr_deref_1943_base_resize_req_0 <= cp_elements(456);
    cp_elements(457) <= ptr_deref_1943_base_resize_ack_0;
    ptr_deref_1943_root_address_inst_req_0 <= cp_elements(457);
    cp_elements(458) <= ptr_deref_1943_root_address_inst_ack_0;
    ptr_deref_1943_addr_0_req_0 <= cp_elements(458);
    cp_elements(459) <= ptr_deref_1943_addr_0_ack_0;
    cp_elements(460) <= ptr_deref_1943_gather_scatter_ack_0;
    ptr_deref_1943_store_0_req_0 <= cp_elements(460);
    cp_elements(461) <= ptr_deref_1943_store_0_ack_0;
    cp_elements(462) <= cp_elements(461);
    ptr_deref_1943_store_0_req_1 <= cp_elements(462);
    cp_elements(463) <= ptr_deref_1943_store_0_ack_1;
    cpelement_group_464 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(465) & cp_elements(466));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(464),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1950_inst_req_0 <= cp_elements(464);
    cp_elements(465) <= cp_elements(271);
    cp_elements(466) <= cp_elements(271);
    cp_elements(467) <= binary_1950_inst_ack_0;
    binary_1950_inst_req_1 <= cp_elements(467);
    cp_elements(468) <= binary_1950_inst_ack_1;
    cpelement_group_469 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(468) & cp_elements(470));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(469),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1954_inst_req_0 <= cp_elements(469);
    cp_elements(470) <= cp_elements(271);
    cp_elements(471) <= type_cast_1954_inst_ack_0;
    cpelement_group_472 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(362) & cp_elements(461) & cp_elements(471) & cp_elements(476));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(472),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1957_gather_scatter_req_0 <= cp_elements(472);
    cp_elements(473) <= cp_elements(362);
    ptr_deref_1957_base_resize_req_0 <= cp_elements(473);
    cp_elements(474) <= ptr_deref_1957_base_resize_ack_0;
    ptr_deref_1957_root_address_inst_req_0 <= cp_elements(474);
    cp_elements(475) <= ptr_deref_1957_root_address_inst_ack_0;
    ptr_deref_1957_addr_0_req_0 <= cp_elements(475);
    cp_elements(476) <= ptr_deref_1957_addr_0_ack_0;
    cp_elements(477) <= ptr_deref_1957_gather_scatter_ack_0;
    ptr_deref_1957_store_0_req_0 <= cp_elements(477);
    cp_elements(478) <= ptr_deref_1957_store_0_ack_0;
    cp_elements(479) <= cp_elements(478);
    ptr_deref_1957_store_0_req_1 <= cp_elements(479);
    cp_elements(480) <= ptr_deref_1957_store_0_ack_1;
    cpelement_group_481 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(482) & cp_elements(483));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(481),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1964_inst_req_0 <= cp_elements(481);
    cp_elements(482) <= cp_elements(271);
    cp_elements(483) <= cp_elements(271);
    cp_elements(484) <= binary_1964_inst_ack_0;
    binary_1964_inst_req_1 <= cp_elements(484);
    cp_elements(485) <= binary_1964_inst_ack_1;
    cpelement_group_486 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(485) & cp_elements(487));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(486),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1968_inst_req_0 <= cp_elements(486);
    cp_elements(487) <= cp_elements(271);
    cp_elements(488) <= type_cast_1968_inst_ack_0;
    cpelement_group_489 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(373) & cp_elements(478) & cp_elements(488) & cp_elements(493));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(489),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1971_gather_scatter_req_0 <= cp_elements(489);
    cp_elements(490) <= cp_elements(373);
    ptr_deref_1971_base_resize_req_0 <= cp_elements(490);
    cp_elements(491) <= ptr_deref_1971_base_resize_ack_0;
    ptr_deref_1971_root_address_inst_req_0 <= cp_elements(491);
    cp_elements(492) <= ptr_deref_1971_root_address_inst_ack_0;
    ptr_deref_1971_addr_0_req_0 <= cp_elements(492);
    cp_elements(493) <= ptr_deref_1971_addr_0_ack_0;
    cp_elements(494) <= ptr_deref_1971_gather_scatter_ack_0;
    ptr_deref_1971_store_0_req_0 <= cp_elements(494);
    cp_elements(495) <= ptr_deref_1971_store_0_ack_0;
    cp_elements(496) <= cp_elements(495);
    ptr_deref_1971_store_0_req_1 <= cp_elements(496);
    cp_elements(497) <= ptr_deref_1971_store_0_ack_1;
    cpelement_group_498 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(499) & cp_elements(500));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(498),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1978_inst_req_0 <= cp_elements(498);
    cp_elements(499) <= cp_elements(271);
    cp_elements(500) <= cp_elements(271);
    cp_elements(501) <= binary_1978_inst_ack_0;
    binary_1978_inst_req_1 <= cp_elements(501);
    cp_elements(502) <= binary_1978_inst_ack_1;
    cpelement_group_503 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(502) & cp_elements(504));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(503),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1982_inst_req_0 <= cp_elements(503);
    cp_elements(504) <= cp_elements(271);
    cp_elements(505) <= type_cast_1982_inst_ack_0;
    cpelement_group_506 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(384) & cp_elements(495) & cp_elements(505) & cp_elements(510));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(506),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1985_gather_scatter_req_0 <= cp_elements(506);
    cp_elements(507) <= cp_elements(384);
    ptr_deref_1985_base_resize_req_0 <= cp_elements(507);
    cp_elements(508) <= ptr_deref_1985_base_resize_ack_0;
    ptr_deref_1985_root_address_inst_req_0 <= cp_elements(508);
    cp_elements(509) <= ptr_deref_1985_root_address_inst_ack_0;
    ptr_deref_1985_addr_0_req_0 <= cp_elements(509);
    cp_elements(510) <= ptr_deref_1985_addr_0_ack_0;
    cp_elements(511) <= ptr_deref_1985_gather_scatter_ack_0;
    ptr_deref_1985_store_0_req_0 <= cp_elements(511);
    cp_elements(512) <= ptr_deref_1985_store_0_ack_0;
    cp_elements(513) <= cp_elements(512);
    ptr_deref_1985_store_0_req_1 <= cp_elements(513);
    cp_elements(514) <= ptr_deref_1985_store_0_ack_1;
    cpelement_group_515 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(516) & cp_elements(517));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(515),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1990_inst_req_0 <= cp_elements(515);
    cp_elements(516) <= cp_elements(271);
    cp_elements(517) <= cp_elements(271);
    cp_elements(518) <= type_cast_1990_inst_ack_0;
    cpelement_group_519 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(395) & cp_elements(512) & cp_elements(518) & cp_elements(523));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(519),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1993_gather_scatter_req_0 <= cp_elements(519);
    cp_elements(520) <= cp_elements(395);
    ptr_deref_1993_base_resize_req_0 <= cp_elements(520);
    cp_elements(521) <= ptr_deref_1993_base_resize_ack_0;
    ptr_deref_1993_root_address_inst_req_0 <= cp_elements(521);
    cp_elements(522) <= ptr_deref_1993_root_address_inst_ack_0;
    ptr_deref_1993_addr_0_req_0 <= cp_elements(522);
    cp_elements(523) <= ptr_deref_1993_addr_0_ack_0;
    cp_elements(524) <= ptr_deref_1993_gather_scatter_ack_0;
    ptr_deref_1993_store_0_req_0 <= cp_elements(524);
    cp_elements(525) <= ptr_deref_1993_store_0_ack_0;
    ptr_deref_1993_store_0_req_1 <= cp_elements(525);
    cp_elements(526) <= ptr_deref_1993_store_0_ack_1;
    cpelement_group_527 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(412) & cp_elements(429) & cp_elements(446) & cp_elements(463) & cp_elements(480) & cp_elements(497) & cp_elements(514) & cp_elements(526));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(527),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(528) <= cp_elements(810);
    cpelement_group_529 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(530) & cp_elements(531));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(529),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2002_inst_req_0 <= cp_elements(529);
    cp_elements(530) <= cp_elements(528);
    cp_elements(531) <= cp_elements(528);
    cp_elements(532) <= binary_2002_inst_ack_0;
    binary_2002_inst_req_1 <= cp_elements(532);
    cp_elements(533) <= binary_2002_inst_ack_1;
    type_cast_1667_inst_req_0 <= cp_elements(533);
    cp_elements(534) <= cp_elements(129);
    cpelement_group_535 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(536) & cp_elements(537));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(535),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2010_inst_req_0 <= cp_elements(535);
    cp_elements(536) <= cp_elements(534);
    cp_elements(537) <= cp_elements(534);
    cp_elements(538) <= binary_2010_inst_ack_0;
    binary_2010_inst_req_1 <= cp_elements(538);
    cp_elements(539) <= binary_2010_inst_ack_1;
    cpelement_group_540 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(539) & cp_elements(541));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(540),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2014_inst_req_0 <= cp_elements(540);
    cp_elements(541) <= cp_elements(534);
    cp_elements(542) <= type_cast_2014_inst_ack_0;
    cp_elements(543) <= cp_elements(534);
    cpelement_group_544 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(543) & cp_elements(553));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(544),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2018_final_reg_req_0 <= cp_elements(544);
    cp_elements(545) <= cp_elements(534);
    array_obj_ref_2018_base_resize_req_0 <= cp_elements(545);
    cp_elements(546) <= cp_elements(534);
    array_obj_ref_2018_index_0_resize_req_0 <= cp_elements(546);
    cp_elements(547) <= array_obj_ref_2018_index_0_resize_ack_0;
    array_obj_ref_2018_index_0_rename_req_0 <= cp_elements(547);
    cp_elements(548) <= array_obj_ref_2018_index_0_rename_ack_0;
    array_obj_ref_2018_offset_inst_req_0 <= cp_elements(548);
    cp_elements(549) <= array_obj_ref_2018_offset_inst_ack_0;
    cp_elements(550) <= array_obj_ref_2018_base_resize_ack_0;
    cpelement_group_551 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(549) & cp_elements(550));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(551),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2018_root_address_inst_req_0 <= cp_elements(551);
    cp_elements(552) <= array_obj_ref_2018_root_address_inst_ack_0;
    array_obj_ref_2018_root_address_inst_req_1 <= cp_elements(552);
    cp_elements(553) <= array_obj_ref_2018_root_address_inst_ack_1;
    cp_elements(554) <= array_obj_ref_2018_final_reg_ack_0;
    cpelement_group_555 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(542) & cp_elements(554) & cp_elements(559));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(555),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2021_gather_scatter_req_0 <= cp_elements(555);
    cp_elements(556) <= cp_elements(554);
    ptr_deref_2021_base_resize_req_0 <= cp_elements(556);
    cp_elements(557) <= ptr_deref_2021_base_resize_ack_0;
    ptr_deref_2021_root_address_inst_req_0 <= cp_elements(557);
    cp_elements(558) <= ptr_deref_2021_root_address_inst_ack_0;
    ptr_deref_2021_addr_0_req_0 <= cp_elements(558);
    cp_elements(559) <= ptr_deref_2021_addr_0_ack_0;
    cp_elements(560) <= ptr_deref_2021_gather_scatter_ack_0;
    ptr_deref_2021_store_0_req_0 <= cp_elements(560);
    cp_elements(561) <= ptr_deref_2021_store_0_ack_0;
    cp_elements(562) <= cp_elements(561);
    ptr_deref_2021_store_0_req_1 <= cp_elements(562);
    cp_elements(563) <= ptr_deref_2021_store_0_ack_1;
    cpelement_group_564 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(565) & cp_elements(566));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(564),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2028_inst_req_0 <= cp_elements(564);
    cp_elements(565) <= cp_elements(534);
    cp_elements(566) <= cp_elements(534);
    cp_elements(567) <= binary_2028_inst_ack_0;
    binary_2028_inst_req_1 <= cp_elements(567);
    cp_elements(568) <= binary_2028_inst_ack_1;
    cpelement_group_569 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(568) & cp_elements(570));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(569),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2032_inst_req_0 <= cp_elements(569);
    cp_elements(570) <= cp_elements(534);
    cp_elements(571) <= type_cast_2032_inst_ack_0;
    cpelement_group_572 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(573) & cp_elements(574));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(572),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2038_inst_req_0 <= cp_elements(572);
    cp_elements(573) <= cp_elements(534);
    cp_elements(574) <= cp_elements(534);
    cp_elements(575) <= binary_2038_inst_ack_0;
    binary_2038_inst_req_1 <= cp_elements(575);
    cp_elements(576) <= binary_2038_inst_ack_1;
    array_obj_ref_2042_index_0_resize_req_0 <= cp_elements(576);
    cp_elements(577) <= cp_elements(534);
    cpelement_group_578 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(577) & cp_elements(586));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(578),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2042_final_reg_req_0 <= cp_elements(578);
    cp_elements(579) <= cp_elements(534);
    array_obj_ref_2042_base_resize_req_0 <= cp_elements(579);
    cp_elements(580) <= array_obj_ref_2042_index_0_resize_ack_0;
    array_obj_ref_2042_index_0_rename_req_0 <= cp_elements(580);
    cp_elements(581) <= array_obj_ref_2042_index_0_rename_ack_0;
    array_obj_ref_2042_offset_inst_req_0 <= cp_elements(581);
    cp_elements(582) <= array_obj_ref_2042_offset_inst_ack_0;
    cp_elements(583) <= array_obj_ref_2042_base_resize_ack_0;
    cpelement_group_584 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(582) & cp_elements(583));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(584),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2042_root_address_inst_req_0 <= cp_elements(584);
    cp_elements(585) <= array_obj_ref_2042_root_address_inst_ack_0;
    array_obj_ref_2042_root_address_inst_req_1 <= cp_elements(585);
    cp_elements(586) <= array_obj_ref_2042_root_address_inst_ack_1;
    cp_elements(587) <= array_obj_ref_2042_final_reg_ack_0;
    cpelement_group_588 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(561) & cp_elements(571) & cp_elements(587) & cp_elements(592));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(588),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2045_gather_scatter_req_0 <= cp_elements(588);
    cp_elements(589) <= cp_elements(587);
    ptr_deref_2045_base_resize_req_0 <= cp_elements(589);
    cp_elements(590) <= ptr_deref_2045_base_resize_ack_0;
    ptr_deref_2045_root_address_inst_req_0 <= cp_elements(590);
    cp_elements(591) <= ptr_deref_2045_root_address_inst_ack_0;
    ptr_deref_2045_addr_0_req_0 <= cp_elements(591);
    cp_elements(592) <= ptr_deref_2045_addr_0_ack_0;
    cp_elements(593) <= ptr_deref_2045_gather_scatter_ack_0;
    ptr_deref_2045_store_0_req_0 <= cp_elements(593);
    cp_elements(594) <= ptr_deref_2045_store_0_ack_0;
    cp_elements(595) <= cp_elements(594);
    ptr_deref_2045_store_0_req_1 <= cp_elements(595);
    cp_elements(596) <= ptr_deref_2045_store_0_ack_1;
    cpelement_group_597 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(598) & cp_elements(599));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(597),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2052_inst_req_0 <= cp_elements(597);
    cp_elements(598) <= cp_elements(534);
    cp_elements(599) <= cp_elements(534);
    cp_elements(600) <= binary_2052_inst_ack_0;
    binary_2052_inst_req_1 <= cp_elements(600);
    cp_elements(601) <= binary_2052_inst_ack_1;
    cpelement_group_602 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(601) & cp_elements(603));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(602),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2056_inst_req_0 <= cp_elements(602);
    cp_elements(603) <= cp_elements(534);
    cp_elements(604) <= type_cast_2056_inst_ack_0;
    cpelement_group_605 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(606) & cp_elements(607));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(605),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2062_inst_req_0 <= cp_elements(605);
    cp_elements(606) <= cp_elements(534);
    cp_elements(607) <= cp_elements(534);
    cp_elements(608) <= binary_2062_inst_ack_0;
    binary_2062_inst_req_1 <= cp_elements(608);
    cp_elements(609) <= binary_2062_inst_ack_1;
    array_obj_ref_2066_index_0_resize_req_0 <= cp_elements(609);
    cp_elements(610) <= cp_elements(534);
    cpelement_group_611 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(610) & cp_elements(619));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(611),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2066_final_reg_req_0 <= cp_elements(611);
    cp_elements(612) <= cp_elements(534);
    array_obj_ref_2066_base_resize_req_0 <= cp_elements(612);
    cp_elements(613) <= array_obj_ref_2066_index_0_resize_ack_0;
    array_obj_ref_2066_index_0_rename_req_0 <= cp_elements(613);
    cp_elements(614) <= array_obj_ref_2066_index_0_rename_ack_0;
    array_obj_ref_2066_offset_inst_req_0 <= cp_elements(614);
    cp_elements(615) <= array_obj_ref_2066_offset_inst_ack_0;
    cp_elements(616) <= array_obj_ref_2066_base_resize_ack_0;
    cpelement_group_617 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(615) & cp_elements(616));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(617),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2066_root_address_inst_req_0 <= cp_elements(617);
    cp_elements(618) <= array_obj_ref_2066_root_address_inst_ack_0;
    array_obj_ref_2066_root_address_inst_req_1 <= cp_elements(618);
    cp_elements(619) <= array_obj_ref_2066_root_address_inst_ack_1;
    cp_elements(620) <= array_obj_ref_2066_final_reg_ack_0;
    cpelement_group_621 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(594) & cp_elements(604) & cp_elements(620) & cp_elements(625));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2069_gather_scatter_req_0 <= cp_elements(621);
    cp_elements(622) <= cp_elements(620);
    ptr_deref_2069_base_resize_req_0 <= cp_elements(622);
    cp_elements(623) <= ptr_deref_2069_base_resize_ack_0;
    ptr_deref_2069_root_address_inst_req_0 <= cp_elements(623);
    cp_elements(624) <= ptr_deref_2069_root_address_inst_ack_0;
    ptr_deref_2069_addr_0_req_0 <= cp_elements(624);
    cp_elements(625) <= ptr_deref_2069_addr_0_ack_0;
    cp_elements(626) <= ptr_deref_2069_gather_scatter_ack_0;
    ptr_deref_2069_store_0_req_0 <= cp_elements(626);
    cp_elements(627) <= ptr_deref_2069_store_0_ack_0;
    cp_elements(628) <= cp_elements(627);
    ptr_deref_2069_store_0_req_1 <= cp_elements(628);
    cp_elements(629) <= ptr_deref_2069_store_0_ack_1;
    cpelement_group_630 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(631) & cp_elements(632));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(630),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2076_inst_req_0 <= cp_elements(630);
    cp_elements(631) <= cp_elements(534);
    cp_elements(632) <= cp_elements(534);
    cp_elements(633) <= binary_2076_inst_ack_0;
    binary_2076_inst_req_1 <= cp_elements(633);
    cp_elements(634) <= binary_2076_inst_ack_1;
    cpelement_group_635 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(634) & cp_elements(636));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(635),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2080_inst_req_0 <= cp_elements(635);
    cp_elements(636) <= cp_elements(534);
    cp_elements(637) <= type_cast_2080_inst_ack_0;
    cpelement_group_638 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(639) & cp_elements(640));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(638),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2086_inst_req_0 <= cp_elements(638);
    cp_elements(639) <= cp_elements(534);
    cp_elements(640) <= cp_elements(534);
    cp_elements(641) <= binary_2086_inst_ack_0;
    binary_2086_inst_req_1 <= cp_elements(641);
    cp_elements(642) <= binary_2086_inst_ack_1;
    array_obj_ref_2090_index_0_resize_req_0 <= cp_elements(642);
    cp_elements(643) <= cp_elements(534);
    cpelement_group_644 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(643) & cp_elements(652));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(644),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2090_final_reg_req_0 <= cp_elements(644);
    cp_elements(645) <= cp_elements(534);
    array_obj_ref_2090_base_resize_req_0 <= cp_elements(645);
    cp_elements(646) <= array_obj_ref_2090_index_0_resize_ack_0;
    array_obj_ref_2090_index_0_rename_req_0 <= cp_elements(646);
    cp_elements(647) <= array_obj_ref_2090_index_0_rename_ack_0;
    array_obj_ref_2090_offset_inst_req_0 <= cp_elements(647);
    cp_elements(648) <= array_obj_ref_2090_offset_inst_ack_0;
    cp_elements(649) <= array_obj_ref_2090_base_resize_ack_0;
    cpelement_group_650 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(648) & cp_elements(649));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(650),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2090_root_address_inst_req_0 <= cp_elements(650);
    cp_elements(651) <= array_obj_ref_2090_root_address_inst_ack_0;
    array_obj_ref_2090_root_address_inst_req_1 <= cp_elements(651);
    cp_elements(652) <= array_obj_ref_2090_root_address_inst_ack_1;
    cp_elements(653) <= array_obj_ref_2090_final_reg_ack_0;
    cpelement_group_654 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(627) & cp_elements(637) & cp_elements(653) & cp_elements(658));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(654),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2093_gather_scatter_req_0 <= cp_elements(654);
    cp_elements(655) <= cp_elements(653);
    ptr_deref_2093_base_resize_req_0 <= cp_elements(655);
    cp_elements(656) <= ptr_deref_2093_base_resize_ack_0;
    ptr_deref_2093_root_address_inst_req_0 <= cp_elements(656);
    cp_elements(657) <= ptr_deref_2093_root_address_inst_ack_0;
    ptr_deref_2093_addr_0_req_0 <= cp_elements(657);
    cp_elements(658) <= ptr_deref_2093_addr_0_ack_0;
    cp_elements(659) <= ptr_deref_2093_gather_scatter_ack_0;
    ptr_deref_2093_store_0_req_0 <= cp_elements(659);
    cp_elements(660) <= ptr_deref_2093_store_0_ack_0;
    cp_elements(661) <= cp_elements(660);
    ptr_deref_2093_store_0_req_1 <= cp_elements(661);
    cp_elements(662) <= ptr_deref_2093_store_0_ack_1;
    cpelement_group_663 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(664) & cp_elements(665));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(663),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2100_inst_req_0 <= cp_elements(663);
    cp_elements(664) <= cp_elements(534);
    cp_elements(665) <= cp_elements(534);
    cp_elements(666) <= binary_2100_inst_ack_0;
    binary_2100_inst_req_1 <= cp_elements(666);
    cp_elements(667) <= binary_2100_inst_ack_1;
    cpelement_group_668 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(667) & cp_elements(669));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(668),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2104_inst_req_0 <= cp_elements(668);
    cp_elements(669) <= cp_elements(534);
    cp_elements(670) <= type_cast_2104_inst_ack_0;
    cpelement_group_671 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(672) & cp_elements(673));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(671),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2110_inst_req_0 <= cp_elements(671);
    cp_elements(672) <= cp_elements(534);
    cp_elements(673) <= cp_elements(534);
    cp_elements(674) <= binary_2110_inst_ack_0;
    binary_2110_inst_req_1 <= cp_elements(674);
    cp_elements(675) <= binary_2110_inst_ack_1;
    array_obj_ref_2114_index_0_resize_req_0 <= cp_elements(675);
    cp_elements(676) <= cp_elements(534);
    cpelement_group_677 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(676) & cp_elements(685));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(677),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2114_final_reg_req_0 <= cp_elements(677);
    cp_elements(678) <= cp_elements(534);
    array_obj_ref_2114_base_resize_req_0 <= cp_elements(678);
    cp_elements(679) <= array_obj_ref_2114_index_0_resize_ack_0;
    array_obj_ref_2114_index_0_rename_req_0 <= cp_elements(679);
    cp_elements(680) <= array_obj_ref_2114_index_0_rename_ack_0;
    array_obj_ref_2114_offset_inst_req_0 <= cp_elements(680);
    cp_elements(681) <= array_obj_ref_2114_offset_inst_ack_0;
    cp_elements(682) <= array_obj_ref_2114_base_resize_ack_0;
    cpelement_group_683 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(681) & cp_elements(682));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(683),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2114_root_address_inst_req_0 <= cp_elements(683);
    cp_elements(684) <= array_obj_ref_2114_root_address_inst_ack_0;
    array_obj_ref_2114_root_address_inst_req_1 <= cp_elements(684);
    cp_elements(685) <= array_obj_ref_2114_root_address_inst_ack_1;
    cp_elements(686) <= array_obj_ref_2114_final_reg_ack_0;
    cpelement_group_687 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(660) & cp_elements(670) & cp_elements(686) & cp_elements(691));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(687),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2117_gather_scatter_req_0 <= cp_elements(687);
    cp_elements(688) <= cp_elements(686);
    ptr_deref_2117_base_resize_req_0 <= cp_elements(688);
    cp_elements(689) <= ptr_deref_2117_base_resize_ack_0;
    ptr_deref_2117_root_address_inst_req_0 <= cp_elements(689);
    cp_elements(690) <= ptr_deref_2117_root_address_inst_ack_0;
    ptr_deref_2117_addr_0_req_0 <= cp_elements(690);
    cp_elements(691) <= ptr_deref_2117_addr_0_ack_0;
    cp_elements(692) <= ptr_deref_2117_gather_scatter_ack_0;
    ptr_deref_2117_store_0_req_0 <= cp_elements(692);
    cp_elements(693) <= ptr_deref_2117_store_0_ack_0;
    cp_elements(694) <= cp_elements(693);
    ptr_deref_2117_store_0_req_1 <= cp_elements(694);
    cp_elements(695) <= ptr_deref_2117_store_0_ack_1;
    cpelement_group_696 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(697) & cp_elements(698));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(696),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2124_inst_req_0 <= cp_elements(696);
    cp_elements(697) <= cp_elements(534);
    cp_elements(698) <= cp_elements(534);
    cp_elements(699) <= binary_2124_inst_ack_0;
    binary_2124_inst_req_1 <= cp_elements(699);
    cp_elements(700) <= binary_2124_inst_ack_1;
    cpelement_group_701 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(700) & cp_elements(702));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(701),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2128_inst_req_0 <= cp_elements(701);
    cp_elements(702) <= cp_elements(534);
    cp_elements(703) <= type_cast_2128_inst_ack_0;
    cpelement_group_704 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(705) & cp_elements(706));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(704),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2134_inst_req_0 <= cp_elements(704);
    cp_elements(705) <= cp_elements(534);
    cp_elements(706) <= cp_elements(534);
    cp_elements(707) <= binary_2134_inst_ack_0;
    binary_2134_inst_req_1 <= cp_elements(707);
    cp_elements(708) <= binary_2134_inst_ack_1;
    array_obj_ref_2138_index_0_resize_req_0 <= cp_elements(708);
    cp_elements(709) <= cp_elements(534);
    cpelement_group_710 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(709) & cp_elements(718));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(710),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2138_final_reg_req_0 <= cp_elements(710);
    cp_elements(711) <= cp_elements(534);
    array_obj_ref_2138_base_resize_req_0 <= cp_elements(711);
    cp_elements(712) <= array_obj_ref_2138_index_0_resize_ack_0;
    array_obj_ref_2138_index_0_rename_req_0 <= cp_elements(712);
    cp_elements(713) <= array_obj_ref_2138_index_0_rename_ack_0;
    array_obj_ref_2138_offset_inst_req_0 <= cp_elements(713);
    cp_elements(714) <= array_obj_ref_2138_offset_inst_ack_0;
    cp_elements(715) <= array_obj_ref_2138_base_resize_ack_0;
    cpelement_group_716 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(714) & cp_elements(715));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(716),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2138_root_address_inst_req_0 <= cp_elements(716);
    cp_elements(717) <= array_obj_ref_2138_root_address_inst_ack_0;
    array_obj_ref_2138_root_address_inst_req_1 <= cp_elements(717);
    cp_elements(718) <= array_obj_ref_2138_root_address_inst_ack_1;
    cp_elements(719) <= array_obj_ref_2138_final_reg_ack_0;
    cpelement_group_720 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(693) & cp_elements(703) & cp_elements(719) & cp_elements(724));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(720),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2141_gather_scatter_req_0 <= cp_elements(720);
    cp_elements(721) <= cp_elements(719);
    ptr_deref_2141_base_resize_req_0 <= cp_elements(721);
    cp_elements(722) <= ptr_deref_2141_base_resize_ack_0;
    ptr_deref_2141_root_address_inst_req_0 <= cp_elements(722);
    cp_elements(723) <= ptr_deref_2141_root_address_inst_ack_0;
    ptr_deref_2141_addr_0_req_0 <= cp_elements(723);
    cp_elements(724) <= ptr_deref_2141_addr_0_ack_0;
    cp_elements(725) <= ptr_deref_2141_gather_scatter_ack_0;
    ptr_deref_2141_store_0_req_0 <= cp_elements(725);
    cp_elements(726) <= ptr_deref_2141_store_0_ack_0;
    cp_elements(727) <= cp_elements(726);
    ptr_deref_2141_store_0_req_1 <= cp_elements(727);
    cp_elements(728) <= ptr_deref_2141_store_0_ack_1;
    cpelement_group_729 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(730) & cp_elements(731));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(729),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2148_inst_req_0 <= cp_elements(729);
    cp_elements(730) <= cp_elements(534);
    cp_elements(731) <= cp_elements(534);
    cp_elements(732) <= binary_2148_inst_ack_0;
    binary_2148_inst_req_1 <= cp_elements(732);
    cp_elements(733) <= binary_2148_inst_ack_1;
    cpelement_group_734 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(733) & cp_elements(735));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(734),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2152_inst_req_0 <= cp_elements(734);
    cp_elements(735) <= cp_elements(534);
    cp_elements(736) <= type_cast_2152_inst_ack_0;
    cpelement_group_737 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(738) & cp_elements(739));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(737),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2158_inst_req_0 <= cp_elements(737);
    cp_elements(738) <= cp_elements(534);
    cp_elements(739) <= cp_elements(534);
    cp_elements(740) <= binary_2158_inst_ack_0;
    binary_2158_inst_req_1 <= cp_elements(740);
    cp_elements(741) <= binary_2158_inst_ack_1;
    array_obj_ref_2162_index_0_resize_req_0 <= cp_elements(741);
    cp_elements(742) <= cp_elements(534);
    cpelement_group_743 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(742) & cp_elements(751));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(743),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2162_final_reg_req_0 <= cp_elements(743);
    cp_elements(744) <= cp_elements(534);
    array_obj_ref_2162_base_resize_req_0 <= cp_elements(744);
    cp_elements(745) <= array_obj_ref_2162_index_0_resize_ack_0;
    array_obj_ref_2162_index_0_rename_req_0 <= cp_elements(745);
    cp_elements(746) <= array_obj_ref_2162_index_0_rename_ack_0;
    array_obj_ref_2162_offset_inst_req_0 <= cp_elements(746);
    cp_elements(747) <= array_obj_ref_2162_offset_inst_ack_0;
    cp_elements(748) <= array_obj_ref_2162_base_resize_ack_0;
    cpelement_group_749 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(747) & cp_elements(748));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(749),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2162_root_address_inst_req_0 <= cp_elements(749);
    cp_elements(750) <= array_obj_ref_2162_root_address_inst_ack_0;
    array_obj_ref_2162_root_address_inst_req_1 <= cp_elements(750);
    cp_elements(751) <= array_obj_ref_2162_root_address_inst_ack_1;
    cp_elements(752) <= array_obj_ref_2162_final_reg_ack_0;
    cpelement_group_753 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(726) & cp_elements(736) & cp_elements(752) & cp_elements(757));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(753),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2165_gather_scatter_req_0 <= cp_elements(753);
    cp_elements(754) <= cp_elements(752);
    ptr_deref_2165_base_resize_req_0 <= cp_elements(754);
    cp_elements(755) <= ptr_deref_2165_base_resize_ack_0;
    ptr_deref_2165_root_address_inst_req_0 <= cp_elements(755);
    cp_elements(756) <= ptr_deref_2165_root_address_inst_ack_0;
    ptr_deref_2165_addr_0_req_0 <= cp_elements(756);
    cp_elements(757) <= ptr_deref_2165_addr_0_ack_0;
    cp_elements(758) <= ptr_deref_2165_gather_scatter_ack_0;
    ptr_deref_2165_store_0_req_0 <= cp_elements(758);
    cp_elements(759) <= ptr_deref_2165_store_0_ack_0;
    cp_elements(760) <= cp_elements(759);
    ptr_deref_2165_store_0_req_1 <= cp_elements(760);
    cp_elements(761) <= ptr_deref_2165_store_0_ack_1;
    cpelement_group_762 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(763) & cp_elements(764));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(762),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2170_inst_req_0 <= cp_elements(762);
    cp_elements(763) <= cp_elements(534);
    cp_elements(764) <= cp_elements(534);
    cp_elements(765) <= type_cast_2170_inst_ack_0;
    cpelement_group_766 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(767) & cp_elements(768));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(766),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2176_inst_req_0 <= cp_elements(766);
    cp_elements(767) <= cp_elements(534);
    cp_elements(768) <= cp_elements(534);
    cp_elements(769) <= binary_2176_inst_ack_0;
    binary_2176_inst_req_1 <= cp_elements(769);
    cp_elements(770) <= binary_2176_inst_ack_1;
    array_obj_ref_2180_index_0_resize_req_0 <= cp_elements(770);
    cp_elements(771) <= cp_elements(534);
    cpelement_group_772 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(771) & cp_elements(780));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(772),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2180_final_reg_req_0 <= cp_elements(772);
    cp_elements(773) <= cp_elements(534);
    array_obj_ref_2180_base_resize_req_0 <= cp_elements(773);
    cp_elements(774) <= array_obj_ref_2180_index_0_resize_ack_0;
    array_obj_ref_2180_index_0_rename_req_0 <= cp_elements(774);
    cp_elements(775) <= array_obj_ref_2180_index_0_rename_ack_0;
    array_obj_ref_2180_offset_inst_req_0 <= cp_elements(775);
    cp_elements(776) <= array_obj_ref_2180_offset_inst_ack_0;
    cp_elements(777) <= array_obj_ref_2180_base_resize_ack_0;
    cpelement_group_778 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(776) & cp_elements(777));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(778),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2180_root_address_inst_req_0 <= cp_elements(778);
    cp_elements(779) <= array_obj_ref_2180_root_address_inst_ack_0;
    array_obj_ref_2180_root_address_inst_req_1 <= cp_elements(779);
    cp_elements(780) <= array_obj_ref_2180_root_address_inst_ack_1;
    cp_elements(781) <= array_obj_ref_2180_final_reg_ack_0;
    cpelement_group_782 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(759) & cp_elements(765) & cp_elements(781) & cp_elements(786));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(782),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2183_gather_scatter_req_0 <= cp_elements(782);
    cp_elements(783) <= cp_elements(781);
    ptr_deref_2183_base_resize_req_0 <= cp_elements(783);
    cp_elements(784) <= ptr_deref_2183_base_resize_ack_0;
    ptr_deref_2183_root_address_inst_req_0 <= cp_elements(784);
    cp_elements(785) <= ptr_deref_2183_root_address_inst_ack_0;
    ptr_deref_2183_addr_0_req_0 <= cp_elements(785);
    cp_elements(786) <= ptr_deref_2183_addr_0_ack_0;
    cp_elements(787) <= ptr_deref_2183_gather_scatter_ack_0;
    ptr_deref_2183_store_0_req_0 <= cp_elements(787);
    cp_elements(788) <= ptr_deref_2183_store_0_ack_0;
    ptr_deref_2183_store_0_req_1 <= cp_elements(788);
    cp_elements(789) <= ptr_deref_2183_store_0_ack_1;
    cpelement_group_790 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(791) & cp_elements(792));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(790),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2190_inst_req_0 <= cp_elements(790);
    cp_elements(791) <= cp_elements(534);
    cp_elements(792) <= cp_elements(534);
    cp_elements(793) <= binary_2190_inst_ack_0;
    binary_2190_inst_req_1 <= cp_elements(793);
    cp_elements(794) <= binary_2190_inst_ack_1;
    cpelement_group_795 : Block -- 
      signal predecessors: BooleanArray(8 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(563) & cp_elements(596) & cp_elements(629) & cp_elements(662) & cp_elements(695) & cp_elements(728) & cp_elements(761) & cp_elements(789) & cp_elements(794));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(795),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(796) <= simple_obj_ref_2198_inst_ack_0;
    simple_obj_ref_2207_inst_req_0 <= cp_elements(796);
    cp_elements(797) <= simple_obj_ref_2207_inst_ack_0;
    simple_obj_ref_2216_inst_req_0 <= cp_elements(797);
    cp_elements(798) <= simple_obj_ref_2216_inst_ack_0;
    cp_elements(799) <= OrReduce(cp_elements(18) & cp_elements(35) & cp_elements(798));
    cp_elements(800) <= cp_elements(799);
    simple_obj_ref_1575_inst_req_0 <= cp_elements(800);
    cp_elements(801) <= false;
    cp_elements(802) <= cp_elements(801);
    cp_elements(803) <= type_cast_1667_inst_ack_0;
    phi_stmt_1661_req_1 <= cp_elements(803);
    cp_elements(804) <= OrReduce(cp_elements(4) & cp_elements(803));
    cp_elements(805) <= cp_elements(804);
    cp_elements(806) <= phi_stmt_1661_ack_0;
    cp_elements(807) <= false;
    cp_elements(808) <= cp_elements(807);
    cp_elements(809) <= OrReduce(cp_elements(6) & cp_elements(7));
    cp_elements(810) <= cp_elements(809);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1623_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1623_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1623_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1628_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1628_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1628_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1633_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1633_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1633_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1638_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1638_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1638_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1647_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1647_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1647_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1652_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1652_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1652_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1657_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1657_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1657_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1860_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1860_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1860_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1860_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1864_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1864_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1864_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1864_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1872_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1872_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1872_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1872_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1876_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1876_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1876_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1876_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1880_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1880_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1880_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1880_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1884_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1884_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1884_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1884_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2042_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2042_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2042_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2042_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2066_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2066_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2066_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2066_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2090_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2090_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2090_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2090_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2114_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2114_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2114_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2114_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2138_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2138_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2138_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2138_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2162_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2162_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2162_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2162_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2180_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2180_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2180_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2180_root_address : std_logic_vector(10 downto 0);
    signal expr_1699_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1699_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_1702_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1702_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal iNsTr_0_1552 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1661 : std_logic_vector(31 downto 0);
    signal iNsTr_11_1680 : std_logic_vector(31 downto 0);
    signal iNsTr_12_1689 : std_logic_vector(31 downto 0);
    signal iNsTr_22_2197 : std_logic_vector(31 downto 0);
    signal iNsTr_24_2206 : std_logic_vector(31 downto 0);
    signal iNsTr_26_2215 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1563 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1574 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1584 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1606 : std_logic_vector(31 downto 0);
    signal ptr_deref_1554_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1554_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1554_word_address_0 : std_logic_vector(3 downto 0);
    signal ptr_deref_1719_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1719_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1719_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1719_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1719_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1719_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1733_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1733_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1733_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1733_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1733_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1733_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1747_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1747_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1747_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1747_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1747_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1747_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1761_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1761_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1761_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1761_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1761_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1761_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1775_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1775_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1775_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1775_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1775_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1775_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1789_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1789_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1789_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1789_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1789_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1789_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1803_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1803_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1803_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1803_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1803_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1803_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1811_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1811_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1811_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1811_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1811_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1811_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1901_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1901_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1901_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1901_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1901_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1901_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1915_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1915_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1915_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1915_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1915_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1915_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1929_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1929_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1929_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1929_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1929_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1929_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1943_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1943_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1943_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1943_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1943_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1943_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1957_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1957_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1957_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1957_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1957_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1957_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1971_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1971_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1971_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1971_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1971_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1971_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1985_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1985_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1985_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1985_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1985_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1985_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1993_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1993_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1993_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1993_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1993_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1993_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2021_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2021_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2021_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2021_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2021_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2021_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2045_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2045_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2045_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2045_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2045_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2045_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2069_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2069_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2069_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2069_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2069_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2069_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2093_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2093_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2093_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2093_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2093_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2093_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2117_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2117_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2117_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2117_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2117_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2117_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2141_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2141_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2141_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2141_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2141_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2141_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2165_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2165_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2183_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2183_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_word_offset_0 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1859_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1859_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1863_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1863_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1867_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1867_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1871_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1871_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1875_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1875_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1879_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1879_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1883_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1883_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1887_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1887_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2017_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2017_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2041_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2041_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2065_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2065_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2089_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2089_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2113_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2113_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2137_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2137_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2161_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2161_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2179_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2179_scaled : std_logic_vector(10 downto 0);
    signal tmp100_1877 : std_logic_vector(31 downto 0);
    signal tmp103_1881 : std_logic_vector(31 downto 0);
    signal tmp106_1885 : std_logic_vector(31 downto 0);
    signal tmp109_1889 : std_logic_vector(31 downto 0);
    signal tmp10_1755 : std_logic_vector(63 downto 0);
    signal tmp113_2019 : std_logic_vector(31 downto 0);
    signal tmp115_2039 : std_logic_vector(31 downto 0);
    signal tmp116_2043 : std_logic_vector(31 downto 0);
    signal tmp118_2063 : std_logic_vector(31 downto 0);
    signal tmp119_2067 : std_logic_vector(31 downto 0);
    signal tmp11_1759 : std_logic_vector(7 downto 0);
    signal tmp121_2087 : std_logic_vector(31 downto 0);
    signal tmp122_2091 : std_logic_vector(31 downto 0);
    signal tmp124_2111 : std_logic_vector(31 downto 0);
    signal tmp125_2115 : std_logic_vector(31 downto 0);
    signal tmp127_2135 : std_logic_vector(31 downto 0);
    signal tmp128_2139 : std_logic_vector(31 downto 0);
    signal tmp130_2159 : std_logic_vector(31 downto 0);
    signal tmp131_2163 : std_logic_vector(31 downto 0);
    signal tmp133_2177 : std_logic_vector(31 downto 0);
    signal tmp134_2181 : std_logic_vector(31 downto 0);
    signal tmp135_2191 : std_logic_vector(31 downto 0);
    signal tmp137_1674 : std_logic_vector(31 downto 0);
    signal tmp138145_1857 : std_logic_vector(31 downto 0);
    signal tmp139146_1851 : std_logic_vector(31 downto 0);
    signal tmp13_1769 : std_logic_vector(63 downto 0);
    signal tmp140147_1845 : std_logic_vector(31 downto 0);
    signal tmp141148_1839 : std_logic_vector(31 downto 0);
    signal tmp142149_1833 : std_logic_vector(31 downto 0);
    signal tmp143150_1827 : std_logic_vector(31 downto 0);
    signal tmp144151_1821 : std_logic_vector(31 downto 0);
    signal tmp14_1773 : std_logic_vector(7 downto 0);
    signal tmp16_1783 : std_logic_vector(63 downto 0);
    signal tmp17_1787 : std_logic_vector(7 downto 0);
    signal tmp19_1797 : std_logic_vector(63 downto 0);
    signal tmp1_1713 : std_logic_vector(63 downto 0);
    signal tmp20_1801 : std_logic_vector(7 downto 0);
    signal tmp22_1809 : std_logic_vector(7 downto 0);
    signal tmp24_1895 : std_logic_vector(63 downto 0);
    signal tmp25_1899 : std_logic_vector(7 downto 0);
    signal tmp27_1909 : std_logic_vector(63 downto 0);
    signal tmp28_1913 : std_logic_vector(7 downto 0);
    signal tmp2_1717 : std_logic_vector(7 downto 0);
    signal tmp2x_xi_1593 : std_logic_vector(0 downto 0);
    signal tmp30_1923 : std_logic_vector(63 downto 0);
    signal tmp31_1927 : std_logic_vector(7 downto 0);
    signal tmp33_1937 : std_logic_vector(63 downto 0);
    signal tmp34_1941 : std_logic_vector(7 downto 0);
    signal tmp36_1951 : std_logic_vector(63 downto 0);
    signal tmp37_1955 : std_logic_vector(7 downto 0);
    signal tmp39_1965 : std_logic_vector(63 downto 0);
    signal tmp40_1969 : std_logic_vector(7 downto 0);
    signal tmp42_1979 : std_logic_vector(63 downto 0);
    signal tmp43_1983 : std_logic_vector(7 downto 0);
    signal tmp45_1991 : std_logic_vector(7 downto 0);
    signal tmp47_2011 : std_logic_vector(63 downto 0);
    signal tmp48_2015 : std_logic_vector(7 downto 0);
    signal tmp4_1727 : std_logic_vector(63 downto 0);
    signal tmp4x_xi_1609 : std_logic_vector(31 downto 0);
    signal tmp50_2029 : std_logic_vector(63 downto 0);
    signal tmp51_2033 : std_logic_vector(7 downto 0);
    signal tmp53_2053 : std_logic_vector(63 downto 0);
    signal tmp54_2057 : std_logic_vector(7 downto 0);
    signal tmp56_2077 : std_logic_vector(63 downto 0);
    signal tmp57_2081 : std_logic_vector(7 downto 0);
    signal tmp59_2101 : std_logic_vector(63 downto 0);
    signal tmp5_1731 : std_logic_vector(7 downto 0);
    signal tmp5x_xi_1614 : std_logic_vector(31 downto 0);
    signal tmp60_2105 : std_logic_vector(7 downto 0);
    signal tmp62_2125 : std_logic_vector(63 downto 0);
    signal tmp63_2129 : std_logic_vector(7 downto 0);
    signal tmp65_2149 : std_logic_vector(63 downto 0);
    signal tmp66_2153 : std_logic_vector(7 downto 0);
    signal tmp68_2171 : std_logic_vector(7 downto 0);
    signal tmp71_1619 : std_logic_vector(31 downto 0);
    signal tmp73_1683 : std_logic_vector(63 downto 0);
    signal tmp74_1692 : std_logic_vector(7 downto 0);
    signal tmp75_1696 : std_logic_vector(31 downto 0);
    signal tmp77_1624 : std_logic_vector(31 downto 0);
    signal tmp78_1629 : std_logic_vector(31 downto 0);
    signal tmp79_1634 : std_logic_vector(31 downto 0);
    signal tmp7_1741 : std_logic_vector(63 downto 0);
    signal tmp80_1639 : std_logic_vector(31 downto 0);
    signal tmp81_1643 : std_logic_vector(31 downto 0);
    signal tmp82_1648 : std_logic_vector(31 downto 0);
    signal tmp83_1653 : std_logic_vector(31 downto 0);
    signal tmp84_1658 : std_logic_vector(31 downto 0);
    signal tmp88_1861 : std_logic_vector(31 downto 0);
    signal tmp8_1745 : std_logic_vector(7 downto 0);
    signal tmp91_1865 : std_logic_vector(31 downto 0);
    signal tmp94_1869 : std_logic_vector(31 downto 0);
    signal tmp97_1873 : std_logic_vector(31 downto 0);
    signal tmp_1566 : std_logic_vector(7 downto 0);
    signal tmpx_xi_1587 : std_logic_vector(7 downto 0);
    signal type_cast_1556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1577_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1591_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1665_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1667_wire : std_logic_vector(31 downto 0);
    signal type_cast_1672_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1711_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1725_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1739_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1753_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1767_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1781_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1795_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1819_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1825_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1831_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1837_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1843_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1849_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1855_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1893_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1907_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1921_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1949_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1963_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1977_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2001_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2009_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2027_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2037_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2051_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2061_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2075_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2085_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2099_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2109_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2123_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2147_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2157_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2175_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2189_wire_constant : std_logic_vector(31 downto 0);
    signal wordx_x0x_xbe_2003 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1623_final_offset <= "00000000001";
    array_obj_ref_1628_final_offset <= "00000000010";
    array_obj_ref_1633_final_offset <= "00000000011";
    array_obj_ref_1638_final_offset <= "00000000100";
    array_obj_ref_1647_final_offset <= "00000000101";
    array_obj_ref_1652_final_offset <= "00000000110";
    array_obj_ref_1657_final_offset <= "00000000111";
    array_obj_ref_1860_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1864_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1868_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1872_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1876_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1880_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1884_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1888_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2018_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2042_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2066_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2090_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2114_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2138_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2162_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2180_offset_scale_factor_0 <= "00000000001";
    expr_1699_wire_constant <= "00000000000000000000000011111111";
    expr_1702_wire_constant <= "00000000000000000000000000000000";
    iNsTr_0_1552 <= "00000000000000000000000000000000";
    iNsTr_11_1680 <= "00000000000000000000000000000000";
    iNsTr_12_1689 <= "00000000000000000000000000000000";
    iNsTr_22_2197 <= "00000000000000000000000000000000";
    iNsTr_24_2206 <= "00000000000000000000000000000000";
    iNsTr_26_2215 <= "00000000000000000000000000000000";
    iNsTr_2_1563 <= "00000000000000000000000000000000";
    iNsTr_4_1574 <= "00000000000000000000000000000000";
    iNsTr_6_1584 <= "00000000000000000000000000000000";
    iNsTr_8_1606 <= "00000000000000000000000000000000";
    ptr_deref_1554_word_address_0 <= "0000";
    ptr_deref_1719_word_offset_0 <= "00000000000";
    ptr_deref_1733_word_offset_0 <= "00000000000";
    ptr_deref_1747_word_offset_0 <= "00000000000";
    ptr_deref_1761_word_offset_0 <= "00000000000";
    ptr_deref_1775_word_offset_0 <= "00000000000";
    ptr_deref_1789_word_offset_0 <= "00000000000";
    ptr_deref_1803_word_offset_0 <= "00000000000";
    ptr_deref_1811_word_offset_0 <= "00000000000";
    ptr_deref_1901_word_offset_0 <= "00000000000";
    ptr_deref_1915_word_offset_0 <= "00000000000";
    ptr_deref_1929_word_offset_0 <= "00000000000";
    ptr_deref_1943_word_offset_0 <= "00000000000";
    ptr_deref_1957_word_offset_0 <= "00000000000";
    ptr_deref_1971_word_offset_0 <= "00000000000";
    ptr_deref_1985_word_offset_0 <= "00000000000";
    ptr_deref_1993_word_offset_0 <= "00000000000";
    ptr_deref_2021_word_offset_0 <= "00000000000";
    ptr_deref_2045_word_offset_0 <= "00000000000";
    ptr_deref_2069_word_offset_0 <= "00000000000";
    ptr_deref_2093_word_offset_0 <= "00000000000";
    ptr_deref_2117_word_offset_0 <= "00000000000";
    ptr_deref_2141_word_offset_0 <= "00000000000";
    ptr_deref_2165_word_offset_0 <= "00000000000";
    ptr_deref_2183_word_offset_0 <= "00000000000";
    type_cast_1556_wire_constant <= "00000001";
    type_cast_1577_wire_constant <= "00000010";
    type_cast_1591_wire_constant <= "00000011";
    type_cast_1665_wire_constant <= "00000000000000000000000000000000";
    type_cast_1672_wire_constant <= "00000000000000000000000000000011";
    type_cast_1711_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1725_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1739_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1753_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1767_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1781_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1795_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1819_wire_constant <= "00000000000000000000000000000001";
    type_cast_1825_wire_constant <= "00000000000000000000000000000010";
    type_cast_1831_wire_constant <= "00000000000000000000000000000011";
    type_cast_1837_wire_constant <= "00000000000000000000000000000100";
    type_cast_1843_wire_constant <= "00000000000000000000000000000101";
    type_cast_1849_wire_constant <= "00000000000000000000000000000110";
    type_cast_1855_wire_constant <= "00000000000000000000000000000111";
    type_cast_1893_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1907_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1921_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1935_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1949_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1963_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1977_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2001_wire_constant <= "00000000000000000000000000000001";
    type_cast_2009_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2027_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2037_wire_constant <= "00000000000000000000000000000001";
    type_cast_2051_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2061_wire_constant <= "00000000000000000000000000000010";
    type_cast_2075_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2085_wire_constant <= "00000000000000000000000000000011";
    type_cast_2099_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2109_wire_constant <= "00000000000000000000000000000100";
    type_cast_2123_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2133_wire_constant <= "00000000000000000000000000000101";
    type_cast_2147_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2157_wire_constant <= "00000000000000000000000000000110";
    type_cast_2175_wire_constant <= "00000000000000000000000000000111";
    type_cast_2189_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1661: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1665_wire_constant & type_cast_1667_wire;
      req <= phi_stmt_1661_req_0 & phi_stmt_1661_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1661_ack_0,
          idata => idata,
          odata => iNsTr_10_1661,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1661
    array_obj_ref_1623_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1623_resized_base_address, req => array_obj_ref_1623_base_resize_req_0, ack => array_obj_ref_1623_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1623_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1623_root_address, dout => tmp77_1624, req => array_obj_ref_1623_final_reg_req_0, ack => array_obj_ref_1623_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1628_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1628_resized_base_address, req => array_obj_ref_1628_base_resize_req_0, ack => array_obj_ref_1628_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1628_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1628_root_address, dout => tmp78_1629, req => array_obj_ref_1628_final_reg_req_0, ack => array_obj_ref_1628_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1633_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1633_resized_base_address, req => array_obj_ref_1633_base_resize_req_0, ack => array_obj_ref_1633_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1633_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1633_root_address, dout => tmp79_1634, req => array_obj_ref_1633_final_reg_req_0, ack => array_obj_ref_1633_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1638_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp5x_xi_1614, dout => array_obj_ref_1638_resized_base_address, req => array_obj_ref_1638_base_resize_req_0, ack => array_obj_ref_1638_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1638_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1638_root_address, dout => tmp80_1639, req => array_obj_ref_1638_final_reg_req_0, ack => array_obj_ref_1638_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1647_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1647_resized_base_address, req => array_obj_ref_1647_base_resize_req_0, ack => array_obj_ref_1647_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1647_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1647_root_address, dout => tmp82_1648, req => array_obj_ref_1647_final_reg_req_0, ack => array_obj_ref_1647_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1652_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1652_resized_base_address, req => array_obj_ref_1652_base_resize_req_0, ack => array_obj_ref_1652_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1652_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1652_root_address, dout => tmp83_1653, req => array_obj_ref_1652_final_reg_req_0, ack => array_obj_ref_1652_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1657_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1657_resized_base_address, req => array_obj_ref_1657_base_resize_req_0, ack => array_obj_ref_1657_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1657_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1657_root_address, dout => tmp84_1658, req => array_obj_ref_1657_final_reg_req_0, ack => array_obj_ref_1657_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1860_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1860_resized_base_address, req => array_obj_ref_1860_base_resize_req_0, ack => array_obj_ref_1860_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1860_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1860_root_address, dout => tmp88_1861, req => array_obj_ref_1860_final_reg_req_0, ack => array_obj_ref_1860_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1860_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp137_1674, dout => simple_obj_ref_1859_resized, req => array_obj_ref_1860_index_0_resize_req_0, ack => array_obj_ref_1860_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1860_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1859_scaled, dout => array_obj_ref_1860_final_offset, req => array_obj_ref_1860_offset_inst_req_0, ack => array_obj_ref_1860_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1864_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1864_resized_base_address, req => array_obj_ref_1864_base_resize_req_0, ack => array_obj_ref_1864_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1864_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1864_root_address, dout => tmp91_1865, req => array_obj_ref_1864_final_reg_req_0, ack => array_obj_ref_1864_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1864_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp144151_1821, dout => simple_obj_ref_1863_resized, req => array_obj_ref_1864_index_0_resize_req_0, ack => array_obj_ref_1864_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1864_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1863_scaled, dout => array_obj_ref_1864_final_offset, req => array_obj_ref_1864_offset_inst_req_0, ack => array_obj_ref_1864_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1868_resized_base_address, req => array_obj_ref_1868_base_resize_req_0, ack => array_obj_ref_1868_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1868_root_address, dout => tmp94_1869, req => array_obj_ref_1868_final_reg_req_0, ack => array_obj_ref_1868_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp143150_1827, dout => simple_obj_ref_1867_resized, req => array_obj_ref_1868_index_0_resize_req_0, ack => array_obj_ref_1868_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1867_scaled, dout => array_obj_ref_1868_final_offset, req => array_obj_ref_1868_offset_inst_req_0, ack => array_obj_ref_1868_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1872_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1872_resized_base_address, req => array_obj_ref_1872_base_resize_req_0, ack => array_obj_ref_1872_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1872_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1872_root_address, dout => tmp97_1873, req => array_obj_ref_1872_final_reg_req_0, ack => array_obj_ref_1872_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1872_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp142149_1833, dout => simple_obj_ref_1871_resized, req => array_obj_ref_1872_index_0_resize_req_0, ack => array_obj_ref_1872_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1872_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1871_scaled, dout => array_obj_ref_1872_final_offset, req => array_obj_ref_1872_offset_inst_req_0, ack => array_obj_ref_1872_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1876_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1876_resized_base_address, req => array_obj_ref_1876_base_resize_req_0, ack => array_obj_ref_1876_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1876_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1876_root_address, dout => tmp100_1877, req => array_obj_ref_1876_final_reg_req_0, ack => array_obj_ref_1876_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1876_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp141148_1839, dout => simple_obj_ref_1875_resized, req => array_obj_ref_1876_index_0_resize_req_0, ack => array_obj_ref_1876_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1876_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1875_scaled, dout => array_obj_ref_1876_final_offset, req => array_obj_ref_1876_offset_inst_req_0, ack => array_obj_ref_1876_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1880_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1880_resized_base_address, req => array_obj_ref_1880_base_resize_req_0, ack => array_obj_ref_1880_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1880_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1880_root_address, dout => tmp103_1881, req => array_obj_ref_1880_final_reg_req_0, ack => array_obj_ref_1880_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1880_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp140147_1845, dout => simple_obj_ref_1879_resized, req => array_obj_ref_1880_index_0_resize_req_0, ack => array_obj_ref_1880_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1880_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1879_scaled, dout => array_obj_ref_1880_final_offset, req => array_obj_ref_1880_offset_inst_req_0, ack => array_obj_ref_1880_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1884_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1884_resized_base_address, req => array_obj_ref_1884_base_resize_req_0, ack => array_obj_ref_1884_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1884_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1884_root_address, dout => tmp106_1885, req => array_obj_ref_1884_final_reg_req_0, ack => array_obj_ref_1884_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1884_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp139146_1851, dout => simple_obj_ref_1883_resized, req => array_obj_ref_1884_index_0_resize_req_0, ack => array_obj_ref_1884_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1884_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1883_scaled, dout => array_obj_ref_1884_final_offset, req => array_obj_ref_1884_offset_inst_req_0, ack => array_obj_ref_1884_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_1888_resized_base_address, req => array_obj_ref_1888_base_resize_req_0, ack => array_obj_ref_1888_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1888_root_address, dout => tmp109_1889, req => array_obj_ref_1888_final_reg_req_0, ack => array_obj_ref_1888_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp138145_1857, dout => simple_obj_ref_1887_resized, req => array_obj_ref_1888_index_0_resize_req_0, ack => array_obj_ref_1888_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1887_scaled, dout => array_obj_ref_1888_final_offset, req => array_obj_ref_1888_offset_inst_req_0, ack => array_obj_ref_1888_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2018_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2018_resized_base_address, req => array_obj_ref_2018_base_resize_req_0, ack => array_obj_ref_2018_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2018_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2018_root_address, dout => tmp113_2019, req => array_obj_ref_2018_final_reg_req_0, ack => array_obj_ref_2018_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2018_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp137_1674, dout => simple_obj_ref_2017_resized, req => array_obj_ref_2018_index_0_resize_req_0, ack => array_obj_ref_2018_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2018_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2017_scaled, dout => array_obj_ref_2018_final_offset, req => array_obj_ref_2018_offset_inst_req_0, ack => array_obj_ref_2018_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2042_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2042_resized_base_address, req => array_obj_ref_2042_base_resize_req_0, ack => array_obj_ref_2042_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2042_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2042_root_address, dout => tmp116_2043, req => array_obj_ref_2042_final_reg_req_0, ack => array_obj_ref_2042_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2042_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp115_2039, dout => simple_obj_ref_2041_resized, req => array_obj_ref_2042_index_0_resize_req_0, ack => array_obj_ref_2042_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2042_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2041_scaled, dout => array_obj_ref_2042_final_offset, req => array_obj_ref_2042_offset_inst_req_0, ack => array_obj_ref_2042_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2066_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2066_resized_base_address, req => array_obj_ref_2066_base_resize_req_0, ack => array_obj_ref_2066_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2066_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2066_root_address, dout => tmp119_2067, req => array_obj_ref_2066_final_reg_req_0, ack => array_obj_ref_2066_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2066_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp118_2063, dout => simple_obj_ref_2065_resized, req => array_obj_ref_2066_index_0_resize_req_0, ack => array_obj_ref_2066_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2066_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2065_scaled, dout => array_obj_ref_2066_final_offset, req => array_obj_ref_2066_offset_inst_req_0, ack => array_obj_ref_2066_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2090_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2090_resized_base_address, req => array_obj_ref_2090_base_resize_req_0, ack => array_obj_ref_2090_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2090_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2090_root_address, dout => tmp122_2091, req => array_obj_ref_2090_final_reg_req_0, ack => array_obj_ref_2090_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2090_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp121_2087, dout => simple_obj_ref_2089_resized, req => array_obj_ref_2090_index_0_resize_req_0, ack => array_obj_ref_2090_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2090_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2089_scaled, dout => array_obj_ref_2090_final_offset, req => array_obj_ref_2090_offset_inst_req_0, ack => array_obj_ref_2090_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2114_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2114_resized_base_address, req => array_obj_ref_2114_base_resize_req_0, ack => array_obj_ref_2114_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2114_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2114_root_address, dout => tmp125_2115, req => array_obj_ref_2114_final_reg_req_0, ack => array_obj_ref_2114_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2114_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_2111, dout => simple_obj_ref_2113_resized, req => array_obj_ref_2114_index_0_resize_req_0, ack => array_obj_ref_2114_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2114_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2113_scaled, dout => array_obj_ref_2114_final_offset, req => array_obj_ref_2114_offset_inst_req_0, ack => array_obj_ref_2114_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2138_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2138_resized_base_address, req => array_obj_ref_2138_base_resize_req_0, ack => array_obj_ref_2138_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2138_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2138_root_address, dout => tmp128_2139, req => array_obj_ref_2138_final_reg_req_0, ack => array_obj_ref_2138_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2138_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp127_2135, dout => simple_obj_ref_2137_resized, req => array_obj_ref_2138_index_0_resize_req_0, ack => array_obj_ref_2138_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2138_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2137_scaled, dout => array_obj_ref_2138_final_offset, req => array_obj_ref_2138_offset_inst_req_0, ack => array_obj_ref_2138_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2162_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2162_resized_base_address, req => array_obj_ref_2162_base_resize_req_0, ack => array_obj_ref_2162_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2162_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2162_root_address, dout => tmp131_2163, req => array_obj_ref_2162_final_reg_req_0, ack => array_obj_ref_2162_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2162_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp130_2159, dout => simple_obj_ref_2161_resized, req => array_obj_ref_2162_index_0_resize_req_0, ack => array_obj_ref_2162_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2162_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2161_scaled, dout => array_obj_ref_2162_final_offset, req => array_obj_ref_2162_offset_inst_req_0, ack => array_obj_ref_2162_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2180_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => array_obj_ref_2180_resized_base_address, req => array_obj_ref_2180_base_resize_req_0, ack => array_obj_ref_2180_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2180_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2180_root_address, dout => tmp134_2181, req => array_obj_ref_2180_final_reg_req_0, ack => array_obj_ref_2180_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2180_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp133_2177, dout => simple_obj_ref_2179_resized, req => array_obj_ref_2180_index_0_resize_req_0, ack => array_obj_ref_2180_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2180_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2179_scaled, dout => array_obj_ref_2180_final_offset, req => array_obj_ref_2180_offset_inst_req_0, ack => array_obj_ref_2180_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1719_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp71_1619, dout => ptr_deref_1719_resized_base_address, req => ptr_deref_1719_base_resize_req_0, ack => ptr_deref_1719_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1733_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp77_1624, dout => ptr_deref_1733_resized_base_address, req => ptr_deref_1733_base_resize_req_0, ack => ptr_deref_1733_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1747_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp78_1629, dout => ptr_deref_1747_resized_base_address, req => ptr_deref_1747_base_resize_req_0, ack => ptr_deref_1747_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1761_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp79_1634, dout => ptr_deref_1761_resized_base_address, req => ptr_deref_1761_base_resize_req_0, ack => ptr_deref_1761_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1775_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp81_1643, dout => ptr_deref_1775_resized_base_address, req => ptr_deref_1775_base_resize_req_0, ack => ptr_deref_1775_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1789_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp82_1648, dout => ptr_deref_1789_resized_base_address, req => ptr_deref_1789_base_resize_req_0, ack => ptr_deref_1789_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1803_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp83_1653, dout => ptr_deref_1803_resized_base_address, req => ptr_deref_1803_base_resize_req_0, ack => ptr_deref_1803_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1811_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp84_1658, dout => ptr_deref_1811_resized_base_address, req => ptr_deref_1811_base_resize_req_0, ack => ptr_deref_1811_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1901_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp88_1861, dout => ptr_deref_1901_resized_base_address, req => ptr_deref_1901_base_resize_req_0, ack => ptr_deref_1901_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1915_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp91_1865, dout => ptr_deref_1915_resized_base_address, req => ptr_deref_1915_base_resize_req_0, ack => ptr_deref_1915_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1929_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp94_1869, dout => ptr_deref_1929_resized_base_address, req => ptr_deref_1929_base_resize_req_0, ack => ptr_deref_1929_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1943_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp97_1873, dout => ptr_deref_1943_resized_base_address, req => ptr_deref_1943_base_resize_req_0, ack => ptr_deref_1943_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1957_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp100_1877, dout => ptr_deref_1957_resized_base_address, req => ptr_deref_1957_base_resize_req_0, ack => ptr_deref_1957_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1971_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp103_1881, dout => ptr_deref_1971_resized_base_address, req => ptr_deref_1971_base_resize_req_0, ack => ptr_deref_1971_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1985_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp106_1885, dout => ptr_deref_1985_resized_base_address, req => ptr_deref_1985_base_resize_req_0, ack => ptr_deref_1985_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1993_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp109_1889, dout => ptr_deref_1993_resized_base_address, req => ptr_deref_1993_base_resize_req_0, ack => ptr_deref_1993_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2021_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp113_2019, dout => ptr_deref_2021_resized_base_address, req => ptr_deref_2021_base_resize_req_0, ack => ptr_deref_2021_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2045_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp116_2043, dout => ptr_deref_2045_resized_base_address, req => ptr_deref_2045_base_resize_req_0, ack => ptr_deref_2045_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2069_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp119_2067, dout => ptr_deref_2069_resized_base_address, req => ptr_deref_2069_base_resize_req_0, ack => ptr_deref_2069_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2093_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp122_2091, dout => ptr_deref_2093_resized_base_address, req => ptr_deref_2093_base_resize_req_0, ack => ptr_deref_2093_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2117_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2115, dout => ptr_deref_2117_resized_base_address, req => ptr_deref_2117_base_resize_req_0, ack => ptr_deref_2117_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2141_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp128_2139, dout => ptr_deref_2141_resized_base_address, req => ptr_deref_2141_base_resize_req_0, ack => ptr_deref_2141_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2165_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp131_2163, dout => ptr_deref_2165_resized_base_address, req => ptr_deref_2165_base_resize_req_0, ack => ptr_deref_2165_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2183_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp134_2181, dout => ptr_deref_2183_resized_base_address, req => ptr_deref_2183_base_resize_req_0, ack => ptr_deref_2183_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1613_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp4x_xi_1609, dout => tmp5x_xi_1614, req => type_cast_1613_inst_req_0, ack => type_cast_1613_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1618_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp4x_xi_1609, dout => tmp71_1619, req => type_cast_1618_inst_req_0, ack => type_cast_1618_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1642_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp80_1639, dout => tmp81_1643, req => type_cast_1642_inst_req_0, ack => type_cast_1642_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1667_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => wordx_x0x_xbe_2003, dout => type_cast_1667_wire, req => type_cast_1667_inst_req_0, ack => type_cast_1667_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1695_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 32, flow_through => false ) 
      port map( din => tmp74_1692, dout => tmp75_1696, req => type_cast_1695_inst_req_0, ack => type_cast_1695_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1716_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp1_1713, dout => tmp2_1717, req => type_cast_1716_inst_req_0, ack => type_cast_1716_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1730_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp4_1727, dout => tmp5_1731, req => type_cast_1730_inst_req_0, ack => type_cast_1730_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1744_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp7_1741, dout => tmp8_1745, req => type_cast_1744_inst_req_0, ack => type_cast_1744_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1758_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp10_1755, dout => tmp11_1759, req => type_cast_1758_inst_req_0, ack => type_cast_1758_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1772_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp13_1769, dout => tmp14_1773, req => type_cast_1772_inst_req_0, ack => type_cast_1772_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1786_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp16_1783, dout => tmp17_1787, req => type_cast_1786_inst_req_0, ack => type_cast_1786_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1800_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp19_1797, dout => tmp20_1801, req => type_cast_1800_inst_req_0, ack => type_cast_1800_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1808_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp73_1683, dout => tmp22_1809, req => type_cast_1808_inst_req_0, ack => type_cast_1808_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1898_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp24_1895, dout => tmp25_1899, req => type_cast_1898_inst_req_0, ack => type_cast_1898_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1912_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp27_1909, dout => tmp28_1913, req => type_cast_1912_inst_req_0, ack => type_cast_1912_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1926_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp30_1923, dout => tmp31_1927, req => type_cast_1926_inst_req_0, ack => type_cast_1926_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1940_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp33_1937, dout => tmp34_1941, req => type_cast_1940_inst_req_0, ack => type_cast_1940_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1954_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp36_1951, dout => tmp37_1955, req => type_cast_1954_inst_req_0, ack => type_cast_1954_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1968_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp39_1965, dout => tmp40_1969, req => type_cast_1968_inst_req_0, ack => type_cast_1968_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1982_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp42_1979, dout => tmp43_1983, req => type_cast_1982_inst_req_0, ack => type_cast_1982_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1990_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp73_1683, dout => tmp45_1991, req => type_cast_1990_inst_req_0, ack => type_cast_1990_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2014_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp47_2011, dout => tmp48_2015, req => type_cast_2014_inst_req_0, ack => type_cast_2014_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2032_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp50_2029, dout => tmp51_2033, req => type_cast_2032_inst_req_0, ack => type_cast_2032_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2056_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp53_2053, dout => tmp54_2057, req => type_cast_2056_inst_req_0, ack => type_cast_2056_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2080_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp56_2077, dout => tmp57_2081, req => type_cast_2080_inst_req_0, ack => type_cast_2080_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2104_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp59_2101, dout => tmp60_2105, req => type_cast_2104_inst_req_0, ack => type_cast_2104_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2128_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp62_2125, dout => tmp63_2129, req => type_cast_2128_inst_req_0, ack => type_cast_2128_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2152_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp65_2149, dout => tmp66_2153, req => type_cast_2152_inst_req_0, ack => type_cast_2152_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2170_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp73_1683, dout => tmp68_2171, req => type_cast_2170_inst_req_0, ack => type_cast_2170_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1860_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1860_index_0_rename_ack_0 <= array_obj_ref_1860_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1859_resized;
      simple_obj_ref_1859_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1864_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1864_index_0_rename_ack_0 <= array_obj_ref_1864_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1863_resized;
      simple_obj_ref_1863_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1868_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1868_index_0_rename_ack_0 <= array_obj_ref_1868_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1867_resized;
      simple_obj_ref_1867_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1872_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1872_index_0_rename_ack_0 <= array_obj_ref_1872_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1871_resized;
      simple_obj_ref_1871_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1876_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1876_index_0_rename_ack_0 <= array_obj_ref_1876_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1875_resized;
      simple_obj_ref_1875_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1880_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1880_index_0_rename_ack_0 <= array_obj_ref_1880_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1879_resized;
      simple_obj_ref_1879_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1884_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1884_index_0_rename_ack_0 <= array_obj_ref_1884_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1883_resized;
      simple_obj_ref_1883_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1888_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1888_index_0_rename_ack_0 <= array_obj_ref_1888_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1887_resized;
      simple_obj_ref_1887_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2018_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2018_index_0_rename_ack_0 <= array_obj_ref_2018_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2017_resized;
      simple_obj_ref_2017_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2042_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2042_index_0_rename_ack_0 <= array_obj_ref_2042_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2041_resized;
      simple_obj_ref_2041_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2066_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2066_index_0_rename_ack_0 <= array_obj_ref_2066_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2065_resized;
      simple_obj_ref_2065_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2090_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2090_index_0_rename_ack_0 <= array_obj_ref_2090_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2089_resized;
      simple_obj_ref_2089_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2114_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2114_index_0_rename_ack_0 <= array_obj_ref_2114_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2113_resized;
      simple_obj_ref_2113_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2138_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2138_index_0_rename_ack_0 <= array_obj_ref_2138_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2137_resized;
      simple_obj_ref_2137_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2162_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2162_index_0_rename_ack_0 <= array_obj_ref_2162_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2161_resized;
      simple_obj_ref_2161_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2180_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2180_index_0_rename_ack_0 <= array_obj_ref_2180_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2179_resized;
      simple_obj_ref_2179_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1554_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1554_gather_scatter_ack_0 <= ptr_deref_1554_gather_scatter_req_0;
      aggregated_sig <= type_cast_1556_wire_constant;
      ptr_deref_1554_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1719_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1719_addr_0_ack_0 <= ptr_deref_1719_addr_0_req_0;
      aggregated_sig <= ptr_deref_1719_root_address;
      ptr_deref_1719_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1719_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1719_gather_scatter_ack_0 <= ptr_deref_1719_gather_scatter_req_0;
      aggregated_sig <= tmp2_1717;
      ptr_deref_1719_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1719_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1719_root_address_inst_ack_0 <= ptr_deref_1719_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1719_resized_base_address;
      ptr_deref_1719_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1733_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1733_addr_0_ack_0 <= ptr_deref_1733_addr_0_req_0;
      aggregated_sig <= ptr_deref_1733_root_address;
      ptr_deref_1733_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1733_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1733_gather_scatter_ack_0 <= ptr_deref_1733_gather_scatter_req_0;
      aggregated_sig <= tmp5_1731;
      ptr_deref_1733_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1733_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1733_root_address_inst_ack_0 <= ptr_deref_1733_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1733_resized_base_address;
      ptr_deref_1733_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1747_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1747_addr_0_ack_0 <= ptr_deref_1747_addr_0_req_0;
      aggregated_sig <= ptr_deref_1747_root_address;
      ptr_deref_1747_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1747_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1747_gather_scatter_ack_0 <= ptr_deref_1747_gather_scatter_req_0;
      aggregated_sig <= tmp8_1745;
      ptr_deref_1747_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1747_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1747_root_address_inst_ack_0 <= ptr_deref_1747_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1747_resized_base_address;
      ptr_deref_1747_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1761_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1761_addr_0_ack_0 <= ptr_deref_1761_addr_0_req_0;
      aggregated_sig <= ptr_deref_1761_root_address;
      ptr_deref_1761_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1761_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1761_gather_scatter_ack_0 <= ptr_deref_1761_gather_scatter_req_0;
      aggregated_sig <= tmp11_1759;
      ptr_deref_1761_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1761_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1761_root_address_inst_ack_0 <= ptr_deref_1761_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1761_resized_base_address;
      ptr_deref_1761_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1775_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1775_addr_0_ack_0 <= ptr_deref_1775_addr_0_req_0;
      aggregated_sig <= ptr_deref_1775_root_address;
      ptr_deref_1775_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1775_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1775_gather_scatter_ack_0 <= ptr_deref_1775_gather_scatter_req_0;
      aggregated_sig <= tmp14_1773;
      ptr_deref_1775_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1775_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1775_root_address_inst_ack_0 <= ptr_deref_1775_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1775_resized_base_address;
      ptr_deref_1775_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1789_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1789_addr_0_ack_0 <= ptr_deref_1789_addr_0_req_0;
      aggregated_sig <= ptr_deref_1789_root_address;
      ptr_deref_1789_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1789_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1789_gather_scatter_ack_0 <= ptr_deref_1789_gather_scatter_req_0;
      aggregated_sig <= tmp17_1787;
      ptr_deref_1789_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1789_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1789_root_address_inst_ack_0 <= ptr_deref_1789_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1789_resized_base_address;
      ptr_deref_1789_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1803_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1803_addr_0_ack_0 <= ptr_deref_1803_addr_0_req_0;
      aggregated_sig <= ptr_deref_1803_root_address;
      ptr_deref_1803_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1803_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1803_gather_scatter_ack_0 <= ptr_deref_1803_gather_scatter_req_0;
      aggregated_sig <= tmp20_1801;
      ptr_deref_1803_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1803_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1803_root_address_inst_ack_0 <= ptr_deref_1803_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1803_resized_base_address;
      ptr_deref_1803_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1811_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1811_addr_0_ack_0 <= ptr_deref_1811_addr_0_req_0;
      aggregated_sig <= ptr_deref_1811_root_address;
      ptr_deref_1811_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1811_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1811_gather_scatter_ack_0 <= ptr_deref_1811_gather_scatter_req_0;
      aggregated_sig <= tmp22_1809;
      ptr_deref_1811_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1811_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1811_root_address_inst_ack_0 <= ptr_deref_1811_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1811_resized_base_address;
      ptr_deref_1811_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1901_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1901_addr_0_ack_0 <= ptr_deref_1901_addr_0_req_0;
      aggregated_sig <= ptr_deref_1901_root_address;
      ptr_deref_1901_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1901_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1901_gather_scatter_ack_0 <= ptr_deref_1901_gather_scatter_req_0;
      aggregated_sig <= tmp25_1899;
      ptr_deref_1901_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1901_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1901_root_address_inst_ack_0 <= ptr_deref_1901_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1901_resized_base_address;
      ptr_deref_1901_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1915_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1915_addr_0_ack_0 <= ptr_deref_1915_addr_0_req_0;
      aggregated_sig <= ptr_deref_1915_root_address;
      ptr_deref_1915_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1915_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1915_gather_scatter_ack_0 <= ptr_deref_1915_gather_scatter_req_0;
      aggregated_sig <= tmp28_1913;
      ptr_deref_1915_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1915_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1915_root_address_inst_ack_0 <= ptr_deref_1915_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1915_resized_base_address;
      ptr_deref_1915_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1929_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1929_addr_0_ack_0 <= ptr_deref_1929_addr_0_req_0;
      aggregated_sig <= ptr_deref_1929_root_address;
      ptr_deref_1929_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1929_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1929_gather_scatter_ack_0 <= ptr_deref_1929_gather_scatter_req_0;
      aggregated_sig <= tmp31_1927;
      ptr_deref_1929_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1929_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1929_root_address_inst_ack_0 <= ptr_deref_1929_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1929_resized_base_address;
      ptr_deref_1929_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1943_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1943_addr_0_ack_0 <= ptr_deref_1943_addr_0_req_0;
      aggregated_sig <= ptr_deref_1943_root_address;
      ptr_deref_1943_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1943_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1943_gather_scatter_ack_0 <= ptr_deref_1943_gather_scatter_req_0;
      aggregated_sig <= tmp34_1941;
      ptr_deref_1943_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1943_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1943_root_address_inst_ack_0 <= ptr_deref_1943_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1943_resized_base_address;
      ptr_deref_1943_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1957_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1957_addr_0_ack_0 <= ptr_deref_1957_addr_0_req_0;
      aggregated_sig <= ptr_deref_1957_root_address;
      ptr_deref_1957_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1957_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1957_gather_scatter_ack_0 <= ptr_deref_1957_gather_scatter_req_0;
      aggregated_sig <= tmp37_1955;
      ptr_deref_1957_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1957_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1957_root_address_inst_ack_0 <= ptr_deref_1957_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1957_resized_base_address;
      ptr_deref_1957_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1971_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1971_addr_0_ack_0 <= ptr_deref_1971_addr_0_req_0;
      aggregated_sig <= ptr_deref_1971_root_address;
      ptr_deref_1971_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1971_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1971_gather_scatter_ack_0 <= ptr_deref_1971_gather_scatter_req_0;
      aggregated_sig <= tmp40_1969;
      ptr_deref_1971_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1971_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1971_root_address_inst_ack_0 <= ptr_deref_1971_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1971_resized_base_address;
      ptr_deref_1971_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1985_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1985_addr_0_ack_0 <= ptr_deref_1985_addr_0_req_0;
      aggregated_sig <= ptr_deref_1985_root_address;
      ptr_deref_1985_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1985_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1985_gather_scatter_ack_0 <= ptr_deref_1985_gather_scatter_req_0;
      aggregated_sig <= tmp43_1983;
      ptr_deref_1985_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1985_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1985_root_address_inst_ack_0 <= ptr_deref_1985_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1985_resized_base_address;
      ptr_deref_1985_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1993_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1993_addr_0_ack_0 <= ptr_deref_1993_addr_0_req_0;
      aggregated_sig <= ptr_deref_1993_root_address;
      ptr_deref_1993_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1993_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1993_gather_scatter_ack_0 <= ptr_deref_1993_gather_scatter_req_0;
      aggregated_sig <= tmp45_1991;
      ptr_deref_1993_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1993_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1993_root_address_inst_ack_0 <= ptr_deref_1993_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1993_resized_base_address;
      ptr_deref_1993_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2021_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2021_addr_0_ack_0 <= ptr_deref_2021_addr_0_req_0;
      aggregated_sig <= ptr_deref_2021_root_address;
      ptr_deref_2021_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2021_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2021_gather_scatter_ack_0 <= ptr_deref_2021_gather_scatter_req_0;
      aggregated_sig <= tmp48_2015;
      ptr_deref_2021_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2021_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2021_root_address_inst_ack_0 <= ptr_deref_2021_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2021_resized_base_address;
      ptr_deref_2021_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2045_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2045_addr_0_ack_0 <= ptr_deref_2045_addr_0_req_0;
      aggregated_sig <= ptr_deref_2045_root_address;
      ptr_deref_2045_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2045_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2045_gather_scatter_ack_0 <= ptr_deref_2045_gather_scatter_req_0;
      aggregated_sig <= tmp51_2033;
      ptr_deref_2045_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2045_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2045_root_address_inst_ack_0 <= ptr_deref_2045_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2045_resized_base_address;
      ptr_deref_2045_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2069_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2069_addr_0_ack_0 <= ptr_deref_2069_addr_0_req_0;
      aggregated_sig <= ptr_deref_2069_root_address;
      ptr_deref_2069_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2069_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2069_gather_scatter_ack_0 <= ptr_deref_2069_gather_scatter_req_0;
      aggregated_sig <= tmp54_2057;
      ptr_deref_2069_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2069_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2069_root_address_inst_ack_0 <= ptr_deref_2069_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2069_resized_base_address;
      ptr_deref_2069_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2093_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2093_addr_0_ack_0 <= ptr_deref_2093_addr_0_req_0;
      aggregated_sig <= ptr_deref_2093_root_address;
      ptr_deref_2093_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2093_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2093_gather_scatter_ack_0 <= ptr_deref_2093_gather_scatter_req_0;
      aggregated_sig <= tmp57_2081;
      ptr_deref_2093_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2093_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2093_root_address_inst_ack_0 <= ptr_deref_2093_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2093_resized_base_address;
      ptr_deref_2093_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2117_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2117_addr_0_ack_0 <= ptr_deref_2117_addr_0_req_0;
      aggregated_sig <= ptr_deref_2117_root_address;
      ptr_deref_2117_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2117_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2117_gather_scatter_ack_0 <= ptr_deref_2117_gather_scatter_req_0;
      aggregated_sig <= tmp60_2105;
      ptr_deref_2117_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2117_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2117_root_address_inst_ack_0 <= ptr_deref_2117_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2117_resized_base_address;
      ptr_deref_2117_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2141_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2141_addr_0_ack_0 <= ptr_deref_2141_addr_0_req_0;
      aggregated_sig <= ptr_deref_2141_root_address;
      ptr_deref_2141_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2141_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2141_gather_scatter_ack_0 <= ptr_deref_2141_gather_scatter_req_0;
      aggregated_sig <= tmp63_2129;
      ptr_deref_2141_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2141_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2141_root_address_inst_ack_0 <= ptr_deref_2141_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2141_resized_base_address;
      ptr_deref_2141_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2165_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2165_addr_0_ack_0 <= ptr_deref_2165_addr_0_req_0;
      aggregated_sig <= ptr_deref_2165_root_address;
      ptr_deref_2165_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2165_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2165_gather_scatter_ack_0 <= ptr_deref_2165_gather_scatter_req_0;
      aggregated_sig <= tmp66_2153;
      ptr_deref_2165_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2165_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2165_root_address_inst_ack_0 <= ptr_deref_2165_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2165_resized_base_address;
      ptr_deref_2165_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2183_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2183_addr_0_ack_0 <= ptr_deref_2183_addr_0_req_0;
      aggregated_sig <= ptr_deref_2183_root_address;
      ptr_deref_2183_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2183_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2183_gather_scatter_ack_0 <= ptr_deref_2183_gather_scatter_req_0;
      aggregated_sig <= tmp68_2171;
      ptr_deref_2183_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2183_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2183_root_address_inst_ack_0 <= ptr_deref_2183_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2183_resized_base_address;
      ptr_deref_2183_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_1594_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp2x_xi_1593;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1594_branch_req_0,
          ack0 => if_stmt_1594_branch_ack_0,
          ack1 => if_stmt_1594_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1697_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1699_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1697_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_1697_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1697_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1702_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1697_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_1697_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1697_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_1699_wire_constant_cmp & expr_1702_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1697_branch_default_req_0,
          ack0 => switch_stmt_1697_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1623_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1623_resized_base_address;
      array_obj_ref_1623_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1623_root_address_inst_req_0,
          ackL => array_obj_ref_1623_root_address_inst_ack_0,
          reqR => array_obj_ref_1623_root_address_inst_req_1,
          ackR => array_obj_ref_1623_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1628_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1628_resized_base_address;
      array_obj_ref_1628_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1628_root_address_inst_req_0,
          ackL => array_obj_ref_1628_root_address_inst_ack_0,
          reqR => array_obj_ref_1628_root_address_inst_req_1,
          ackR => array_obj_ref_1628_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1633_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1633_resized_base_address;
      array_obj_ref_1633_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1633_root_address_inst_req_0,
          ackL => array_obj_ref_1633_root_address_inst_ack_0,
          reqR => array_obj_ref_1633_root_address_inst_req_1,
          ackR => array_obj_ref_1633_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1638_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1638_resized_base_address;
      array_obj_ref_1638_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1638_root_address_inst_req_0,
          ackL => array_obj_ref_1638_root_address_inst_ack_0,
          reqR => array_obj_ref_1638_root_address_inst_req_1,
          ackR => array_obj_ref_1638_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1647_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1647_resized_base_address;
      array_obj_ref_1647_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000101",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1647_root_address_inst_req_0,
          ackL => array_obj_ref_1647_root_address_inst_ack_0,
          reqR => array_obj_ref_1647_root_address_inst_req_1,
          ackR => array_obj_ref_1647_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1652_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1652_resized_base_address;
      array_obj_ref_1652_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000110",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1652_root_address_inst_req_0,
          ackL => array_obj_ref_1652_root_address_inst_ack_0,
          reqR => array_obj_ref_1652_root_address_inst_req_1,
          ackR => array_obj_ref_1652_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1657_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1657_resized_base_address;
      array_obj_ref_1657_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000111",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1657_root_address_inst_req_0,
          ackL => array_obj_ref_1657_root_address_inst_ack_0,
          reqR => array_obj_ref_1657_root_address_inst_req_1,
          ackR => array_obj_ref_1657_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_2018_root_address_inst array_obj_ref_1860_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2018_final_offset & array_obj_ref_2018_resized_base_address & array_obj_ref_1860_final_offset & array_obj_ref_1860_resized_base_address;
      array_obj_ref_2018_root_address <= data_out(21 downto 11);
      array_obj_ref_1860_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_2018_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1860_root_address_inst_req_0;
      array_obj_ref_2018_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1860_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_2018_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1860_root_address_inst_req_1;
      array_obj_ref_2018_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1860_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_2042_root_address_inst array_obj_ref_1864_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2042_final_offset & array_obj_ref_2042_resized_base_address & array_obj_ref_1864_final_offset & array_obj_ref_1864_resized_base_address;
      array_obj_ref_2042_root_address <= data_out(21 downto 11);
      array_obj_ref_1864_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_2042_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1864_root_address_inst_req_0;
      array_obj_ref_2042_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1864_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_2042_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1864_root_address_inst_req_1;
      array_obj_ref_2042_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1864_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_2066_root_address_inst array_obj_ref_1868_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2066_final_offset & array_obj_ref_2066_resized_base_address & array_obj_ref_1868_final_offset & array_obj_ref_1868_resized_base_address;
      array_obj_ref_2066_root_address <= data_out(21 downto 11);
      array_obj_ref_1868_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_2066_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1868_root_address_inst_req_0;
      array_obj_ref_2066_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1868_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_2066_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1868_root_address_inst_req_1;
      array_obj_ref_2066_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1868_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_2090_root_address_inst array_obj_ref_1872_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2090_final_offset & array_obj_ref_2090_resized_base_address & array_obj_ref_1872_final_offset & array_obj_ref_1872_resized_base_address;
      array_obj_ref_2090_root_address <= data_out(21 downto 11);
      array_obj_ref_1872_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_2090_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1872_root_address_inst_req_0;
      array_obj_ref_2090_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1872_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_2090_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1872_root_address_inst_req_1;
      array_obj_ref_2090_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1872_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1876_root_address_inst array_obj_ref_2114_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1876_final_offset & array_obj_ref_1876_resized_base_address & array_obj_ref_2114_final_offset & array_obj_ref_2114_resized_base_address;
      array_obj_ref_1876_root_address <= data_out(21 downto 11);
      array_obj_ref_2114_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1876_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_2114_root_address_inst_req_0;
      array_obj_ref_1876_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_2114_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1876_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_2114_root_address_inst_req_1;
      array_obj_ref_1876_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_2114_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1880_root_address_inst array_obj_ref_2138_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1880_final_offset & array_obj_ref_1880_resized_base_address & array_obj_ref_2138_final_offset & array_obj_ref_2138_resized_base_address;
      array_obj_ref_1880_root_address <= data_out(21 downto 11);
      array_obj_ref_2138_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1880_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_2138_root_address_inst_req_0;
      array_obj_ref_1880_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_2138_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1880_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_2138_root_address_inst_req_1;
      array_obj_ref_1880_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_2138_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_1884_root_address_inst array_obj_ref_2162_root_address_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1884_final_offset & array_obj_ref_1884_resized_base_address & array_obj_ref_2162_final_offset & array_obj_ref_2162_resized_base_address;
      array_obj_ref_1884_root_address <= data_out(21 downto 11);
      array_obj_ref_2162_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1884_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_2162_root_address_inst_req_0;
      array_obj_ref_1884_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_2162_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1884_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_2162_root_address_inst_req_1;
      array_obj_ref_1884_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_2162_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_1888_root_address_inst array_obj_ref_2180_root_address_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1888_final_offset & array_obj_ref_1888_resized_base_address & array_obj_ref_2180_final_offset & array_obj_ref_2180_resized_base_address;
      array_obj_ref_1888_root_address <= data_out(21 downto 11);
      array_obj_ref_2180_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1888_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_2180_root_address_inst_req_0;
      array_obj_ref_1888_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_2180_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1888_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_2180_root_address_inst_req_1;
      array_obj_ref_1888_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_2180_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1592_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xi_1587;
      tmp2x_xi_1593 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1592_inst_req_0,
          ackL => binary_1592_inst_ack_0,
          reqR => binary_1592_inst_req_1,
          ackR => binary_1592_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1673_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_1661;
      tmp137_1674 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1673_inst_req_0,
          ackL => binary_1673_inst_ack_0,
          reqR => binary_1673_inst_req_1,
          ackR => binary_1673_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1712_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp1_1713 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1712_inst_req_0,
          ackL => binary_1712_inst_ack_0,
          reqR => binary_1712_inst_req_1,
          ackR => binary_1712_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1726_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp4_1727 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1726_inst_req_0,
          ackL => binary_1726_inst_ack_0,
          reqR => binary_1726_inst_req_1,
          ackR => binary_1726_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1740_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp7_1741 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1740_inst_req_0,
          ackL => binary_1740_inst_ack_0,
          reqR => binary_1740_inst_req_1,
          ackR => binary_1740_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1754_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp10_1755 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1754_inst_req_0,
          ackL => binary_1754_inst_ack_0,
          reqR => binary_1754_inst_req_1,
          ackR => binary_1754_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1768_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp13_1769 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1768_inst_req_0,
          ackL => binary_1768_inst_ack_0,
          reqR => binary_1768_inst_req_1,
          ackR => binary_1768_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1782_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp16_1783 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1782_inst_req_0,
          ackL => binary_1782_inst_ack_0,
          reqR => binary_1782_inst_req_1,
          ackR => binary_1782_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1796_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp19_1797 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1796_inst_req_0,
          ackL => binary_1796_inst_ack_0,
          reqR => binary_1796_inst_req_1,
          ackR => binary_1796_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1820_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp144151_1821 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1820_inst_req_0,
          ackL => binary_1820_inst_ack_0,
          reqR => binary_1820_inst_req_1,
          ackR => binary_1820_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1826_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp143150_1827 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1826_inst_req_0,
          ackL => binary_1826_inst_ack_0,
          reqR => binary_1826_inst_req_1,
          ackR => binary_1826_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1832_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp142149_1833 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1832_inst_req_0,
          ackL => binary_1832_inst_ack_0,
          reqR => binary_1832_inst_req_1,
          ackR => binary_1832_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_1838_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp141148_1839 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1838_inst_req_0,
          ackL => binary_1838_inst_ack_0,
          reqR => binary_1838_inst_req_1,
          ackR => binary_1838_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_1844_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp140147_1845 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1844_inst_req_0,
          ackL => binary_1844_inst_ack_0,
          reqR => binary_1844_inst_req_1,
          ackR => binary_1844_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_1850_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp139146_1851 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1850_inst_req_0,
          ackL => binary_1850_inst_ack_0,
          reqR => binary_1850_inst_req_1,
          ackR => binary_1850_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_1856_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp138145_1857 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1856_inst_req_0,
          ackL => binary_1856_inst_ack_0,
          reqR => binary_1856_inst_req_1,
          ackR => binary_1856_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_1894_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp24_1895 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1894_inst_req_0,
          ackL => binary_1894_inst_ack_0,
          reqR => binary_1894_inst_req_1,
          ackR => binary_1894_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_1908_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp27_1909 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1908_inst_req_0,
          ackL => binary_1908_inst_ack_0,
          reqR => binary_1908_inst_req_1,
          ackR => binary_1908_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_1922_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp30_1923 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1922_inst_req_0,
          ackL => binary_1922_inst_ack_0,
          reqR => binary_1922_inst_req_1,
          ackR => binary_1922_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_1936_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp33_1937 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1936_inst_req_0,
          ackL => binary_1936_inst_ack_0,
          reqR => binary_1936_inst_req_1,
          ackR => binary_1936_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_1950_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp36_1951 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1950_inst_req_0,
          ackL => binary_1950_inst_ack_0,
          reqR => binary_1950_inst_req_1,
          ackR => binary_1950_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_1964_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp39_1965 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1964_inst_req_0,
          ackL => binary_1964_inst_ack_0,
          reqR => binary_1964_inst_req_1,
          ackR => binary_1964_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_1978_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp42_1979 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1978_inst_req_0,
          ackL => binary_1978_inst_ack_0,
          reqR => binary_1978_inst_req_1,
          ackR => binary_1978_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_2002_inst binary_2190_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_10_1661 & iNsTr_10_1661;
      wordx_x0x_xbe_2003 <= data_out(63 downto 32);
      tmp135_2191 <= data_out(31 downto 0);
      reqL(1) <= binary_2002_inst_req_0;
      reqL(0) <= binary_2190_inst_req_0;
      binary_2002_inst_ack_0 <= ackL(1);
      binary_2190_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_2002_inst_req_1;
      reqR(0) <= binary_2190_inst_req_1;
      binary_2002_inst_ack_1 <= ackR(1);
      binary_2190_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_2010_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp47_2011 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2010_inst_req_0,
          ackL => binary_2010_inst_ack_0,
          reqR => binary_2010_inst_req_1,
          ackR => binary_2010_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_2028_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp50_2029 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2028_inst_req_0,
          ackL => binary_2028_inst_ack_0,
          reqR => binary_2028_inst_req_1,
          ackR => binary_2028_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_2038_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp115_2039 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2038_inst_req_0,
          ackL => binary_2038_inst_ack_0,
          reqR => binary_2038_inst_req_1,
          ackR => binary_2038_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_2052_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp53_2053 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2052_inst_req_0,
          ackL => binary_2052_inst_ack_0,
          reqR => binary_2052_inst_req_1,
          ackR => binary_2052_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_2062_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp118_2063 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2062_inst_req_0,
          ackL => binary_2062_inst_ack_0,
          reqR => binary_2062_inst_req_1,
          ackR => binary_2062_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_2076_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp56_2077 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2076_inst_req_0,
          ackL => binary_2076_inst_ack_0,
          reqR => binary_2076_inst_req_1,
          ackR => binary_2076_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_2086_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp121_2087 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2086_inst_req_0,
          ackL => binary_2086_inst_ack_0,
          reqR => binary_2086_inst_req_1,
          ackR => binary_2086_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_2100_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp59_2101 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2100_inst_req_0,
          ackL => binary_2100_inst_ack_0,
          reqR => binary_2100_inst_req_1,
          ackR => binary_2100_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_2110_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp124_2111 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2110_inst_req_0,
          ackL => binary_2110_inst_ack_0,
          reqR => binary_2110_inst_req_1,
          ackR => binary_2110_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_2124_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp62_2125 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2124_inst_req_0,
          ackL => binary_2124_inst_ack_0,
          reqR => binary_2124_inst_req_1,
          ackR => binary_2124_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_2134_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp127_2135 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2134_inst_req_0,
          ackL => binary_2134_inst_ack_0,
          reqR => binary_2134_inst_req_1,
          ackR => binary_2134_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_2148_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp73_1683;
      tmp65_2149 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2148_inst_req_0,
          ackL => binary_2148_inst_ack_0,
          reqR => binary_2148_inst_req_1,
          ackR => binary_2148_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_2158_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp130_2159 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2158_inst_req_0,
          ackL => binary_2158_inst_ack_0,
          reqR => binary_2158_inst_req_1,
          ackR => binary_2158_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_2176_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp137_1674;
      tmp133_2177 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2176_inst_req_0,
          ackL => binary_2176_inst_ack_0,
          reqR => binary_2176_inst_req_1,
          ackR => binary_2176_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : switch_stmt_1697_select_expr_0 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp75_1696;
      expr_1699_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1697_select_expr_0_req_0,
          ackL => switch_stmt_1697_select_expr_0_ack_0,
          reqR => switch_stmt_1697_select_expr_0_req_1,
          ackR => switch_stmt_1697_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : switch_stmt_1697_select_expr_1 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp75_1696;
      expr_1702_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1697_select_expr_1_req_0,
          ackL => switch_stmt_1697_select_expr_1_ack_0,
          reqR => switch_stmt_1697_select_expr_1_req_1,
          ackR => switch_stmt_1697_select_expr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared store operator group (0) : ptr_deref_1554_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1554_store_0_req_0;
      ptr_deref_1554_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1554_store_0_req_1;
      ptr_deref_1554_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1554_word_address_0;
      data_in <= ptr_deref_1554_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(3 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1901_store_0 ptr_deref_2021_store_0 ptr_deref_1719_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1901_store_0_req_0;
      reqL(1) <= ptr_deref_2021_store_0_req_0;
      reqL(0) <= ptr_deref_1719_store_0_req_0;
      ptr_deref_1901_store_0_ack_0 <= ackL(2);
      ptr_deref_2021_store_0_ack_0 <= ackL(1);
      ptr_deref_1719_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1901_store_0_req_1;
      reqR(1) <= ptr_deref_2021_store_0_req_1;
      reqR(0) <= ptr_deref_1719_store_0_req_1;
      ptr_deref_1901_store_0_ack_1 <= ackR(2);
      ptr_deref_2021_store_0_ack_1 <= ackR(1);
      ptr_deref_1719_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1901_word_address_0 & ptr_deref_2021_word_address_0 & ptr_deref_1719_word_address_0;
      data_in <= ptr_deref_1901_data_0 & ptr_deref_2021_data_0 & ptr_deref_1719_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(7),
          mack => memory_space_3_sr_ack(7),
          maddr => memory_space_3_sr_addr(87 downto 77),
          mdata => memory_space_3_sr_data(63 downto 56),
          mtag => memory_space_3_sr_tag(15 downto 14),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(7),
          mack => memory_space_3_sc_ack(7),
          mtag => memory_space_3_sc_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_1915_store_0 ptr_deref_2045_store_0 ptr_deref_1733_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1915_store_0_req_0;
      reqL(1) <= ptr_deref_2045_store_0_req_0;
      reqL(0) <= ptr_deref_1733_store_0_req_0;
      ptr_deref_1915_store_0_ack_0 <= ackL(2);
      ptr_deref_2045_store_0_ack_0 <= ackL(1);
      ptr_deref_1733_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1915_store_0_req_1;
      reqR(1) <= ptr_deref_2045_store_0_req_1;
      reqR(0) <= ptr_deref_1733_store_0_req_1;
      ptr_deref_1915_store_0_ack_1 <= ackR(2);
      ptr_deref_2045_store_0_ack_1 <= ackR(1);
      ptr_deref_1733_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1915_word_address_0 & ptr_deref_2045_word_address_0 & ptr_deref_1733_word_address_0;
      data_in <= ptr_deref_1915_data_0 & ptr_deref_2045_data_0 & ptr_deref_1733_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(6),
          mack => memory_space_3_sr_ack(6),
          maddr => memory_space_3_sr_addr(76 downto 66),
          mdata => memory_space_3_sr_data(55 downto 48),
          mtag => memory_space_3_sr_tag(13 downto 12),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(6),
          mack => memory_space_3_sc_ack(6),
          mtag => memory_space_3_sc_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_1747_store_0 ptr_deref_1929_store_0 ptr_deref_2069_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1747_store_0_req_0;
      reqL(1) <= ptr_deref_1929_store_0_req_0;
      reqL(0) <= ptr_deref_2069_store_0_req_0;
      ptr_deref_1747_store_0_ack_0 <= ackL(2);
      ptr_deref_1929_store_0_ack_0 <= ackL(1);
      ptr_deref_2069_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1747_store_0_req_1;
      reqR(1) <= ptr_deref_1929_store_0_req_1;
      reqR(0) <= ptr_deref_2069_store_0_req_1;
      ptr_deref_1747_store_0_ack_1 <= ackR(2);
      ptr_deref_1929_store_0_ack_1 <= ackR(1);
      ptr_deref_2069_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1747_word_address_0 & ptr_deref_1929_word_address_0 & ptr_deref_2069_word_address_0;
      data_in <= ptr_deref_1747_data_0 & ptr_deref_1929_data_0 & ptr_deref_2069_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(5),
          mack => memory_space_3_sr_ack(5),
          maddr => memory_space_3_sr_addr(65 downto 55),
          mdata => memory_space_3_sr_data(47 downto 40),
          mtag => memory_space_3_sr_tag(11 downto 10),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(5),
          mack => memory_space_3_sc_ack(5),
          mtag => memory_space_3_sc_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_1943_store_0 ptr_deref_1761_store_0 ptr_deref_2093_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1943_store_0_req_0;
      reqL(1) <= ptr_deref_1761_store_0_req_0;
      reqL(0) <= ptr_deref_2093_store_0_req_0;
      ptr_deref_1943_store_0_ack_0 <= ackL(2);
      ptr_deref_1761_store_0_ack_0 <= ackL(1);
      ptr_deref_2093_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1943_store_0_req_1;
      reqR(1) <= ptr_deref_1761_store_0_req_1;
      reqR(0) <= ptr_deref_2093_store_0_req_1;
      ptr_deref_1943_store_0_ack_1 <= ackR(2);
      ptr_deref_1761_store_0_ack_1 <= ackR(1);
      ptr_deref_2093_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1943_word_address_0 & ptr_deref_1761_word_address_0 & ptr_deref_2093_word_address_0;
      data_in <= ptr_deref_1943_data_0 & ptr_deref_1761_data_0 & ptr_deref_2093_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(4),
          mack => memory_space_3_sr_ack(4),
          maddr => memory_space_3_sr_addr(54 downto 44),
          mdata => memory_space_3_sr_data(39 downto 32),
          mtag => memory_space_3_sr_tag(9 downto 8),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(4),
          mack => memory_space_3_sc_ack(4),
          mtag => memory_space_3_sc_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_1957_store_0 ptr_deref_2117_store_0 ptr_deref_1775_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1957_store_0_req_0;
      reqL(1) <= ptr_deref_2117_store_0_req_0;
      reqL(0) <= ptr_deref_1775_store_0_req_0;
      ptr_deref_1957_store_0_ack_0 <= ackL(2);
      ptr_deref_2117_store_0_ack_0 <= ackL(1);
      ptr_deref_1775_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1957_store_0_req_1;
      reqR(1) <= ptr_deref_2117_store_0_req_1;
      reqR(0) <= ptr_deref_1775_store_0_req_1;
      ptr_deref_1957_store_0_ack_1 <= ackR(2);
      ptr_deref_2117_store_0_ack_1 <= ackR(1);
      ptr_deref_1775_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1957_word_address_0 & ptr_deref_2117_word_address_0 & ptr_deref_1775_word_address_0;
      data_in <= ptr_deref_1957_data_0 & ptr_deref_2117_data_0 & ptr_deref_1775_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(3),
          mack => memory_space_3_sr_ack(3),
          maddr => memory_space_3_sr_addr(43 downto 33),
          mdata => memory_space_3_sr_data(31 downto 24),
          mtag => memory_space_3_sr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(3),
          mack => memory_space_3_sc_ack(3),
          mtag => memory_space_3_sc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_1971_store_0 ptr_deref_2141_store_0 ptr_deref_1789_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1971_store_0_req_0;
      reqL(1) <= ptr_deref_2141_store_0_req_0;
      reqL(0) <= ptr_deref_1789_store_0_req_0;
      ptr_deref_1971_store_0_ack_0 <= ackL(2);
      ptr_deref_2141_store_0_ack_0 <= ackL(1);
      ptr_deref_1789_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1971_store_0_req_1;
      reqR(1) <= ptr_deref_2141_store_0_req_1;
      reqR(0) <= ptr_deref_1789_store_0_req_1;
      ptr_deref_1971_store_0_ack_1 <= ackR(2);
      ptr_deref_2141_store_0_ack_1 <= ackR(1);
      ptr_deref_1789_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1971_word_address_0 & ptr_deref_2141_word_address_0 & ptr_deref_1789_word_address_0;
      data_in <= ptr_deref_1971_data_0 & ptr_deref_2141_data_0 & ptr_deref_1789_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(2),
          mack => memory_space_3_sr_ack(2),
          maddr => memory_space_3_sr_addr(32 downto 22),
          mdata => memory_space_3_sr_data(23 downto 16),
          mtag => memory_space_3_sr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(2),
          mack => memory_space_3_sc_ack(2),
          mtag => memory_space_3_sc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_1985_store_0 ptr_deref_2165_store_0 ptr_deref_1803_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1985_store_0_req_0;
      reqL(1) <= ptr_deref_2165_store_0_req_0;
      reqL(0) <= ptr_deref_1803_store_0_req_0;
      ptr_deref_1985_store_0_ack_0 <= ackL(2);
      ptr_deref_2165_store_0_ack_0 <= ackL(1);
      ptr_deref_1803_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1985_store_0_req_1;
      reqR(1) <= ptr_deref_2165_store_0_req_1;
      reqR(0) <= ptr_deref_1803_store_0_req_1;
      ptr_deref_1985_store_0_ack_1 <= ackR(2);
      ptr_deref_2165_store_0_ack_1 <= ackR(1);
      ptr_deref_1803_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1985_word_address_0 & ptr_deref_2165_word_address_0 & ptr_deref_1803_word_address_0;
      data_in <= ptr_deref_1985_data_0 & ptr_deref_2165_data_0 & ptr_deref_1803_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(1),
          mack => memory_space_3_sr_ack(1),
          maddr => memory_space_3_sr_addr(21 downto 11),
          mdata => memory_space_3_sr_data(15 downto 8),
          mtag => memory_space_3_sr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(1),
          mack => memory_space_3_sc_ack(1),
          mtag => memory_space_3_sc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared store operator group (8) : ptr_deref_1993_store_0 ptr_deref_1811_store_0 ptr_deref_2183_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1993_store_0_req_0;
      reqL(1) <= ptr_deref_1811_store_0_req_0;
      reqL(0) <= ptr_deref_2183_store_0_req_0;
      ptr_deref_1993_store_0_ack_0 <= ackL(2);
      ptr_deref_1811_store_0_ack_0 <= ackL(1);
      ptr_deref_2183_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1993_store_0_req_1;
      reqR(1) <= ptr_deref_1811_store_0_req_1;
      reqR(0) <= ptr_deref_2183_store_0_req_1;
      ptr_deref_1993_store_0_ack_1 <= ackR(2);
      ptr_deref_1811_store_0_ack_1 <= ackR(1);
      ptr_deref_2183_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1993_word_address_0 & ptr_deref_1811_word_address_0 & ptr_deref_2183_word_address_0;
      data_in <= ptr_deref_1993_data_0 & ptr_deref_1811_data_0 & ptr_deref_2183_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(10 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    -- shared inport operator group (0) : simple_obj_ref_1565_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1565_inst_req_0;
      simple_obj_ref_1565_inst_ack_0 <= ack(0);
      tmp_1566 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => start_wrapper_input_pipe_read_req(0),
          oack => start_wrapper_input_pipe_read_ack(0),
          odata => start_wrapper_input_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1586_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1586_inst_req_0;
      simple_obj_ref_1586_inst_ack_0 <= ack(0);
      tmpx_xi_1587 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_ack_pipe_read_req(0),
          oack => free_queue_ack_pipe_read_ack(0),
          odata => free_queue_ack_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_1608_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1608_inst_req_0;
      simple_obj_ref_1608_inst_ack_0 <= ack(0);
      tmp4x_xi_1609 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_get_pipe_read_req(0),
          oack => free_queue_get_pipe_read_ack(0),
          odata => free_queue_get_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_1682_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1682_inst_req_0;
      simple_obj_ref_1682_inst_ack_0 <= ack(0);
      tmp73_1683 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_1691_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1691_inst_req_0;
      simple_obj_ref_1691_inst_ack_0 <= ack(0);
      tmp74_1692 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_ctrl_pipe_read_req(0),
          oack => in_ctrl_pipe_read_ack(0),
          odata => in_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : simple_obj_ref_1575_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1575_inst_req_0;
      simple_obj_ref_1575_inst_ack_0 <= ack(0);
      data_in <= type_cast_1577_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_2198_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2198_inst_req_0;
      simple_obj_ref_2198_inst_ack_0 <= ack(0);
      data_in <= tmp4x_xi_1609;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => midpipe_pipe_write_req(0),
          oack => midpipe_pipe_write_ack(0),
          odata => midpipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_2207_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2207_inst_req_0;
      simple_obj_ref_2207_inst_ack_0 <= ack(0);
      data_in <= tmp74_1692;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => last_ctrl_pipe_write_req(0),
          oack => last_ctrl_pipe_write_ack(0),
          odata => last_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : simple_obj_ref_2216_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2216_inst_req_0;
      simple_obj_ref_2216_inst_ack_0 <= ack(0);
      data_in <= tmp135_2191;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => pkt_length_pipe_write_req(0),
          oack => pkt_length_pipe_write_ack(0),
          odata => pkt_length_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_output is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_3_lr_req : out  std_logic_vector(7 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(87 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(15 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(7 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(15 downto 0);
    midpipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    midpipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    midpipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    last_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    last_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    last_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    pkt_length_pipe_read_req : out  std_logic_vector(0 downto 0);
    pkt_length_pipe_read_ack : in   std_logic_vector(0 downto 0);
    pkt_length_pipe_read_data : in   std_logic_vector(31 downto 0);
    start_wrapper_output_pipe_read_req : out  std_logic_vector(0 downto 0);
    start_wrapper_output_pipe_read_ack : in   std_logic_vector(0 downto 0);
    start_wrapper_output_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
    op_lut_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    op_lut_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    op_lut_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    op_lut_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_output;
architecture Default of wrapper_output is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_output_CP_10224_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_2505_base_resize_req_0 : boolean;
  signal binary_2681_inst_req_0 : boolean;
  signal ptr_deref_2395_addr_0_ack_0 : boolean;
  signal ptr_deref_2273_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2619_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2286_load_0_req_0 : boolean;
  signal type_cast_2277_inst_req_0 : boolean;
  signal array_obj_ref_2269_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_2458_inst_req_0 : boolean;
  signal binary_2425_inst_req_0 : boolean;
  signal array_obj_ref_2282_final_reg_ack_0 : boolean;
  signal ptr_deref_2395_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2282_base_resize_ack_0 : boolean;
  signal ptr_deref_2505_gather_scatter_ack_0 : boolean;
  signal binary_2430_inst_ack_1 : boolean;
  signal binary_2386_inst_req_1 : boolean;
  signal ptr_deref_2395_root_address_inst_req_0 : boolean;
  signal binary_2386_inst_ack_0 : boolean;
  signal binary_2430_inst_req_1 : boolean;
  signal array_obj_ref_2501_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_2255_inst_ack_0 : boolean;
  signal array_obj_ref_2282_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2395_gather_scatter_req_0 : boolean;
  signal ptr_deref_2376_load_0_ack_1 : boolean;
  signal simple_obj_ref_2264_inst_req_0 : boolean;
  signal ptr_deref_2395_load_0_req_0 : boolean;
  signal ptr_deref_2286_root_address_inst_ack_0 : boolean;
  signal binary_2440_inst_req_1 : boolean;
  signal binary_2629_inst_req_1 : boolean;
  signal simple_obj_ref_2448_inst_ack_0 : boolean;
  signal binary_2435_inst_req_0 : boolean;
  signal ptr_deref_2505_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2505_load_0_req_0 : boolean;
  signal ptr_deref_2619_load_0_req_1 : boolean;
  signal ptr_deref_2643_load_0_req_1 : boolean;
  signal binary_2430_inst_ack_0 : boolean;
  signal binary_2435_inst_ack_1 : boolean;
  signal ptr_deref_2619_load_0_ack_0 : boolean;
  signal ptr_deref_2395_load_0_ack_1 : boolean;
  signal ptr_deref_2505_base_resize_ack_0 : boolean;
  signal binary_2440_inst_ack_0 : boolean;
  signal binary_2465_inst_ack_1 : boolean;
  signal binary_2435_inst_req_1 : boolean;
  signal ptr_deref_2395_addr_0_req_0 : boolean;
  signal ptr_deref_2505_root_address_inst_req_0 : boolean;
  signal binary_2386_inst_ack_1 : boolean;
  signal simple_obj_ref_2264_inst_ack_0 : boolean;
  signal binary_2465_inst_req_1 : boolean;
  signal binary_2430_inst_req_0 : boolean;
  signal ptr_deref_2619_gather_scatter_req_0 : boolean;
  signal ptr_deref_2395_load_0_req_1 : boolean;
  signal binary_2440_inst_req_0 : boolean;
  signal ptr_deref_2286_addr_0_ack_0 : boolean;
  signal array_obj_ref_2269_final_reg_ack_0 : boolean;
  signal type_cast_2277_inst_ack_0 : boolean;
  signal ptr_deref_2273_load_0_req_1 : boolean;
  signal binary_2435_inst_ack_0 : boolean;
  signal ptr_deref_2286_load_0_ack_1 : boolean;
  signal ptr_deref_2643_load_0_ack_1 : boolean;
  signal ptr_deref_2286_base_resize_req_0 : boolean;
  signal ptr_deref_2273_load_0_ack_1 : boolean;
  signal ptr_deref_2286_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2269_base_resize_req_0 : boolean;
  signal binary_2425_inst_req_1 : boolean;
  signal ptr_deref_2273_base_resize_ack_0 : boolean;
  signal binary_2515_inst_req_1 : boolean;
  signal binary_2296_inst_req_0 : boolean;
  signal array_obj_ref_2269_final_reg_req_0 : boolean;
  signal array_obj_ref_2282_root_address_inst_req_0 : boolean;
  signal ptr_deref_2505_load_0_ack_0 : boolean;
  signal ptr_deref_2273_addr_0_ack_0 : boolean;
  signal array_obj_ref_2282_root_address_inst_ack_0 : boolean;
  signal binary_2296_inst_req_1 : boolean;
  signal ptr_deref_2273_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2501_base_resize_req_0 : boolean;
  signal ptr_deref_2286_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2519_offset_inst_ack_0 : boolean;
  signal binary_2465_inst_req_0 : boolean;
  signal ptr_deref_2286_load_0_req_1 : boolean;
  signal ptr_deref_2273_addr_0_req_0 : boolean;
  signal ptr_deref_2273_root_address_inst_req_0 : boolean;
  signal type_cast_2290_inst_ack_0 : boolean;
  signal array_obj_ref_2269_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2501_base_resize_ack_0 : boolean;
  signal ptr_deref_2273_base_resize_req_0 : boolean;
  signal array_obj_ref_2501_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_2242_inst_req_0 : boolean;
  signal ptr_deref_2286_base_resize_ack_0 : boolean;
  signal binary_2671_inst_req_0 : boolean;
  signal ptr_deref_2643_gather_scatter_ack_0 : boolean;
  signal binary_2605_inst_ack_1 : boolean;
  signal array_obj_ref_2269_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_2242_inst_ack_0 : boolean;
  signal ptr_deref_2286_addr_0_req_0 : boolean;
  signal array_obj_ref_2657_offset_inst_ack_0 : boolean;
  signal binary_2465_inst_ack_0 : boolean;
  signal ptr_deref_2376_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2269_base_resize_ack_0 : boolean;
  signal binary_2605_inst_ack_0 : boolean;
  signal array_obj_ref_2282_root_address_inst_req_1 : boolean;
  signal binary_2386_inst_req_0 : boolean;
  signal binary_2420_inst_req_0 : boolean;
  signal ptr_deref_2286_load_0_ack_0 : boolean;
  signal ptr_deref_2286_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2501_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2301_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2657_offset_inst_req_0 : boolean;
  signal binary_2296_inst_ack_1 : boolean;
  signal ptr_deref_2305_addr_0_req_0 : boolean;
  signal ptr_deref_2305_addr_0_ack_0 : boolean;
  signal ptr_deref_2305_base_resize_req_0 : boolean;
  signal array_obj_ref_2301_final_reg_req_0 : boolean;
  signal array_obj_ref_2301_final_reg_ack_0 : boolean;
  signal binary_2605_inst_req_1 : boolean;
  signal array_obj_ref_2269_root_address_inst_ack_1 : boolean;
  signal type_cast_2246_inst_req_0 : boolean;
  signal binary_2420_inst_ack_1 : boolean;
  signal type_cast_2290_inst_req_0 : boolean;
  signal simple_obj_ref_2448_inst_req_0 : boolean;
  signal ptr_deref_2273_gather_scatter_req_0 : boolean;
  signal ptr_deref_2395_base_resize_ack_0 : boolean;
  signal ptr_deref_2376_load_0_ack_0 : boolean;
  signal binary_2420_inst_req_1 : boolean;
  signal type_cast_2246_inst_ack_0 : boolean;
  signal ptr_deref_2305_load_0_ack_1 : boolean;
  signal ptr_deref_2305_gather_scatter_req_0 : boolean;
  signal ptr_deref_2505_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2391_root_address_inst_req_1 : boolean;
  signal binary_2425_inst_ack_1 : boolean;
  signal binary_2515_inst_ack_0 : boolean;
  signal ptr_deref_2273_load_0_req_0 : boolean;
  signal ptr_deref_2376_gather_scatter_ack_0 : boolean;
  signal binary_2410_inst_ack_1 : boolean;
  signal binary_2497_inst_ack_1 : boolean;
  signal binary_2410_inst_req_1 : boolean;
  signal array_obj_ref_2301_base_resize_req_0 : boolean;
  signal array_obj_ref_2501_offset_inst_req_0 : boolean;
  signal array_obj_ref_2301_base_resize_ack_0 : boolean;
  signal array_obj_ref_2282_final_reg_req_0 : boolean;
  signal array_obj_ref_2301_root_address_inst_req_0 : boolean;
  signal ptr_deref_2395_load_0_ack_0 : boolean;
  signal array_obj_ref_2391_root_address_inst_ack_1 : boolean;
  signal binary_2605_inst_req_0 : boolean;
  signal array_obj_ref_2501_final_reg_ack_0 : boolean;
  signal ptr_deref_2305_root_address_inst_req_0 : boolean;
  signal ptr_deref_2305_root_address_inst_ack_0 : boolean;
  signal binary_2296_inst_ack_0 : boolean;
  signal binary_2420_inst_ack_0 : boolean;
  signal array_obj_ref_2391_root_address_inst_ack_0 : boolean;
  signal binary_2497_inst_ack_0 : boolean;
  signal binary_2410_inst_ack_0 : boolean;
  signal ptr_deref_2376_load_0_req_1 : boolean;
  signal binary_2440_inst_ack_1 : boolean;
  signal binary_2315_inst_ack_0 : boolean;
  signal binary_2315_inst_req_1 : boolean;
  signal binary_2315_inst_ack_1 : boolean;
  signal ptr_deref_2305_load_0_req_1 : boolean;
  signal ptr_deref_2376_load_0_req_0 : boolean;
  signal array_obj_ref_2501_offset_inst_ack_0 : boolean;
  signal ptr_deref_2273_load_0_ack_0 : boolean;
  signal array_obj_ref_2391_final_reg_ack_0 : boolean;
  signal binary_2686_inst_req_0 : boolean;
  signal binary_2497_inst_req_0 : boolean;
  signal binary_2410_inst_req_0 : boolean;
  signal ptr_deref_2505_addr_0_ack_0 : boolean;
  signal array_obj_ref_2501_final_reg_req_0 : boolean;
  signal array_obj_ref_2391_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2519_index_0_resize_req_0 : boolean;
  signal ptr_deref_2643_load_0_req_0 : boolean;
  signal ptr_deref_2505_addr_0_req_0 : boolean;
  signal array_obj_ref_2391_final_reg_req_0 : boolean;
  signal binary_2415_inst_ack_1 : boolean;
  signal array_obj_ref_2501_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2643_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2501_index_0_resize_req_0 : boolean;
  signal binary_2415_inst_req_1 : boolean;
  signal ptr_deref_2505_load_0_req_1 : boolean;
  signal binary_2415_inst_req_0 : boolean;
  signal ptr_deref_2305_base_resize_ack_0 : boolean;
  signal array_obj_ref_2301_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2501_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2301_root_address_inst_req_1 : boolean;
  signal binary_2415_inst_ack_0 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal binary_2497_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal binary_2425_inst_ack_0 : boolean;
  signal array_obj_ref_2282_base_resize_req_0 : boolean;
  signal simple_obj_ref_2255_inst_req_0 : boolean;
  signal ptr_deref_2305_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2519_offset_inst_req_0 : boolean;
  signal simple_obj_ref_2458_inst_ack_0 : boolean;
  signal ptr_deref_2395_base_resize_req_0 : boolean;
  signal ptr_deref_2305_load_0_req_0 : boolean;
  signal ptr_deref_2305_load_0_ack_0 : boolean;
  signal binary_2315_inst_req_0 : boolean;
  signal ptr_deref_2619_load_0_ack_1 : boolean;
  signal binary_2405_inst_ack_1 : boolean;
  signal binary_2491_inst_ack_1 : boolean;
  signal binary_2405_inst_req_1 : boolean;
  signal binary_2491_inst_req_1 : boolean;
  signal binary_2405_inst_ack_0 : boolean;
  signal binary_2491_inst_ack_0 : boolean;
  signal array_obj_ref_2320_base_resize_req_0 : boolean;
  signal binary_2491_inst_req_0 : boolean;
  signal array_obj_ref_2320_base_resize_ack_0 : boolean;
  signal ptr_deref_2643_addr_0_ack_0 : boolean;
  signal array_obj_ref_2391_base_resize_ack_0 : boolean;
  signal binary_2405_inst_req_0 : boolean;
  signal array_obj_ref_2320_root_address_inst_req_0 : boolean;
  signal ptr_deref_2643_base_resize_ack_0 : boolean;
  signal type_cast_2665_inst_req_0 : boolean;
  signal ptr_deref_2523_base_resize_req_0 : boolean;
  signal ptr_deref_2523_base_resize_ack_0 : boolean;
  signal ptr_deref_2523_root_address_inst_req_0 : boolean;
  signal ptr_deref_2523_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2619_base_resize_ack_0 : boolean;
  signal ptr_deref_2523_addr_0_req_0 : boolean;
  signal ptr_deref_2523_addr_0_ack_0 : boolean;
  signal ptr_deref_2619_base_resize_req_0 : boolean;
  signal array_obj_ref_2501_root_address_inst_req_1 : boolean;
  signal binary_2696_inst_ack_0 : boolean;
  signal array_obj_ref_2519_final_reg_ack_0 : boolean;
  signal ptr_deref_2643_load_0_ack_0 : boolean;
  signal binary_2706_inst_ack_1 : boolean;
  signal ptr_deref_2619_load_0_req_0 : boolean;
  signal if_stmt_2714_branch_req_0 : boolean;
  signal array_obj_ref_2519_base_resize_req_0 : boolean;
  signal array_obj_ref_2519_root_address_inst_req_0 : boolean;
  signal ptr_deref_2619_addr_0_req_0 : boolean;
  signal array_obj_ref_2519_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2643_addr_0_req_0 : boolean;
  signal simple_obj_ref_2721_inst_ack_0 : boolean;
  signal array_obj_ref_2519_root_address_inst_req_1 : boolean;
  signal type_cast_2599_inst_req_0 : boolean;
  signal array_obj_ref_2519_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2619_addr_0_ack_0 : boolean;
  signal binary_2629_inst_ack_0 : boolean;
  signal ptr_deref_2619_root_address_inst_ack_0 : boolean;
  signal type_cast_2380_inst_req_0 : boolean;
  signal array_obj_ref_2519_final_reg_req_0 : boolean;
  signal binary_2515_inst_ack_1 : boolean;
  signal binary_2706_inst_req_0 : boolean;
  signal type_cast_2380_inst_ack_0 : boolean;
  signal ptr_deref_2619_root_address_inst_req_0 : boolean;
  signal ptr_deref_2643_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2643_root_address_inst_req_0 : boolean;
  signal type_cast_2665_inst_ack_0 : boolean;
  signal binary_2696_inst_ack_1 : boolean;
  signal array_obj_ref_2519_base_resize_ack_0 : boolean;
  signal simple_obj_ref_2231_inst_req_0 : boolean;
  signal simple_obj_ref_2231_inst_ack_0 : boolean;
  signal array_obj_ref_2320_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2320_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2320_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2519_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2519_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2391_base_resize_req_0 : boolean;
  signal array_obj_ref_2501_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2320_final_reg_req_0 : boolean;
  signal array_obj_ref_2320_final_reg_ack_0 : boolean;
  signal array_obj_ref_2519_index_0_resize_ack_0 : boolean;
  signal binary_2485_inst_ack_1 : boolean;
  signal binary_2485_inst_req_1 : boolean;
  signal binary_2485_inst_ack_0 : boolean;
  signal type_cast_2399_inst_ack_0 : boolean;
  signal binary_2485_inst_req_0 : boolean;
  signal type_cast_2399_inst_req_0 : boolean;
  signal type_cast_2509_inst_ack_0 : boolean;
  signal ptr_deref_2324_base_resize_req_0 : boolean;
  signal ptr_deref_2324_base_resize_ack_0 : boolean;
  signal binary_2515_inst_req_0 : boolean;
  signal ptr_deref_2324_root_address_inst_req_0 : boolean;
  signal ptr_deref_2324_root_address_inst_ack_0 : boolean;
  signal type_cast_2509_inst_req_0 : boolean;
  signal ptr_deref_2324_addr_0_req_0 : boolean;
  signal ptr_deref_2324_addr_0_ack_0 : boolean;
  signal ptr_deref_2324_load_0_req_0 : boolean;
  signal ptr_deref_2324_load_0_ack_0 : boolean;
  signal type_cast_2480_inst_ack_0 : boolean;
  signal ptr_deref_2324_load_0_req_1 : boolean;
  signal type_cast_2480_inst_req_0 : boolean;
  signal ptr_deref_2324_load_0_ack_1 : boolean;
  signal ptr_deref_2505_load_0_ack_1 : boolean;
  signal ptr_deref_2324_gather_scatter_req_0 : boolean;
  signal ptr_deref_2324_gather_scatter_ack_0 : boolean;
  signal type_cast_2599_inst_ack_0 : boolean;
  signal array_obj_ref_2657_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2395_gather_scatter_ack_0 : boolean;
  signal type_cast_2328_inst_req_0 : boolean;
  signal type_cast_2328_inst_ack_0 : boolean;
  signal binary_2686_inst_req_1 : boolean;
  signal binary_2629_inst_ack_1 : boolean;
  signal binary_2334_inst_req_0 : boolean;
  signal binary_2334_inst_ack_0 : boolean;
  signal binary_2334_inst_req_1 : boolean;
  signal binary_2334_inst_ack_1 : boolean;
  signal binary_2676_inst_req_1 : boolean;
  signal binary_2611_inst_req_0 : boolean;
  signal binary_2611_inst_ack_0 : boolean;
  signal type_cast_2647_inst_req_0 : boolean;
  signal array_obj_ref_2339_base_resize_req_0 : boolean;
  signal type_cast_2647_inst_ack_0 : boolean;
  signal array_obj_ref_2339_base_resize_ack_0 : boolean;
  signal array_obj_ref_2339_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2657_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2339_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2339_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2339_root_address_inst_ack_1 : boolean;
  signal binary_2696_inst_req_0 : boolean;
  signal array_obj_ref_2339_final_reg_req_0 : boolean;
  signal array_obj_ref_2339_final_reg_ack_0 : boolean;
  signal binary_2653_inst_req_0 : boolean;
  signal binary_2676_inst_ack_1 : boolean;
  signal ptr_deref_2343_base_resize_req_0 : boolean;
  signal ptr_deref_2343_base_resize_ack_0 : boolean;
  signal binary_2686_inst_ack_1 : boolean;
  signal ptr_deref_2343_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2657_index_0_rename_ack_0 : boolean;
  signal ptr_deref_2343_root_address_inst_ack_0 : boolean;
  signal binary_2653_inst_ack_0 : boolean;
  signal ptr_deref_2343_addr_0_req_0 : boolean;
  signal ptr_deref_2343_addr_0_ack_0 : boolean;
  signal array_obj_ref_2657_index_0_resize_req_0 : boolean;
  signal binary_2653_inst_req_1 : boolean;
  signal ptr_deref_2343_load_0_req_0 : boolean;
  signal ptr_deref_2343_load_0_ack_0 : boolean;
  signal ptr_deref_2343_load_0_req_1 : boolean;
  signal binary_2611_inst_req_1 : boolean;
  signal ptr_deref_2343_load_0_ack_1 : boolean;
  signal ptr_deref_2343_gather_scatter_req_0 : boolean;
  signal ptr_deref_2343_gather_scatter_ack_0 : boolean;
  signal binary_2653_inst_ack_1 : boolean;
  signal type_cast_2623_inst_req_0 : boolean;
  signal type_cast_2623_inst_ack_0 : boolean;
  signal binary_2611_inst_ack_1 : boolean;
  signal binary_2696_inst_req_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal binary_2686_inst_ack_0 : boolean;
  signal binary_2353_inst_req_0 : boolean;
  signal binary_2353_inst_ack_0 : boolean;
  signal binary_2353_inst_req_1 : boolean;
  signal binary_2353_inst_ack_1 : boolean;
  signal array_obj_ref_2358_base_resize_req_0 : boolean;
  signal array_obj_ref_2358_base_resize_ack_0 : boolean;
  signal binary_2629_inst_req_0 : boolean;
  signal array_obj_ref_2358_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2358_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2358_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2358_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2358_final_reg_req_0 : boolean;
  signal array_obj_ref_2358_final_reg_ack_0 : boolean;
  signal ptr_deref_2362_base_resize_req_0 : boolean;
  signal ptr_deref_2362_base_resize_ack_0 : boolean;
  signal ptr_deref_2362_root_address_inst_req_0 : boolean;
  signal ptr_deref_2362_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2362_addr_0_req_0 : boolean;
  signal ptr_deref_2362_addr_0_ack_0 : boolean;
  signal ptr_deref_2362_load_0_req_0 : boolean;
  signal ptr_deref_2362_load_0_ack_0 : boolean;
  signal ptr_deref_2362_load_0_req_1 : boolean;
  signal ptr_deref_2362_load_0_ack_1 : boolean;
  signal ptr_deref_2362_gather_scatter_req_0 : boolean;
  signal ptr_deref_2362_gather_scatter_ack_0 : boolean;
  signal type_cast_2366_inst_req_0 : boolean;
  signal type_cast_2366_inst_ack_0 : boolean;
  signal binary_2372_inst_req_0 : boolean;
  signal binary_2372_inst_ack_0 : boolean;
  signal binary_2372_inst_req_1 : boolean;
  signal binary_2372_inst_ack_1 : boolean;
  signal ptr_deref_2376_base_resize_req_0 : boolean;
  signal ptr_deref_2376_base_resize_ack_0 : boolean;
  signal ptr_deref_2376_root_address_inst_req_0 : boolean;
  signal ptr_deref_2376_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2376_addr_0_req_0 : boolean;
  signal ptr_deref_2376_addr_0_ack_0 : boolean;
  signal ptr_deref_2523_load_0_req_0 : boolean;
  signal ptr_deref_2643_base_resize_req_0 : boolean;
  signal ptr_deref_2523_load_0_ack_0 : boolean;
  signal ptr_deref_2523_load_0_req_1 : boolean;
  signal ptr_deref_2523_load_0_ack_1 : boolean;
  signal ptr_deref_2523_gather_scatter_req_0 : boolean;
  signal ptr_deref_2523_gather_scatter_ack_0 : boolean;
  signal binary_2701_inst_req_1 : boolean;
  signal binary_2701_inst_ack_0 : boolean;
  signal binary_2706_inst_req_1 : boolean;
  signal binary_2706_inst_ack_0 : boolean;
  signal type_cast_2527_inst_req_0 : boolean;
  signal type_cast_2527_inst_ack_0 : boolean;
  signal if_stmt_2714_branch_ack_1 : boolean;
  signal binary_2533_inst_req_0 : boolean;
  signal binary_2533_inst_ack_0 : boolean;
  signal binary_2533_inst_req_1 : boolean;
  signal binary_2533_inst_ack_1 : boolean;
  signal array_obj_ref_2639_final_reg_ack_0 : boolean;
  signal binary_2539_inst_req_0 : boolean;
  signal binary_2539_inst_ack_0 : boolean;
  signal array_obj_ref_2639_final_reg_req_0 : boolean;
  signal binary_2539_inst_req_1 : boolean;
  signal binary_2539_inst_ack_1 : boolean;
  signal array_obj_ref_2639_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2639_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2639_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2639_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2615_final_reg_ack_0 : boolean;
  signal array_obj_ref_2543_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2543_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2615_final_reg_req_0 : boolean;
  signal binary_2691_inst_ack_1 : boolean;
  signal array_obj_ref_2543_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2543_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2543_offset_inst_req_0 : boolean;
  signal array_obj_ref_2543_offset_inst_ack_0 : boolean;
  signal binary_2691_inst_req_1 : boolean;
  signal array_obj_ref_2543_base_resize_req_0 : boolean;
  signal array_obj_ref_2543_base_resize_ack_0 : boolean;
  signal simple_obj_ref_2721_inst_req_0 : boolean;
  signal array_obj_ref_2615_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2639_base_resize_ack_0 : boolean;
  signal binary_2691_inst_ack_0 : boolean;
  signal array_obj_ref_2543_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2543_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2639_base_resize_req_0 : boolean;
  signal array_obj_ref_2543_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2543_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2615_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2543_final_reg_req_0 : boolean;
  signal array_obj_ref_2543_final_reg_ack_0 : boolean;
  signal array_obj_ref_2615_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2661_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2661_gather_scatter_req_0 : boolean;
  signal ptr_deref_2661_load_0_ack_1 : boolean;
  signal ptr_deref_2661_load_0_req_1 : boolean;
  signal array_obj_ref_2639_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2639_offset_inst_req_0 : boolean;
  signal array_obj_ref_2615_root_address_inst_req_0 : boolean;
  signal binary_2691_inst_req_0 : boolean;
  signal ptr_deref_2547_base_resize_req_0 : boolean;
  signal ptr_deref_2547_base_resize_ack_0 : boolean;
  signal ptr_deref_2547_root_address_inst_req_0 : boolean;
  signal ptr_deref_2547_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2547_addr_0_req_0 : boolean;
  signal ptr_deref_2661_load_0_ack_0 : boolean;
  signal ptr_deref_2547_addr_0_ack_0 : boolean;
  signal binary_2701_inst_ack_1 : boolean;
  signal ptr_deref_2661_load_0_req_0 : boolean;
  signal ptr_deref_2547_load_0_req_0 : boolean;
  signal array_obj_ref_2639_index_0_rename_ack_0 : boolean;
  signal ptr_deref_2547_load_0_ack_0 : boolean;
  signal ptr_deref_2547_load_0_req_1 : boolean;
  signal array_obj_ref_2639_index_0_rename_req_0 : boolean;
  signal ptr_deref_2547_load_0_ack_1 : boolean;
  signal ptr_deref_2547_gather_scatter_req_0 : boolean;
  signal ptr_deref_2547_gather_scatter_ack_0 : boolean;
  signal binary_2701_inst_req_0 : boolean;
  signal array_obj_ref_2615_base_resize_ack_0 : boolean;
  signal array_obj_ref_2639_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2639_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2615_base_resize_req_0 : boolean;
  signal type_cast_2551_inst_req_0 : boolean;
  signal ptr_deref_2661_addr_0_ack_0 : boolean;
  signal type_cast_2551_inst_ack_0 : boolean;
  signal binary_2676_inst_ack_0 : boolean;
  signal ptr_deref_2661_addr_0_req_0 : boolean;
  signal array_obj_ref_2615_offset_inst_ack_0 : boolean;
  signal binary_2557_inst_req_0 : boolean;
  signal ptr_deref_2661_root_address_inst_ack_0 : boolean;
  signal binary_2557_inst_ack_0 : boolean;
  signal ptr_deref_2661_root_address_inst_req_0 : boolean;
  signal binary_2557_inst_req_1 : boolean;
  signal binary_2557_inst_ack_1 : boolean;
  signal if_stmt_2714_branch_ack_0 : boolean;
  signal array_obj_ref_2615_offset_inst_req_0 : boolean;
  signal ptr_deref_2661_base_resize_ack_0 : boolean;
  signal ptr_deref_2661_base_resize_req_0 : boolean;
  signal binary_2563_inst_req_0 : boolean;
  signal binary_2563_inst_ack_0 : boolean;
  signal binary_2563_inst_req_1 : boolean;
  signal binary_2563_inst_ack_1 : boolean;
  signal array_obj_ref_2615_index_0_rename_ack_0 : boolean;
  signal binary_2635_inst_ack_1 : boolean;
  signal array_obj_ref_2615_index_0_rename_req_0 : boolean;
  signal binary_2635_inst_req_1 : boolean;
  signal binary_2635_inst_ack_0 : boolean;
  signal binary_2635_inst_req_0 : boolean;
  signal binary_2681_inst_ack_1 : boolean;
  signal binary_2676_inst_req_0 : boolean;
  signal array_obj_ref_2657_final_reg_ack_0 : boolean;
  signal array_obj_ref_2567_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2657_final_reg_req_0 : boolean;
  signal array_obj_ref_2567_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2567_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2567_index_0_rename_ack_0 : boolean;
  signal binary_2681_inst_req_1 : boolean;
  signal binary_2671_inst_ack_1 : boolean;
  signal array_obj_ref_2615_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2567_offset_inst_req_0 : boolean;
  signal array_obj_ref_2657_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2567_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2615_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2657_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2657_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2567_base_resize_req_0 : boolean;
  signal array_obj_ref_2657_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2567_base_resize_ack_0 : boolean;
  signal binary_2681_inst_ack_0 : boolean;
  signal binary_2671_inst_req_1 : boolean;
  signal array_obj_ref_2567_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2567_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2567_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2657_base_resize_ack_0 : boolean;
  signal array_obj_ref_2567_root_address_inst_ack_1 : boolean;
  signal binary_2671_inst_ack_0 : boolean;
  signal array_obj_ref_2657_base_resize_req_0 : boolean;
  signal array_obj_ref_2567_final_reg_req_0 : boolean;
  signal array_obj_ref_2567_final_reg_ack_0 : boolean;
  signal ptr_deref_2571_base_resize_req_0 : boolean;
  signal ptr_deref_2571_base_resize_ack_0 : boolean;
  signal ptr_deref_2571_root_address_inst_req_0 : boolean;
  signal ptr_deref_2571_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2571_addr_0_req_0 : boolean;
  signal ptr_deref_2571_addr_0_ack_0 : boolean;
  signal ptr_deref_2571_load_0_req_0 : boolean;
  signal ptr_deref_2571_load_0_ack_0 : boolean;
  signal ptr_deref_2571_load_0_req_1 : boolean;
  signal ptr_deref_2571_load_0_ack_1 : boolean;
  signal ptr_deref_2571_gather_scatter_req_0 : boolean;
  signal ptr_deref_2571_gather_scatter_ack_0 : boolean;
  signal type_cast_2575_inst_req_0 : boolean;
  signal type_cast_2575_inst_ack_0 : boolean;
  signal binary_2581_inst_req_0 : boolean;
  signal binary_2581_inst_ack_0 : boolean;
  signal binary_2581_inst_req_1 : boolean;
  signal binary_2581_inst_ack_1 : boolean;
  signal binary_2587_inst_req_0 : boolean;
  signal binary_2587_inst_ack_0 : boolean;
  signal binary_2587_inst_req_1 : boolean;
  signal binary_2587_inst_ack_1 : boolean;
  signal array_obj_ref_2591_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2591_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2591_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2591_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2591_offset_inst_req_0 : boolean;
  signal array_obj_ref_2591_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2591_base_resize_req_0 : boolean;
  signal array_obj_ref_2591_base_resize_ack_0 : boolean;
  signal array_obj_ref_2591_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2591_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2591_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2591_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2591_final_reg_req_0 : boolean;
  signal array_obj_ref_2591_final_reg_ack_0 : boolean;
  signal ptr_deref_2595_base_resize_req_0 : boolean;
  signal ptr_deref_2595_base_resize_ack_0 : boolean;
  signal ptr_deref_2595_root_address_inst_req_0 : boolean;
  signal ptr_deref_2595_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2595_addr_0_req_0 : boolean;
  signal ptr_deref_2595_addr_0_ack_0 : boolean;
  signal ptr_deref_2595_load_0_req_0 : boolean;
  signal ptr_deref_2595_load_0_ack_0 : boolean;
  signal ptr_deref_2595_load_0_req_1 : boolean;
  signal ptr_deref_2595_load_0_ack_1 : boolean;
  signal ptr_deref_2595_gather_scatter_req_0 : boolean;
  signal ptr_deref_2595_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_2731_inst_req_0 : boolean;
  signal simple_obj_ref_2731_inst_ack_0 : boolean;
  signal binary_2738_inst_req_0 : boolean;
  signal binary_2738_inst_ack_0 : boolean;
  signal binary_2738_inst_req_1 : boolean;
  signal binary_2738_inst_ack_1 : boolean;
  signal simple_obj_ref_2742_inst_req_0 : boolean;
  signal simple_obj_ref_2742_inst_ack_0 : boolean;
  signal simple_obj_ref_2751_inst_req_0 : boolean;
  signal simple_obj_ref_2751_inst_ack_0 : boolean;
  signal simple_obj_ref_2760_inst_req_0 : boolean;
  signal simple_obj_ref_2760_inst_ack_0 : boolean;
  signal simple_obj_ref_2770_inst_req_0 : boolean;
  signal simple_obj_ref_2770_inst_ack_0 : boolean;
  signal phi_stmt_2469_req_1 : boolean;
  signal type_cast_2473_inst_req_0 : boolean;
  signal type_cast_2473_inst_ack_0 : boolean;
  signal phi_stmt_2469_req_0 : boolean;
  signal phi_stmt_2469_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_output_CP_10224: Block -- control-path 
    signal cp_elements: BooleanArray(529 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    simple_obj_ref_2231_inst_req_0 <= cp_elements(0);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(500);
    cp_elements(3) <= OrReduce(cp_elements(507) & cp_elements(529));
    simple_obj_ref_2721_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= simple_obj_ref_2231_inst_ack_0;
    cp_elements(5) <= simple_obj_ref_2242_inst_ack_0;
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(8) & cp_elements(9));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2246_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= cp_elements(6);
    cp_elements(9) <= cp_elements(6);
    cp_elements(10) <= type_cast_2246_inst_ack_0;
    simple_obj_ref_2255_inst_req_0 <= cp_elements(10);
    cp_elements(11) <= simple_obj_ref_2255_inst_ack_0;
    simple_obj_ref_2264_inst_req_0 <= cp_elements(11);
    cp_elements(12) <= simple_obj_ref_2264_inst_ack_0;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= cp_elements(13);
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(19));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2269_final_reg_req_0 <= cp_elements(15);
    cp_elements(16) <= cp_elements(13);
    array_obj_ref_2269_base_resize_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_2269_base_resize_ack_0;
    array_obj_ref_2269_root_address_inst_req_0 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_2269_root_address_inst_ack_0;
    array_obj_ref_2269_root_address_inst_req_1 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_2269_root_address_inst_ack_1;
    cp_elements(20) <= array_obj_ref_2269_final_reg_ack_0;
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(20) & cp_elements(25));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2273_load_0_req_0 <= cp_elements(21);
    cp_elements(22) <= cp_elements(20);
    ptr_deref_2273_base_resize_req_0 <= cp_elements(22);
    cp_elements(23) <= ptr_deref_2273_base_resize_ack_0;
    ptr_deref_2273_root_address_inst_req_0 <= cp_elements(23);
    cp_elements(24) <= ptr_deref_2273_root_address_inst_ack_0;
    ptr_deref_2273_addr_0_req_0 <= cp_elements(24);
    cp_elements(25) <= ptr_deref_2273_addr_0_ack_0;
    cp_elements(26) <= ptr_deref_2273_load_0_ack_0;
    ptr_deref_2273_load_0_req_1 <= cp_elements(26);
    cp_elements(27) <= ptr_deref_2273_load_0_ack_1;
    ptr_deref_2273_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= ptr_deref_2273_gather_scatter_ack_0;
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(28) & cp_elements(30));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2277_inst_req_0 <= cp_elements(29);
    cp_elements(30) <= cp_elements(13);
    cp_elements(31) <= type_cast_2277_inst_ack_0;
    cp_elements(32) <= cp_elements(13);
    cpelement_group_33 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(37));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(33),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2282_final_reg_req_0 <= cp_elements(33);
    cp_elements(34) <= cp_elements(13);
    array_obj_ref_2282_base_resize_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_2282_base_resize_ack_0;
    array_obj_ref_2282_root_address_inst_req_0 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_2282_root_address_inst_ack_0;
    array_obj_ref_2282_root_address_inst_req_1 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_2282_root_address_inst_ack_1;
    cp_elements(38) <= array_obj_ref_2282_final_reg_ack_0;
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(38) & cp_elements(43));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2286_load_0_req_0 <= cp_elements(39);
    cp_elements(40) <= cp_elements(38);
    ptr_deref_2286_base_resize_req_0 <= cp_elements(40);
    cp_elements(41) <= ptr_deref_2286_base_resize_ack_0;
    ptr_deref_2286_root_address_inst_req_0 <= cp_elements(41);
    cp_elements(42) <= ptr_deref_2286_root_address_inst_ack_0;
    ptr_deref_2286_addr_0_req_0 <= cp_elements(42);
    cp_elements(43) <= ptr_deref_2286_addr_0_ack_0;
    cp_elements(44) <= ptr_deref_2286_load_0_ack_0;
    ptr_deref_2286_load_0_req_1 <= cp_elements(44);
    cp_elements(45) <= ptr_deref_2286_load_0_ack_1;
    ptr_deref_2286_gather_scatter_req_0 <= cp_elements(45);
    cp_elements(46) <= ptr_deref_2286_gather_scatter_ack_0;
    cpelement_group_47 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(46) & cp_elements(48));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(47),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2290_inst_req_0 <= cp_elements(47);
    cp_elements(48) <= cp_elements(13);
    cp_elements(49) <= type_cast_2290_inst_ack_0;
    cpelement_group_50 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(49) & cp_elements(51));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(50),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2296_inst_req_0 <= cp_elements(50);
    cp_elements(51) <= cp_elements(13);
    cp_elements(52) <= binary_2296_inst_ack_0;
    binary_2296_inst_req_1 <= cp_elements(52);
    cp_elements(53) <= binary_2296_inst_ack_1;
    cp_elements(54) <= cp_elements(13);
    cpelement_group_55 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(54) & cp_elements(59));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(55),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2301_final_reg_req_0 <= cp_elements(55);
    cp_elements(56) <= cp_elements(13);
    array_obj_ref_2301_base_resize_req_0 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_2301_base_resize_ack_0;
    array_obj_ref_2301_root_address_inst_req_0 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_2301_root_address_inst_ack_0;
    array_obj_ref_2301_root_address_inst_req_1 <= cp_elements(58);
    cp_elements(59) <= array_obj_ref_2301_root_address_inst_ack_1;
    cp_elements(60) <= array_obj_ref_2301_final_reg_ack_0;
    cpelement_group_61 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(65));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(61),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2305_load_0_req_0 <= cp_elements(61);
    cp_elements(62) <= cp_elements(60);
    ptr_deref_2305_base_resize_req_0 <= cp_elements(62);
    cp_elements(63) <= ptr_deref_2305_base_resize_ack_0;
    ptr_deref_2305_root_address_inst_req_0 <= cp_elements(63);
    cp_elements(64) <= ptr_deref_2305_root_address_inst_ack_0;
    ptr_deref_2305_addr_0_req_0 <= cp_elements(64);
    cp_elements(65) <= ptr_deref_2305_addr_0_ack_0;
    cp_elements(66) <= ptr_deref_2305_load_0_ack_0;
    ptr_deref_2305_load_0_req_1 <= cp_elements(66);
    cp_elements(67) <= ptr_deref_2305_load_0_ack_1;
    ptr_deref_2305_gather_scatter_req_0 <= cp_elements(67);
    cp_elements(68) <= ptr_deref_2305_gather_scatter_ack_0;
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(70));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2309_inst_req_0 <= cp_elements(69);
    cp_elements(70) <= cp_elements(13);
    cp_elements(71) <= type_cast_2309_inst_ack_0;
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(73));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2315_inst_req_0 <= cp_elements(72);
    cp_elements(73) <= cp_elements(13);
    cp_elements(74) <= binary_2315_inst_ack_0;
    binary_2315_inst_req_1 <= cp_elements(74);
    cp_elements(75) <= binary_2315_inst_ack_1;
    cp_elements(76) <= cp_elements(13);
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(81));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2320_final_reg_req_0 <= cp_elements(77);
    cp_elements(78) <= cp_elements(13);
    array_obj_ref_2320_base_resize_req_0 <= cp_elements(78);
    cp_elements(79) <= array_obj_ref_2320_base_resize_ack_0;
    array_obj_ref_2320_root_address_inst_req_0 <= cp_elements(79);
    cp_elements(80) <= array_obj_ref_2320_root_address_inst_ack_0;
    array_obj_ref_2320_root_address_inst_req_1 <= cp_elements(80);
    cp_elements(81) <= array_obj_ref_2320_root_address_inst_ack_1;
    cp_elements(82) <= array_obj_ref_2320_final_reg_ack_0;
    cpelement_group_83 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(87));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(83),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2324_load_0_req_0 <= cp_elements(83);
    cp_elements(84) <= cp_elements(82);
    ptr_deref_2324_base_resize_req_0 <= cp_elements(84);
    cp_elements(85) <= ptr_deref_2324_base_resize_ack_0;
    ptr_deref_2324_root_address_inst_req_0 <= cp_elements(85);
    cp_elements(86) <= ptr_deref_2324_root_address_inst_ack_0;
    ptr_deref_2324_addr_0_req_0 <= cp_elements(86);
    cp_elements(87) <= ptr_deref_2324_addr_0_ack_0;
    cp_elements(88) <= ptr_deref_2324_load_0_ack_0;
    ptr_deref_2324_load_0_req_1 <= cp_elements(88);
    cp_elements(89) <= ptr_deref_2324_load_0_ack_1;
    ptr_deref_2324_gather_scatter_req_0 <= cp_elements(89);
    cp_elements(90) <= ptr_deref_2324_gather_scatter_ack_0;
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(90) & cp_elements(92));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2328_inst_req_0 <= cp_elements(91);
    cp_elements(92) <= cp_elements(13);
    cp_elements(93) <= type_cast_2328_inst_ack_0;
    cpelement_group_94 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(94),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2334_inst_req_0 <= cp_elements(94);
    cp_elements(95) <= cp_elements(13);
    cp_elements(96) <= binary_2334_inst_ack_0;
    binary_2334_inst_req_1 <= cp_elements(96);
    cp_elements(97) <= binary_2334_inst_ack_1;
    cp_elements(98) <= cp_elements(13);
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(98) & cp_elements(103));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2339_final_reg_req_0 <= cp_elements(99);
    cp_elements(100) <= cp_elements(13);
    array_obj_ref_2339_base_resize_req_0 <= cp_elements(100);
    cp_elements(101) <= array_obj_ref_2339_base_resize_ack_0;
    array_obj_ref_2339_root_address_inst_req_0 <= cp_elements(101);
    cp_elements(102) <= array_obj_ref_2339_root_address_inst_ack_0;
    array_obj_ref_2339_root_address_inst_req_1 <= cp_elements(102);
    cp_elements(103) <= array_obj_ref_2339_root_address_inst_ack_1;
    cp_elements(104) <= array_obj_ref_2339_final_reg_ack_0;
    cpelement_group_105 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(104) & cp_elements(109));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(105),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2343_load_0_req_0 <= cp_elements(105);
    cp_elements(106) <= cp_elements(104);
    ptr_deref_2343_base_resize_req_0 <= cp_elements(106);
    cp_elements(107) <= ptr_deref_2343_base_resize_ack_0;
    ptr_deref_2343_root_address_inst_req_0 <= cp_elements(107);
    cp_elements(108) <= ptr_deref_2343_root_address_inst_ack_0;
    ptr_deref_2343_addr_0_req_0 <= cp_elements(108);
    cp_elements(109) <= ptr_deref_2343_addr_0_ack_0;
    cp_elements(110) <= ptr_deref_2343_load_0_ack_0;
    ptr_deref_2343_load_0_req_1 <= cp_elements(110);
    cp_elements(111) <= ptr_deref_2343_load_0_ack_1;
    ptr_deref_2343_gather_scatter_req_0 <= cp_elements(111);
    cp_elements(112) <= ptr_deref_2343_gather_scatter_ack_0;
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(112) & cp_elements(114));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2347_inst_req_0 <= cp_elements(113);
    cp_elements(114) <= cp_elements(13);
    cp_elements(115) <= type_cast_2347_inst_ack_0;
    cpelement_group_116 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(115) & cp_elements(117));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(116),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2353_inst_req_0 <= cp_elements(116);
    cp_elements(117) <= cp_elements(13);
    cp_elements(118) <= binary_2353_inst_ack_0;
    binary_2353_inst_req_1 <= cp_elements(118);
    cp_elements(119) <= binary_2353_inst_ack_1;
    cp_elements(120) <= cp_elements(13);
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(120) & cp_elements(125));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2358_final_reg_req_0 <= cp_elements(121);
    cp_elements(122) <= cp_elements(13);
    array_obj_ref_2358_base_resize_req_0 <= cp_elements(122);
    cp_elements(123) <= array_obj_ref_2358_base_resize_ack_0;
    array_obj_ref_2358_root_address_inst_req_0 <= cp_elements(123);
    cp_elements(124) <= array_obj_ref_2358_root_address_inst_ack_0;
    array_obj_ref_2358_root_address_inst_req_1 <= cp_elements(124);
    cp_elements(125) <= array_obj_ref_2358_root_address_inst_ack_1;
    cp_elements(126) <= array_obj_ref_2358_final_reg_ack_0;
    cpelement_group_127 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(126) & cp_elements(131));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(127),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2362_load_0_req_0 <= cp_elements(127);
    cp_elements(128) <= cp_elements(126);
    ptr_deref_2362_base_resize_req_0 <= cp_elements(128);
    cp_elements(129) <= ptr_deref_2362_base_resize_ack_0;
    ptr_deref_2362_root_address_inst_req_0 <= cp_elements(129);
    cp_elements(130) <= ptr_deref_2362_root_address_inst_ack_0;
    ptr_deref_2362_addr_0_req_0 <= cp_elements(130);
    cp_elements(131) <= ptr_deref_2362_addr_0_ack_0;
    cp_elements(132) <= ptr_deref_2362_load_0_ack_0;
    ptr_deref_2362_load_0_req_1 <= cp_elements(132);
    cp_elements(133) <= ptr_deref_2362_load_0_ack_1;
    ptr_deref_2362_gather_scatter_req_0 <= cp_elements(133);
    cp_elements(134) <= ptr_deref_2362_gather_scatter_ack_0;
    cpelement_group_135 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(136));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(135),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2366_inst_req_0 <= cp_elements(135);
    cp_elements(136) <= cp_elements(13);
    cp_elements(137) <= type_cast_2366_inst_ack_0;
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(139));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2372_inst_req_0 <= cp_elements(138);
    cp_elements(139) <= cp_elements(13);
    cp_elements(140) <= binary_2372_inst_ack_0;
    binary_2372_inst_req_1 <= cp_elements(140);
    cp_elements(141) <= binary_2372_inst_ack_1;
    cpelement_group_142 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(147));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(142),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2376_load_0_req_0 <= cp_elements(142);
    cp_elements(143) <= cp_elements(13);
    cp_elements(144) <= cp_elements(143);
    ptr_deref_2376_base_resize_req_0 <= cp_elements(144);
    cp_elements(145) <= ptr_deref_2376_base_resize_ack_0;
    ptr_deref_2376_root_address_inst_req_0 <= cp_elements(145);
    cp_elements(146) <= ptr_deref_2376_root_address_inst_ack_0;
    ptr_deref_2376_addr_0_req_0 <= cp_elements(146);
    cp_elements(147) <= ptr_deref_2376_addr_0_ack_0;
    cp_elements(148) <= ptr_deref_2376_load_0_ack_0;
    ptr_deref_2376_load_0_req_1 <= cp_elements(148);
    cp_elements(149) <= ptr_deref_2376_load_0_ack_1;
    ptr_deref_2376_gather_scatter_req_0 <= cp_elements(149);
    cp_elements(150) <= ptr_deref_2376_gather_scatter_ack_0;
    cpelement_group_151 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(150) & cp_elements(152));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(151),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2380_inst_req_0 <= cp_elements(151);
    cp_elements(152) <= cp_elements(13);
    cp_elements(153) <= type_cast_2380_inst_ack_0;
    cpelement_group_154 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(153) & cp_elements(155));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(154),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2386_inst_req_0 <= cp_elements(154);
    cp_elements(155) <= cp_elements(13);
    cp_elements(156) <= binary_2386_inst_ack_0;
    binary_2386_inst_req_1 <= cp_elements(156);
    cp_elements(157) <= binary_2386_inst_ack_1;
    cp_elements(158) <= cp_elements(13);
    cpelement_group_159 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(158) & cp_elements(163));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(159),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2391_final_reg_req_0 <= cp_elements(159);
    cp_elements(160) <= cp_elements(13);
    array_obj_ref_2391_base_resize_req_0 <= cp_elements(160);
    cp_elements(161) <= array_obj_ref_2391_base_resize_ack_0;
    array_obj_ref_2391_root_address_inst_req_0 <= cp_elements(161);
    cp_elements(162) <= array_obj_ref_2391_root_address_inst_ack_0;
    array_obj_ref_2391_root_address_inst_req_1 <= cp_elements(162);
    cp_elements(163) <= array_obj_ref_2391_root_address_inst_ack_1;
    cp_elements(164) <= array_obj_ref_2391_final_reg_ack_0;
    cpelement_group_165 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(164) & cp_elements(169));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(165),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2395_load_0_req_0 <= cp_elements(165);
    cp_elements(166) <= cp_elements(164);
    ptr_deref_2395_base_resize_req_0 <= cp_elements(166);
    cp_elements(167) <= ptr_deref_2395_base_resize_ack_0;
    ptr_deref_2395_root_address_inst_req_0 <= cp_elements(167);
    cp_elements(168) <= ptr_deref_2395_root_address_inst_ack_0;
    ptr_deref_2395_addr_0_req_0 <= cp_elements(168);
    cp_elements(169) <= ptr_deref_2395_addr_0_ack_0;
    cp_elements(170) <= ptr_deref_2395_load_0_ack_0;
    ptr_deref_2395_load_0_req_1 <= cp_elements(170);
    cp_elements(171) <= ptr_deref_2395_load_0_ack_1;
    ptr_deref_2395_gather_scatter_req_0 <= cp_elements(171);
    cp_elements(172) <= ptr_deref_2395_gather_scatter_ack_0;
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2399_inst_req_0 <= cp_elements(173);
    cp_elements(174) <= cp_elements(13);
    cp_elements(175) <= type_cast_2399_inst_ack_0;
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2405_inst_req_0 <= cp_elements(176);
    cp_elements(177) <= cp_elements(13);
    cp_elements(178) <= binary_2405_inst_ack_0;
    binary_2405_inst_req_1 <= cp_elements(178);
    cp_elements(179) <= binary_2405_inst_ack_1;
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(31) & cp_elements(53) & cp_elements(181));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2410_inst_req_0 <= cp_elements(180);
    cp_elements(181) <= cp_elements(13);
    cp_elements(182) <= binary_2410_inst_ack_0;
    binary_2410_inst_req_1 <= cp_elements(182);
    cp_elements(183) <= binary_2410_inst_ack_1;
    cpelement_group_184 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(183) & cp_elements(185));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(184),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2415_inst_req_0 <= cp_elements(184);
    cp_elements(185) <= cp_elements(13);
    cp_elements(186) <= binary_2415_inst_ack_0;
    binary_2415_inst_req_1 <= cp_elements(186);
    cp_elements(187) <= binary_2415_inst_ack_1;
    cpelement_group_188 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(97) & cp_elements(187) & cp_elements(189));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(188),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2420_inst_req_0 <= cp_elements(188);
    cp_elements(189) <= cp_elements(13);
    cp_elements(190) <= binary_2420_inst_ack_0;
    binary_2420_inst_req_1 <= cp_elements(190);
    cp_elements(191) <= binary_2420_inst_ack_1;
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(119) & cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2425_inst_req_0 <= cp_elements(192);
    cp_elements(193) <= cp_elements(13);
    cp_elements(194) <= binary_2425_inst_ack_0;
    binary_2425_inst_req_1 <= cp_elements(194);
    cp_elements(195) <= binary_2425_inst_ack_1;
    cpelement_group_196 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(141) & cp_elements(195) & cp_elements(197));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(196),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2430_inst_req_0 <= cp_elements(196);
    cp_elements(197) <= cp_elements(13);
    cp_elements(198) <= binary_2430_inst_ack_0;
    binary_2430_inst_req_1 <= cp_elements(198);
    cp_elements(199) <= binary_2430_inst_ack_1;
    cpelement_group_200 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(157) & cp_elements(199) & cp_elements(201));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2435_inst_req_0 <= cp_elements(200);
    cp_elements(201) <= cp_elements(13);
    cp_elements(202) <= binary_2435_inst_ack_0;
    binary_2435_inst_req_1 <= cp_elements(202);
    cp_elements(203) <= binary_2435_inst_ack_1;
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(203) & cp_elements(205));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2440_inst_req_0 <= cp_elements(204);
    cp_elements(205) <= cp_elements(13);
    cp_elements(206) <= binary_2440_inst_ack_0;
    binary_2440_inst_req_1 <= cp_elements(206);
    cp_elements(207) <= binary_2440_inst_ack_1;
    simple_obj_ref_2448_inst_req_0 <= cp_elements(207);
    cp_elements(208) <= simple_obj_ref_2448_inst_ack_0;
    simple_obj_ref_2458_inst_req_0 <= cp_elements(208);
    cp_elements(209) <= simple_obj_ref_2458_inst_ack_0;
    cp_elements(210) <= cp_elements(209);
    cpelement_group_211 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(212) & cp_elements(213));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2465_inst_req_0 <= cp_elements(211);
    cp_elements(212) <= cp_elements(210);
    cp_elements(213) <= cp_elements(210);
    cp_elements(214) <= binary_2465_inst_ack_0;
    binary_2465_inst_req_1 <= cp_elements(214);
    cp_elements(215) <= binary_2465_inst_ack_1;
    phi_stmt_2469_req_1 <= cp_elements(215);
    cp_elements(216) <= cp_elements(527);
    cpelement_group_217 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(219));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(217),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2480_inst_req_0 <= cp_elements(217);
    cp_elements(218) <= cp_elements(216);
    cp_elements(219) <= cp_elements(216);
    cp_elements(220) <= type_cast_2480_inst_ack_0;
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(222) & cp_elements(223) & cp_elements(224));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2485_inst_req_0 <= cp_elements(221);
    cp_elements(222) <= cp_elements(216);
    cp_elements(223) <= cp_elements(220);
    cp_elements(224) <= cp_elements(216);
    cp_elements(225) <= binary_2485_inst_ack_0;
    binary_2485_inst_req_1 <= cp_elements(225);
    cp_elements(226) <= binary_2485_inst_ack_1;
    cpelement_group_227 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(228) & cp_elements(229));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(227),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2491_inst_req_0 <= cp_elements(227);
    cp_elements(228) <= cp_elements(216);
    cp_elements(229) <= cp_elements(220);
    cp_elements(230) <= binary_2491_inst_ack_0;
    binary_2491_inst_req_1 <= cp_elements(230);
    cp_elements(231) <= binary_2491_inst_ack_1;
    cpelement_group_232 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(233) & cp_elements(234));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(232),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2497_inst_req_0 <= cp_elements(232);
    cp_elements(233) <= cp_elements(216);
    cp_elements(234) <= cp_elements(231);
    cp_elements(235) <= binary_2497_inst_ack_0;
    binary_2497_inst_req_1 <= cp_elements(235);
    cp_elements(236) <= binary_2497_inst_ack_1;
    array_obj_ref_2501_index_0_resize_req_0 <= cp_elements(236);
    cp_elements(237) <= cp_elements(216);
    cpelement_group_238 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(237) & cp_elements(246));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(238),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2501_final_reg_req_0 <= cp_elements(238);
    cp_elements(239) <= cp_elements(216);
    array_obj_ref_2501_base_resize_req_0 <= cp_elements(239);
    cp_elements(240) <= array_obj_ref_2501_index_0_resize_ack_0;
    array_obj_ref_2501_index_0_rename_req_0 <= cp_elements(240);
    cp_elements(241) <= array_obj_ref_2501_index_0_rename_ack_0;
    array_obj_ref_2501_offset_inst_req_0 <= cp_elements(241);
    cp_elements(242) <= array_obj_ref_2501_offset_inst_ack_0;
    cp_elements(243) <= array_obj_ref_2501_base_resize_ack_0;
    cpelement_group_244 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(242) & cp_elements(243));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(244),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2501_root_address_inst_req_0 <= cp_elements(244);
    cp_elements(245) <= array_obj_ref_2501_root_address_inst_ack_0;
    array_obj_ref_2501_root_address_inst_req_1 <= cp_elements(245);
    cp_elements(246) <= array_obj_ref_2501_root_address_inst_ack_1;
    cp_elements(247) <= array_obj_ref_2501_final_reg_ack_0;
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(247) & cp_elements(252));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2505_load_0_req_0 <= cp_elements(248);
    cp_elements(249) <= cp_elements(247);
    ptr_deref_2505_base_resize_req_0 <= cp_elements(249);
    cp_elements(250) <= ptr_deref_2505_base_resize_ack_0;
    ptr_deref_2505_root_address_inst_req_0 <= cp_elements(250);
    cp_elements(251) <= ptr_deref_2505_root_address_inst_ack_0;
    ptr_deref_2505_addr_0_req_0 <= cp_elements(251);
    cp_elements(252) <= ptr_deref_2505_addr_0_ack_0;
    cp_elements(253) <= ptr_deref_2505_load_0_ack_0;
    ptr_deref_2505_load_0_req_1 <= cp_elements(253);
    cp_elements(254) <= ptr_deref_2505_load_0_ack_1;
    ptr_deref_2505_gather_scatter_req_0 <= cp_elements(254);
    cp_elements(255) <= ptr_deref_2505_gather_scatter_ack_0;
    cpelement_group_256 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(255) & cp_elements(257));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(256),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2509_inst_req_0 <= cp_elements(256);
    cp_elements(257) <= cp_elements(216);
    cp_elements(258) <= type_cast_2509_inst_ack_0;
    cpelement_group_259 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(260) & cp_elements(261));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2515_inst_req_0 <= cp_elements(259);
    cp_elements(260) <= cp_elements(216);
    cp_elements(261) <= cp_elements(231);
    cp_elements(262) <= binary_2515_inst_ack_0;
    binary_2515_inst_req_1 <= cp_elements(262);
    cp_elements(263) <= binary_2515_inst_ack_1;
    array_obj_ref_2519_index_0_resize_req_0 <= cp_elements(263);
    cp_elements(264) <= cp_elements(216);
    cpelement_group_265 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(264) & cp_elements(273));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(265),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2519_final_reg_req_0 <= cp_elements(265);
    cp_elements(266) <= cp_elements(216);
    array_obj_ref_2519_base_resize_req_0 <= cp_elements(266);
    cp_elements(267) <= array_obj_ref_2519_index_0_resize_ack_0;
    array_obj_ref_2519_index_0_rename_req_0 <= cp_elements(267);
    cp_elements(268) <= array_obj_ref_2519_index_0_rename_ack_0;
    array_obj_ref_2519_offset_inst_req_0 <= cp_elements(268);
    cp_elements(269) <= array_obj_ref_2519_offset_inst_ack_0;
    cp_elements(270) <= array_obj_ref_2519_base_resize_ack_0;
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(269) & cp_elements(270));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2519_root_address_inst_req_0 <= cp_elements(271);
    cp_elements(272) <= array_obj_ref_2519_root_address_inst_ack_0;
    array_obj_ref_2519_root_address_inst_req_1 <= cp_elements(272);
    cp_elements(273) <= array_obj_ref_2519_root_address_inst_ack_1;
    cp_elements(274) <= array_obj_ref_2519_final_reg_ack_0;
    cpelement_group_275 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(279));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(275),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2523_load_0_req_0 <= cp_elements(275);
    cp_elements(276) <= cp_elements(274);
    ptr_deref_2523_base_resize_req_0 <= cp_elements(276);
    cp_elements(277) <= ptr_deref_2523_base_resize_ack_0;
    ptr_deref_2523_root_address_inst_req_0 <= cp_elements(277);
    cp_elements(278) <= ptr_deref_2523_root_address_inst_ack_0;
    ptr_deref_2523_addr_0_req_0 <= cp_elements(278);
    cp_elements(279) <= ptr_deref_2523_addr_0_ack_0;
    cp_elements(280) <= ptr_deref_2523_load_0_ack_0;
    ptr_deref_2523_load_0_req_1 <= cp_elements(280);
    cp_elements(281) <= ptr_deref_2523_load_0_ack_1;
    ptr_deref_2523_gather_scatter_req_0 <= cp_elements(281);
    cp_elements(282) <= ptr_deref_2523_gather_scatter_ack_0;
    cpelement_group_283 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(282) & cp_elements(284));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(283),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2527_inst_req_0 <= cp_elements(283);
    cp_elements(284) <= cp_elements(216);
    cp_elements(285) <= type_cast_2527_inst_ack_0;
    cpelement_group_286 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(285) & cp_elements(287));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(286),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2533_inst_req_0 <= cp_elements(286);
    cp_elements(287) <= cp_elements(216);
    cp_elements(288) <= binary_2533_inst_ack_0;
    binary_2533_inst_req_1 <= cp_elements(288);
    cp_elements(289) <= binary_2533_inst_ack_1;
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(292));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2539_inst_req_0 <= cp_elements(290);
    cp_elements(291) <= cp_elements(216);
    cp_elements(292) <= cp_elements(231);
    cp_elements(293) <= binary_2539_inst_ack_0;
    binary_2539_inst_req_1 <= cp_elements(293);
    cp_elements(294) <= binary_2539_inst_ack_1;
    array_obj_ref_2543_index_0_resize_req_0 <= cp_elements(294);
    cp_elements(295) <= cp_elements(216);
    cpelement_group_296 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(295) & cp_elements(304));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(296),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2543_final_reg_req_0 <= cp_elements(296);
    cp_elements(297) <= cp_elements(216);
    array_obj_ref_2543_base_resize_req_0 <= cp_elements(297);
    cp_elements(298) <= array_obj_ref_2543_index_0_resize_ack_0;
    array_obj_ref_2543_index_0_rename_req_0 <= cp_elements(298);
    cp_elements(299) <= array_obj_ref_2543_index_0_rename_ack_0;
    array_obj_ref_2543_offset_inst_req_0 <= cp_elements(299);
    cp_elements(300) <= array_obj_ref_2543_offset_inst_ack_0;
    cp_elements(301) <= array_obj_ref_2543_base_resize_ack_0;
    cpelement_group_302 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(300) & cp_elements(301));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(302),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2543_root_address_inst_req_0 <= cp_elements(302);
    cp_elements(303) <= array_obj_ref_2543_root_address_inst_ack_0;
    array_obj_ref_2543_root_address_inst_req_1 <= cp_elements(303);
    cp_elements(304) <= array_obj_ref_2543_root_address_inst_ack_1;
    cp_elements(305) <= array_obj_ref_2543_final_reg_ack_0;
    cpelement_group_306 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(305) & cp_elements(310));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(306),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2547_load_0_req_0 <= cp_elements(306);
    cp_elements(307) <= cp_elements(305);
    ptr_deref_2547_base_resize_req_0 <= cp_elements(307);
    cp_elements(308) <= ptr_deref_2547_base_resize_ack_0;
    ptr_deref_2547_root_address_inst_req_0 <= cp_elements(308);
    cp_elements(309) <= ptr_deref_2547_root_address_inst_ack_0;
    ptr_deref_2547_addr_0_req_0 <= cp_elements(309);
    cp_elements(310) <= ptr_deref_2547_addr_0_ack_0;
    cp_elements(311) <= ptr_deref_2547_load_0_ack_0;
    ptr_deref_2547_load_0_req_1 <= cp_elements(311);
    cp_elements(312) <= ptr_deref_2547_load_0_ack_1;
    ptr_deref_2547_gather_scatter_req_0 <= cp_elements(312);
    cp_elements(313) <= ptr_deref_2547_gather_scatter_ack_0;
    cpelement_group_314 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(315));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(314),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2551_inst_req_0 <= cp_elements(314);
    cp_elements(315) <= cp_elements(216);
    cp_elements(316) <= type_cast_2551_inst_ack_0;
    cpelement_group_317 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(316) & cp_elements(318));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(317),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2557_inst_req_0 <= cp_elements(317);
    cp_elements(318) <= cp_elements(216);
    cp_elements(319) <= binary_2557_inst_ack_0;
    binary_2557_inst_req_1 <= cp_elements(319);
    cp_elements(320) <= binary_2557_inst_ack_1;
    cpelement_group_321 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(322) & cp_elements(323));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(321),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2563_inst_req_0 <= cp_elements(321);
    cp_elements(322) <= cp_elements(216);
    cp_elements(323) <= cp_elements(231);
    cp_elements(324) <= binary_2563_inst_ack_0;
    binary_2563_inst_req_1 <= cp_elements(324);
    cp_elements(325) <= binary_2563_inst_ack_1;
    array_obj_ref_2567_index_0_resize_req_0 <= cp_elements(325);
    cp_elements(326) <= cp_elements(216);
    cpelement_group_327 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(326) & cp_elements(335));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(327),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2567_final_reg_req_0 <= cp_elements(327);
    cp_elements(328) <= cp_elements(216);
    array_obj_ref_2567_base_resize_req_0 <= cp_elements(328);
    cp_elements(329) <= array_obj_ref_2567_index_0_resize_ack_0;
    array_obj_ref_2567_index_0_rename_req_0 <= cp_elements(329);
    cp_elements(330) <= array_obj_ref_2567_index_0_rename_ack_0;
    array_obj_ref_2567_offset_inst_req_0 <= cp_elements(330);
    cp_elements(331) <= array_obj_ref_2567_offset_inst_ack_0;
    cp_elements(332) <= array_obj_ref_2567_base_resize_ack_0;
    cpelement_group_333 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(331) & cp_elements(332));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(333),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2567_root_address_inst_req_0 <= cp_elements(333);
    cp_elements(334) <= array_obj_ref_2567_root_address_inst_ack_0;
    array_obj_ref_2567_root_address_inst_req_1 <= cp_elements(334);
    cp_elements(335) <= array_obj_ref_2567_root_address_inst_ack_1;
    cp_elements(336) <= array_obj_ref_2567_final_reg_ack_0;
    cpelement_group_337 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(336) & cp_elements(341));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(337),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2571_load_0_req_0 <= cp_elements(337);
    cp_elements(338) <= cp_elements(336);
    ptr_deref_2571_base_resize_req_0 <= cp_elements(338);
    cp_elements(339) <= ptr_deref_2571_base_resize_ack_0;
    ptr_deref_2571_root_address_inst_req_0 <= cp_elements(339);
    cp_elements(340) <= ptr_deref_2571_root_address_inst_ack_0;
    ptr_deref_2571_addr_0_req_0 <= cp_elements(340);
    cp_elements(341) <= ptr_deref_2571_addr_0_ack_0;
    cp_elements(342) <= ptr_deref_2571_load_0_ack_0;
    ptr_deref_2571_load_0_req_1 <= cp_elements(342);
    cp_elements(343) <= ptr_deref_2571_load_0_ack_1;
    ptr_deref_2571_gather_scatter_req_0 <= cp_elements(343);
    cp_elements(344) <= ptr_deref_2571_gather_scatter_ack_0;
    cpelement_group_345 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(344) & cp_elements(346));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(345),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2575_inst_req_0 <= cp_elements(345);
    cp_elements(346) <= cp_elements(216);
    cp_elements(347) <= type_cast_2575_inst_ack_0;
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(349));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2581_inst_req_0 <= cp_elements(348);
    cp_elements(349) <= cp_elements(216);
    cp_elements(350) <= binary_2581_inst_ack_0;
    binary_2581_inst_req_1 <= cp_elements(350);
    cp_elements(351) <= binary_2581_inst_ack_1;
    cpelement_group_352 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(353) & cp_elements(354));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(352),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2587_inst_req_0 <= cp_elements(352);
    cp_elements(353) <= cp_elements(216);
    cp_elements(354) <= cp_elements(231);
    cp_elements(355) <= binary_2587_inst_ack_0;
    binary_2587_inst_req_1 <= cp_elements(355);
    cp_elements(356) <= binary_2587_inst_ack_1;
    array_obj_ref_2591_index_0_resize_req_0 <= cp_elements(356);
    cp_elements(357) <= cp_elements(216);
    cpelement_group_358 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(357) & cp_elements(366));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(358),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2591_final_reg_req_0 <= cp_elements(358);
    cp_elements(359) <= cp_elements(216);
    array_obj_ref_2591_base_resize_req_0 <= cp_elements(359);
    cp_elements(360) <= array_obj_ref_2591_index_0_resize_ack_0;
    array_obj_ref_2591_index_0_rename_req_0 <= cp_elements(360);
    cp_elements(361) <= array_obj_ref_2591_index_0_rename_ack_0;
    array_obj_ref_2591_offset_inst_req_0 <= cp_elements(361);
    cp_elements(362) <= array_obj_ref_2591_offset_inst_ack_0;
    cp_elements(363) <= array_obj_ref_2591_base_resize_ack_0;
    cpelement_group_364 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(362) & cp_elements(363));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2591_root_address_inst_req_0 <= cp_elements(364);
    cp_elements(365) <= array_obj_ref_2591_root_address_inst_ack_0;
    array_obj_ref_2591_root_address_inst_req_1 <= cp_elements(365);
    cp_elements(366) <= array_obj_ref_2591_root_address_inst_ack_1;
    cp_elements(367) <= array_obj_ref_2591_final_reg_ack_0;
    cpelement_group_368 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(367) & cp_elements(372));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(368),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2595_load_0_req_0 <= cp_elements(368);
    cp_elements(369) <= cp_elements(367);
    ptr_deref_2595_base_resize_req_0 <= cp_elements(369);
    cp_elements(370) <= ptr_deref_2595_base_resize_ack_0;
    ptr_deref_2595_root_address_inst_req_0 <= cp_elements(370);
    cp_elements(371) <= ptr_deref_2595_root_address_inst_ack_0;
    ptr_deref_2595_addr_0_req_0 <= cp_elements(371);
    cp_elements(372) <= ptr_deref_2595_addr_0_ack_0;
    cp_elements(373) <= ptr_deref_2595_load_0_ack_0;
    ptr_deref_2595_load_0_req_1 <= cp_elements(373);
    cp_elements(374) <= ptr_deref_2595_load_0_ack_1;
    ptr_deref_2595_gather_scatter_req_0 <= cp_elements(374);
    cp_elements(375) <= ptr_deref_2595_gather_scatter_ack_0;
    cpelement_group_376 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(375) & cp_elements(377));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(376),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2599_inst_req_0 <= cp_elements(376);
    cp_elements(377) <= cp_elements(216);
    cp_elements(378) <= type_cast_2599_inst_ack_0;
    cpelement_group_379 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(378) & cp_elements(380));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(379),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2605_inst_req_0 <= cp_elements(379);
    cp_elements(380) <= cp_elements(216);
    cp_elements(381) <= binary_2605_inst_ack_0;
    binary_2605_inst_req_1 <= cp_elements(381);
    cp_elements(382) <= binary_2605_inst_ack_1;
    cpelement_group_383 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(384) & cp_elements(385));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(383),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2611_inst_req_0 <= cp_elements(383);
    cp_elements(384) <= cp_elements(216);
    cp_elements(385) <= cp_elements(231);
    cp_elements(386) <= binary_2611_inst_ack_0;
    binary_2611_inst_req_1 <= cp_elements(386);
    cp_elements(387) <= binary_2611_inst_ack_1;
    array_obj_ref_2615_index_0_resize_req_0 <= cp_elements(387);
    cp_elements(388) <= cp_elements(216);
    cpelement_group_389 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(388) & cp_elements(397));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(389),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2615_final_reg_req_0 <= cp_elements(389);
    cp_elements(390) <= cp_elements(216);
    array_obj_ref_2615_base_resize_req_0 <= cp_elements(390);
    cp_elements(391) <= array_obj_ref_2615_index_0_resize_ack_0;
    array_obj_ref_2615_index_0_rename_req_0 <= cp_elements(391);
    cp_elements(392) <= array_obj_ref_2615_index_0_rename_ack_0;
    array_obj_ref_2615_offset_inst_req_0 <= cp_elements(392);
    cp_elements(393) <= array_obj_ref_2615_offset_inst_ack_0;
    cp_elements(394) <= array_obj_ref_2615_base_resize_ack_0;
    cpelement_group_395 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(393) & cp_elements(394));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(395),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2615_root_address_inst_req_0 <= cp_elements(395);
    cp_elements(396) <= array_obj_ref_2615_root_address_inst_ack_0;
    array_obj_ref_2615_root_address_inst_req_1 <= cp_elements(396);
    cp_elements(397) <= array_obj_ref_2615_root_address_inst_ack_1;
    cp_elements(398) <= array_obj_ref_2615_final_reg_ack_0;
    cpelement_group_399 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(398) & cp_elements(403));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(399),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2619_load_0_req_0 <= cp_elements(399);
    cp_elements(400) <= cp_elements(398);
    ptr_deref_2619_base_resize_req_0 <= cp_elements(400);
    cp_elements(401) <= ptr_deref_2619_base_resize_ack_0;
    ptr_deref_2619_root_address_inst_req_0 <= cp_elements(401);
    cp_elements(402) <= ptr_deref_2619_root_address_inst_ack_0;
    ptr_deref_2619_addr_0_req_0 <= cp_elements(402);
    cp_elements(403) <= ptr_deref_2619_addr_0_ack_0;
    cp_elements(404) <= ptr_deref_2619_load_0_ack_0;
    ptr_deref_2619_load_0_req_1 <= cp_elements(404);
    cp_elements(405) <= ptr_deref_2619_load_0_ack_1;
    ptr_deref_2619_gather_scatter_req_0 <= cp_elements(405);
    cp_elements(406) <= ptr_deref_2619_gather_scatter_ack_0;
    cpelement_group_407 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(406) & cp_elements(408));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(407),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2623_inst_req_0 <= cp_elements(407);
    cp_elements(408) <= cp_elements(216);
    cp_elements(409) <= type_cast_2623_inst_ack_0;
    cpelement_group_410 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(409) & cp_elements(411));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(410),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2629_inst_req_0 <= cp_elements(410);
    cp_elements(411) <= cp_elements(216);
    cp_elements(412) <= binary_2629_inst_ack_0;
    binary_2629_inst_req_1 <= cp_elements(412);
    cp_elements(413) <= binary_2629_inst_ack_1;
    cpelement_group_414 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(415) & cp_elements(416));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(414),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2635_inst_req_0 <= cp_elements(414);
    cp_elements(415) <= cp_elements(216);
    cp_elements(416) <= cp_elements(231);
    cp_elements(417) <= binary_2635_inst_ack_0;
    binary_2635_inst_req_1 <= cp_elements(417);
    cp_elements(418) <= binary_2635_inst_ack_1;
    array_obj_ref_2639_index_0_resize_req_0 <= cp_elements(418);
    cp_elements(419) <= cp_elements(216);
    cpelement_group_420 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(419) & cp_elements(428));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(420),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2639_final_reg_req_0 <= cp_elements(420);
    cp_elements(421) <= cp_elements(216);
    array_obj_ref_2639_base_resize_req_0 <= cp_elements(421);
    cp_elements(422) <= array_obj_ref_2639_index_0_resize_ack_0;
    array_obj_ref_2639_index_0_rename_req_0 <= cp_elements(422);
    cp_elements(423) <= array_obj_ref_2639_index_0_rename_ack_0;
    array_obj_ref_2639_offset_inst_req_0 <= cp_elements(423);
    cp_elements(424) <= array_obj_ref_2639_offset_inst_ack_0;
    cp_elements(425) <= array_obj_ref_2639_base_resize_ack_0;
    cpelement_group_426 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(424) & cp_elements(425));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(426),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2639_root_address_inst_req_0 <= cp_elements(426);
    cp_elements(427) <= array_obj_ref_2639_root_address_inst_ack_0;
    array_obj_ref_2639_root_address_inst_req_1 <= cp_elements(427);
    cp_elements(428) <= array_obj_ref_2639_root_address_inst_ack_1;
    cp_elements(429) <= array_obj_ref_2639_final_reg_ack_0;
    cpelement_group_430 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(429) & cp_elements(434));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(430),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2643_load_0_req_0 <= cp_elements(430);
    cp_elements(431) <= cp_elements(429);
    ptr_deref_2643_base_resize_req_0 <= cp_elements(431);
    cp_elements(432) <= ptr_deref_2643_base_resize_ack_0;
    ptr_deref_2643_root_address_inst_req_0 <= cp_elements(432);
    cp_elements(433) <= ptr_deref_2643_root_address_inst_ack_0;
    ptr_deref_2643_addr_0_req_0 <= cp_elements(433);
    cp_elements(434) <= ptr_deref_2643_addr_0_ack_0;
    cp_elements(435) <= ptr_deref_2643_load_0_ack_0;
    ptr_deref_2643_load_0_req_1 <= cp_elements(435);
    cp_elements(436) <= ptr_deref_2643_load_0_ack_1;
    ptr_deref_2643_gather_scatter_req_0 <= cp_elements(436);
    cp_elements(437) <= ptr_deref_2643_gather_scatter_ack_0;
    cpelement_group_438 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(437) & cp_elements(439));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(438),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2647_inst_req_0 <= cp_elements(438);
    cp_elements(439) <= cp_elements(216);
    cp_elements(440) <= type_cast_2647_inst_ack_0;
    cpelement_group_441 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(440) & cp_elements(442));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(441),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2653_inst_req_0 <= cp_elements(441);
    cp_elements(442) <= cp_elements(216);
    cp_elements(443) <= binary_2653_inst_ack_0;
    binary_2653_inst_req_1 <= cp_elements(443);
    cp_elements(444) <= binary_2653_inst_ack_1;
    cp_elements(445) <= cp_elements(216);
    cpelement_group_446 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(445) & cp_elements(455));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(446),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2657_final_reg_req_0 <= cp_elements(446);
    cp_elements(447) <= cp_elements(216);
    array_obj_ref_2657_base_resize_req_0 <= cp_elements(447);
    cp_elements(448) <= cp_elements(231);
    array_obj_ref_2657_index_0_resize_req_0 <= cp_elements(448);
    cp_elements(449) <= array_obj_ref_2657_index_0_resize_ack_0;
    array_obj_ref_2657_index_0_rename_req_0 <= cp_elements(449);
    cp_elements(450) <= array_obj_ref_2657_index_0_rename_ack_0;
    array_obj_ref_2657_offset_inst_req_0 <= cp_elements(450);
    cp_elements(451) <= array_obj_ref_2657_offset_inst_ack_0;
    cp_elements(452) <= array_obj_ref_2657_base_resize_ack_0;
    cpelement_group_453 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(451) & cp_elements(452));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(453),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2657_root_address_inst_req_0 <= cp_elements(453);
    cp_elements(454) <= array_obj_ref_2657_root_address_inst_ack_0;
    array_obj_ref_2657_root_address_inst_req_1 <= cp_elements(454);
    cp_elements(455) <= array_obj_ref_2657_root_address_inst_ack_1;
    cp_elements(456) <= array_obj_ref_2657_final_reg_ack_0;
    cpelement_group_457 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(456) & cp_elements(461));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(457),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2661_load_0_req_0 <= cp_elements(457);
    cp_elements(458) <= cp_elements(456);
    ptr_deref_2661_base_resize_req_0 <= cp_elements(458);
    cp_elements(459) <= ptr_deref_2661_base_resize_ack_0;
    ptr_deref_2661_root_address_inst_req_0 <= cp_elements(459);
    cp_elements(460) <= ptr_deref_2661_root_address_inst_ack_0;
    ptr_deref_2661_addr_0_req_0 <= cp_elements(460);
    cp_elements(461) <= ptr_deref_2661_addr_0_ack_0;
    cp_elements(462) <= ptr_deref_2661_load_0_ack_0;
    ptr_deref_2661_load_0_req_1 <= cp_elements(462);
    cp_elements(463) <= ptr_deref_2661_load_0_ack_1;
    ptr_deref_2661_gather_scatter_req_0 <= cp_elements(463);
    cp_elements(464) <= ptr_deref_2661_gather_scatter_ack_0;
    cpelement_group_465 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(464) & cp_elements(466));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(465),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2665_inst_req_0 <= cp_elements(465);
    cp_elements(466) <= cp_elements(216);
    cp_elements(467) <= type_cast_2665_inst_ack_0;
    cpelement_group_468 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(467) & cp_elements(469));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(468),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2671_inst_req_0 <= cp_elements(468);
    cp_elements(469) <= cp_elements(216);
    cp_elements(470) <= binary_2671_inst_ack_0;
    binary_2671_inst_req_1 <= cp_elements(470);
    cp_elements(471) <= binary_2671_inst_ack_1;
    cpelement_group_472 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(258) & cp_elements(289) & cp_elements(473));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(472),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2676_inst_req_0 <= cp_elements(472);
    cp_elements(473) <= cp_elements(216);
    cp_elements(474) <= binary_2676_inst_ack_0;
    binary_2676_inst_req_1 <= cp_elements(474);
    cp_elements(475) <= binary_2676_inst_ack_1;
    cpelement_group_476 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(320) & cp_elements(475) & cp_elements(477));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(476),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2681_inst_req_0 <= cp_elements(476);
    cp_elements(477) <= cp_elements(216);
    cp_elements(478) <= binary_2681_inst_ack_0;
    binary_2681_inst_req_1 <= cp_elements(478);
    cp_elements(479) <= binary_2681_inst_ack_1;
    cpelement_group_480 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(351) & cp_elements(479) & cp_elements(481));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(480),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2686_inst_req_0 <= cp_elements(480);
    cp_elements(481) <= cp_elements(216);
    cp_elements(482) <= binary_2686_inst_ack_0;
    binary_2686_inst_req_1 <= cp_elements(482);
    cp_elements(483) <= binary_2686_inst_ack_1;
    cpelement_group_484 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(382) & cp_elements(483) & cp_elements(485));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(484),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2691_inst_req_0 <= cp_elements(484);
    cp_elements(485) <= cp_elements(216);
    cp_elements(486) <= binary_2691_inst_ack_0;
    binary_2691_inst_req_1 <= cp_elements(486);
    cp_elements(487) <= binary_2691_inst_ack_1;
    cpelement_group_488 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(413) & cp_elements(487) & cp_elements(489));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(488),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2696_inst_req_0 <= cp_elements(488);
    cp_elements(489) <= cp_elements(216);
    cp_elements(490) <= binary_2696_inst_ack_0;
    binary_2696_inst_req_1 <= cp_elements(490);
    cp_elements(491) <= binary_2696_inst_ack_1;
    cpelement_group_492 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(444) & cp_elements(491) & cp_elements(493));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(492),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2701_inst_req_0 <= cp_elements(492);
    cp_elements(493) <= cp_elements(216);
    cp_elements(494) <= binary_2701_inst_ack_0;
    binary_2701_inst_req_1 <= cp_elements(494);
    cp_elements(495) <= binary_2701_inst_ack_1;
    cpelement_group_496 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(471) & cp_elements(495) & cp_elements(497));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(496),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2706_inst_req_0 <= cp_elements(496);
    cp_elements(497) <= cp_elements(216);
    cp_elements(498) <= binary_2706_inst_ack_0;
    binary_2706_inst_req_1 <= cp_elements(498);
    cp_elements(499) <= binary_2706_inst_ack_1;
    cpelement_group_500 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(226) & cp_elements(499));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(500),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(501) <= cp_elements(2);
    cp_elements(502) <= false;
    cp_elements(503) <= cp_elements(502);
    cp_elements(504) <= cp_elements(2);
    if_stmt_2714_branch_req_0 <= cp_elements(504);
    cp_elements(505) <= cp_elements(504);
    cp_elements(506) <= cp_elements(505);
    cp_elements(507) <= if_stmt_2714_branch_ack_1;
    cp_elements(508) <= cp_elements(505);
    cp_elements(509) <= if_stmt_2714_branch_ack_0;
    simple_obj_ref_2742_inst_req_0 <= cp_elements(509);
    cp_elements(510) <= simple_obj_ref_2721_inst_ack_0;
    simple_obj_ref_2731_inst_req_0 <= cp_elements(510);
    cp_elements(511) <= simple_obj_ref_2731_inst_ack_0;
    cp_elements(512) <= cp_elements(511);
    cpelement_group_513 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(514) & cp_elements(515));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(513),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2738_inst_req_0 <= cp_elements(513);
    cp_elements(514) <= cp_elements(512);
    cp_elements(515) <= cp_elements(512);
    cp_elements(516) <= binary_2738_inst_ack_0;
    binary_2738_inst_req_1 <= cp_elements(516);
    cp_elements(517) <= binary_2738_inst_ack_1;
    type_cast_2473_inst_req_0 <= cp_elements(517);
    cp_elements(518) <= simple_obj_ref_2742_inst_ack_0;
    simple_obj_ref_2751_inst_req_0 <= cp_elements(518);
    cp_elements(519) <= simple_obj_ref_2751_inst_ack_0;
    simple_obj_ref_2760_inst_req_0 <= cp_elements(519);
    cp_elements(520) <= simple_obj_ref_2760_inst_ack_0;
    simple_obj_ref_2770_inst_req_0 <= cp_elements(520);
    cp_elements(521) <= simple_obj_ref_2770_inst_ack_0;
    cp_elements(522) <= OrReduce(cp_elements(4) & cp_elements(521));
    cp_elements(523) <= cp_elements(522);
    simple_obj_ref_2242_inst_req_0 <= cp_elements(523);
    cp_elements(524) <= type_cast_2473_inst_ack_0;
    phi_stmt_2469_req_0 <= cp_elements(524);
    cp_elements(525) <= OrReduce(cp_elements(215) & cp_elements(524));
    cp_elements(526) <= cp_elements(525);
    cp_elements(527) <= phi_stmt_2469_ack_0;
    cp_elements(528) <= false;
    cp_elements(529) <= cp_elements(528);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2269_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2269_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2269_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2282_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2282_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2282_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2301_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2301_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2301_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2320_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2320_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2320_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2339_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2339_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2339_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2358_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2358_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2358_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2391_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2391_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2391_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2501_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2501_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2501_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2501_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2519_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2519_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2519_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2519_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2543_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2543_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2543_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2543_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2567_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2567_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2567_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2567_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2591_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2591_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2591_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2591_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2615_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2615_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2615_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2615_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2639_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2639_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2639_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2639_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2657_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2657_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2657_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2657_root_address : std_logic_vector(10 downto 0);
    signal iNsTr_0_2229 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2713 : std_logic_vector(31 downto 0);
    signal iNsTr_13_2730 : std_logic_vector(31 downto 0);
    signal iNsTr_17_2750 : std_logic_vector(31 downto 0);
    signal iNsTr_19_2759 : std_logic_vector(31 downto 0);
    signal iNsTr_21_2769 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2240 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2253 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2262 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2447 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2457 : std_logic_vector(31 downto 0);
    signal indvar_2469 : std_logic_vector(15 downto 0);
    signal ins38_2441 : std_logic_vector(63 downto 0);
    signal ins77_2707 : std_logic_vector(63 downto 0);
    signal mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_2411 : std_logic_vector(63 downto 0);
    signal mask17x_xmaskedx_xmaskedx_xmasked_2416 : std_logic_vector(63 downto 0);
    signal mask22x_xmaskedx_xmaskedx_xmasked_2421 : std_logic_vector(63 downto 0);
    signal mask27x_xmaskedx_xmasked_2426 : std_logic_vector(63 downto 0);
    signal mask32x_xmasked_2431 : std_logic_vector(63 downto 0);
    signal mask37_2436 : std_logic_vector(63 downto 0);
    signal mask51_2677 : std_logic_vector(63 downto 0);
    signal mask56_2682 : std_logic_vector(63 downto 0);
    signal mask61x_xmaskedx_xmasked_2687 : std_logic_vector(63 downto 0);
    signal mask66x_xmaskedx_xmasked_2692 : std_logic_vector(63 downto 0);
    signal mask71x_xmasked_2697 : std_logic_vector(63 downto 0);
    signal mask76_2702 : std_logic_vector(63 downto 0);
    signal phitmp_2739 : std_logic_vector(15 downto 0);
    signal ptr_deref_2273_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2273_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2273_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2273_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2273_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2286_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2286_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2286_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2286_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2286_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2305_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2305_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2305_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2305_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2305_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2324_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2324_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2324_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2324_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2324_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2343_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2343_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2343_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2343_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2343_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2362_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2362_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2362_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2362_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2362_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2376_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2376_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2376_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2376_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2376_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2395_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2395_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2395_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2395_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2395_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2505_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2505_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2505_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2505_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2505_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2523_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2523_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2523_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2523_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2523_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2547_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2547_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2547_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2547_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2547_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2571_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2571_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2571_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2571_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2571_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2595_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2595_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2595_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2595_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2595_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2619_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2619_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2619_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2619_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2619_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2643_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2643_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2643_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2643_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2643_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2661_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2661_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2661_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2661_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2661_word_offset_0 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2500_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2500_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2518_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2518_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2542_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2542_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2566_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2566_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2590_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2590_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2614_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2614_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2638_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2638_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2656_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2656_scaled : std_logic_vector(10 downto 0);
    signal tmp10_2310 : std_logic_vector(63 downto 0);
    signal tmp11_2316 : std_logic_vector(63 downto 0);
    signal tmp124_2243 : std_logic_vector(31 downto 0);
    signal tmp125_2247 : std_logic_vector(31 downto 0);
    signal tmp126_2256 : std_logic_vector(31 downto 0);
    signal tmp127_2265 : std_logic_vector(7 downto 0);
    signal tmp128_2270 : std_logic_vector(31 downto 0);
    signal tmp129_2274 : std_logic_vector(7 downto 0);
    signal tmp130_2283 : std_logic_vector(31 downto 0);
    signal tmp131_2287 : std_logic_vector(7 downto 0);
    signal tmp132_2302 : std_logic_vector(31 downto 0);
    signal tmp133_2306 : std_logic_vector(7 downto 0);
    signal tmp134_2321 : std_logic_vector(31 downto 0);
    signal tmp135_2325 : std_logic_vector(7 downto 0);
    signal tmp136_2340 : std_logic_vector(31 downto 0);
    signal tmp137_2344 : std_logic_vector(7 downto 0);
    signal tmp138_2359 : std_logic_vector(31 downto 0);
    signal tmp139_2363 : std_logic_vector(7 downto 0);
    signal tmp140_2377 : std_logic_vector(7 downto 0);
    signal tmp141_2392 : std_logic_vector(31 downto 0);
    signal tmp142_2396 : std_logic_vector(7 downto 0);
    signal tmp144_2481 : std_logic_vector(31 downto 0);
    signal tmp145_2466 : std_logic_vector(31 downto 0);
    signal tmp146_2486 : std_logic_vector(0 downto 0);
    signal tmp149_2492 : std_logic_vector(31 downto 0);
    signal tmp150_2498 : std_logic_vector(31 downto 0);
    signal tmp151_2502 : std_logic_vector(31 downto 0);
    signal tmp152_2506 : std_logic_vector(7 downto 0);
    signal tmp155_2516 : std_logic_vector(31 downto 0);
    signal tmp156_2520 : std_logic_vector(31 downto 0);
    signal tmp157_2524 : std_logic_vector(7 downto 0);
    signal tmp15_2329 : std_logic_vector(63 downto 0);
    signal tmp160_2540 : std_logic_vector(31 downto 0);
    signal tmp161_2544 : std_logic_vector(31 downto 0);
    signal tmp162_2548 : std_logic_vector(7 downto 0);
    signal tmp165_2564 : std_logic_vector(31 downto 0);
    signal tmp166_2568 : std_logic_vector(31 downto 0);
    signal tmp167_2572 : std_logic_vector(7 downto 0);
    signal tmp16_2335 : std_logic_vector(63 downto 0);
    signal tmp170_2588 : std_logic_vector(31 downto 0);
    signal tmp171_2592 : std_logic_vector(31 downto 0);
    signal tmp172_2596 : std_logic_vector(7 downto 0);
    signal tmp175_2612 : std_logic_vector(31 downto 0);
    signal tmp176_2616 : std_logic_vector(31 downto 0);
    signal tmp177_2620 : std_logic_vector(7 downto 0);
    signal tmp180_2636 : std_logic_vector(31 downto 0);
    signal tmp181_2640 : std_logic_vector(31 downto 0);
    signal tmp182_2644 : std_logic_vector(7 downto 0);
    signal tmp185_2658 : std_logic_vector(31 downto 0);
    signal tmp186_2662 : std_logic_vector(7 downto 0);
    signal tmp20_2348 : std_logic_vector(63 downto 0);
    signal tmp21_2354 : std_logic_vector(63 downto 0);
    signal tmp25_2367 : std_logic_vector(63 downto 0);
    signal tmp26_2373 : std_logic_vector(63 downto 0);
    signal tmp30_2381 : std_logic_vector(63 downto 0);
    signal tmp31_2387 : std_logic_vector(63 downto 0);
    signal tmp35_2400 : std_logic_vector(63 downto 0);
    signal tmp36_2406 : std_logic_vector(63 downto 0);
    signal tmp3_2278 : std_logic_vector(63 downto 0);
    signal tmp40_2510 : std_logic_vector(63 downto 0);
    signal tmp44_2528 : std_logic_vector(63 downto 0);
    signal tmp45_2534 : std_logic_vector(63 downto 0);
    signal tmp49_2552 : std_logic_vector(63 downto 0);
    signal tmp50_2558 : std_logic_vector(63 downto 0);
    signal tmp54_2576 : std_logic_vector(63 downto 0);
    signal tmp55_2582 : std_logic_vector(63 downto 0);
    signal tmp59_2600 : std_logic_vector(63 downto 0);
    signal tmp5_2291 : std_logic_vector(63 downto 0);
    signal tmp60_2606 : std_logic_vector(63 downto 0);
    signal tmp64_2624 : std_logic_vector(63 downto 0);
    signal tmp65_2630 : std_logic_vector(63 downto 0);
    signal tmp69_2648 : std_logic_vector(63 downto 0);
    signal tmp6_2297 : std_logic_vector(63 downto 0);
    signal tmp70_2654 : std_logic_vector(63 downto 0);
    signal tmp74_2666 : std_logic_vector(63 downto 0);
    signal tmp75_2672 : std_logic_vector(63 downto 0);
    signal tmp_2232 : std_logic_vector(7 downto 0);
    signal type_cast_2295_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2314_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2333_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2352_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2371_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2385_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2404_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2450_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2464_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2473_wire : std_logic_vector(15 downto 0);
    signal type_cast_2476_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2490_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2496_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2514_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2538_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2556_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2562_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2580_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2586_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2604_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2610_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2628_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2634_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2652_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2670_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2723_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2737_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2762_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_2269_final_offset <= "00000000111";
    array_obj_ref_2282_final_offset <= "00000000110";
    array_obj_ref_2301_final_offset <= "00000000101";
    array_obj_ref_2320_final_offset <= "00000000100";
    array_obj_ref_2339_final_offset <= "00000000011";
    array_obj_ref_2358_final_offset <= "00000000010";
    array_obj_ref_2391_final_offset <= "00000000001";
    array_obj_ref_2501_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2519_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2543_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2567_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2591_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2615_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2639_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2657_offset_scale_factor_0 <= "00000000001";
    iNsTr_0_2229 <= "00000000000000000000000000000000";
    iNsTr_10_2713 <= "00000000000000000000000000000000";
    iNsTr_13_2730 <= "00000000000000000000000000000000";
    iNsTr_17_2750 <= "00000000000000000000000000000000";
    iNsTr_19_2759 <= "00000000000000000000000000000000";
    iNsTr_21_2769 <= "00000000000000000000000000000000";
    iNsTr_2_2240 <= "00000000000000000000000000000000";
    iNsTr_3_2253 <= "00000000000000000000000000000000";
    iNsTr_4_2262 <= "00000000000000000000000000000000";
    iNsTr_5_2447 <= "00000000000000000000000000000000";
    iNsTr_7_2457 <= "00000000000000000000000000000000";
    ptr_deref_2273_word_offset_0 <= "00000000000";
    ptr_deref_2286_word_offset_0 <= "00000000000";
    ptr_deref_2305_word_offset_0 <= "00000000000";
    ptr_deref_2324_word_offset_0 <= "00000000000";
    ptr_deref_2343_word_offset_0 <= "00000000000";
    ptr_deref_2362_word_offset_0 <= "00000000000";
    ptr_deref_2376_word_offset_0 <= "00000000000";
    ptr_deref_2395_word_offset_0 <= "00000000000";
    ptr_deref_2505_word_offset_0 <= "00000000000";
    ptr_deref_2523_word_offset_0 <= "00000000000";
    ptr_deref_2547_word_offset_0 <= "00000000000";
    ptr_deref_2571_word_offset_0 <= "00000000000";
    ptr_deref_2595_word_offset_0 <= "00000000000";
    ptr_deref_2619_word_offset_0 <= "00000000000";
    ptr_deref_2643_word_offset_0 <= "00000000000";
    ptr_deref_2661_word_offset_0 <= "00000000000";
    type_cast_2295_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2314_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2352_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2371_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2385_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2404_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2450_wire_constant <= "11111111";
    type_cast_2464_wire_constant <= "11111111111111111111111111111111";
    type_cast_2476_wire_constant <= "0000000000000001";
    type_cast_2490_wire_constant <= "00000000000000000000000000000011";
    type_cast_2496_wire_constant <= "00000000000000000000000000000111";
    type_cast_2514_wire_constant <= "00000000000000000000000000000110";
    type_cast_2532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2538_wire_constant <= "00000000000000000000000000000101";
    type_cast_2556_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2562_wire_constant <= "00000000000000000000000000000100";
    type_cast_2580_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2586_wire_constant <= "00000000000000000000000000000011";
    type_cast_2604_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2610_wire_constant <= "00000000000000000000000000000010";
    type_cast_2628_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2634_wire_constant <= "00000000000000000000000000000001";
    type_cast_2652_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2670_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2723_wire_constant <= "00000000";
    type_cast_2737_wire_constant <= "0000000000000001";
    type_cast_2762_wire_constant <= "00000001";
    phi_stmt_2469: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2473_wire & type_cast_2476_wire_constant;
      req <= phi_stmt_2469_req_0 & phi_stmt_2469_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2469_ack_0,
          idata => idata,
          odata => indvar_2469,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2469
    array_obj_ref_2269_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2269_resized_base_address, req => array_obj_ref_2269_base_resize_req_0, ack => array_obj_ref_2269_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2269_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2269_root_address, dout => tmp128_2270, req => array_obj_ref_2269_final_reg_req_0, ack => array_obj_ref_2269_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2282_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2282_resized_base_address, req => array_obj_ref_2282_base_resize_req_0, ack => array_obj_ref_2282_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2282_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2282_root_address, dout => tmp130_2283, req => array_obj_ref_2282_final_reg_req_0, ack => array_obj_ref_2282_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2301_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2301_resized_base_address, req => array_obj_ref_2301_base_resize_req_0, ack => array_obj_ref_2301_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2301_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2301_root_address, dout => tmp132_2302, req => array_obj_ref_2301_final_reg_req_0, ack => array_obj_ref_2301_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2320_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2320_resized_base_address, req => array_obj_ref_2320_base_resize_req_0, ack => array_obj_ref_2320_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2320_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2320_root_address, dout => tmp134_2321, req => array_obj_ref_2320_final_reg_req_0, ack => array_obj_ref_2320_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2339_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2339_resized_base_address, req => array_obj_ref_2339_base_resize_req_0, ack => array_obj_ref_2339_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2339_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2339_root_address, dout => tmp136_2340, req => array_obj_ref_2339_final_reg_req_0, ack => array_obj_ref_2339_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2358_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2358_resized_base_address, req => array_obj_ref_2358_base_resize_req_0, ack => array_obj_ref_2358_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2358_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2358_root_address, dout => tmp138_2359, req => array_obj_ref_2358_final_reg_req_0, ack => array_obj_ref_2358_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2391_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2391_resized_base_address, req => array_obj_ref_2391_base_resize_req_0, ack => array_obj_ref_2391_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2391_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2391_root_address, dout => tmp141_2392, req => array_obj_ref_2391_final_reg_req_0, ack => array_obj_ref_2391_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2501_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2501_resized_base_address, req => array_obj_ref_2501_base_resize_req_0, ack => array_obj_ref_2501_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2501_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2501_root_address, dout => tmp151_2502, req => array_obj_ref_2501_final_reg_req_0, ack => array_obj_ref_2501_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2501_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp150_2498, dout => simple_obj_ref_2500_resized, req => array_obj_ref_2501_index_0_resize_req_0, ack => array_obj_ref_2501_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2501_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2500_scaled, dout => array_obj_ref_2501_final_offset, req => array_obj_ref_2501_offset_inst_req_0, ack => array_obj_ref_2501_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2519_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2519_resized_base_address, req => array_obj_ref_2519_base_resize_req_0, ack => array_obj_ref_2519_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2519_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2519_root_address, dout => tmp156_2520, req => array_obj_ref_2519_final_reg_req_0, ack => array_obj_ref_2519_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2519_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp155_2516, dout => simple_obj_ref_2518_resized, req => array_obj_ref_2519_index_0_resize_req_0, ack => array_obj_ref_2519_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2519_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2518_scaled, dout => array_obj_ref_2519_final_offset, req => array_obj_ref_2519_offset_inst_req_0, ack => array_obj_ref_2519_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2543_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2543_resized_base_address, req => array_obj_ref_2543_base_resize_req_0, ack => array_obj_ref_2543_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2543_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2543_root_address, dout => tmp161_2544, req => array_obj_ref_2543_final_reg_req_0, ack => array_obj_ref_2543_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2543_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp160_2540, dout => simple_obj_ref_2542_resized, req => array_obj_ref_2543_index_0_resize_req_0, ack => array_obj_ref_2543_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2543_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2542_scaled, dout => array_obj_ref_2543_final_offset, req => array_obj_ref_2543_offset_inst_req_0, ack => array_obj_ref_2543_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2567_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2567_resized_base_address, req => array_obj_ref_2567_base_resize_req_0, ack => array_obj_ref_2567_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2567_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2567_root_address, dout => tmp166_2568, req => array_obj_ref_2567_final_reg_req_0, ack => array_obj_ref_2567_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2567_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp165_2564, dout => simple_obj_ref_2566_resized, req => array_obj_ref_2567_index_0_resize_req_0, ack => array_obj_ref_2567_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2567_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2566_scaled, dout => array_obj_ref_2567_final_offset, req => array_obj_ref_2567_offset_inst_req_0, ack => array_obj_ref_2567_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2591_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2591_resized_base_address, req => array_obj_ref_2591_base_resize_req_0, ack => array_obj_ref_2591_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2591_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2591_root_address, dout => tmp171_2592, req => array_obj_ref_2591_final_reg_req_0, ack => array_obj_ref_2591_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2591_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp170_2588, dout => simple_obj_ref_2590_resized, req => array_obj_ref_2591_index_0_resize_req_0, ack => array_obj_ref_2591_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2591_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2590_scaled, dout => array_obj_ref_2591_final_offset, req => array_obj_ref_2591_offset_inst_req_0, ack => array_obj_ref_2591_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2615_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2615_resized_base_address, req => array_obj_ref_2615_base_resize_req_0, ack => array_obj_ref_2615_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2615_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2615_root_address, dout => tmp176_2616, req => array_obj_ref_2615_final_reg_req_0, ack => array_obj_ref_2615_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2615_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp175_2612, dout => simple_obj_ref_2614_resized, req => array_obj_ref_2615_index_0_resize_req_0, ack => array_obj_ref_2615_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2615_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2614_scaled, dout => array_obj_ref_2615_final_offset, req => array_obj_ref_2615_offset_inst_req_0, ack => array_obj_ref_2615_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2639_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2639_resized_base_address, req => array_obj_ref_2639_base_resize_req_0, ack => array_obj_ref_2639_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2639_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2639_root_address, dout => tmp181_2640, req => array_obj_ref_2639_final_reg_req_0, ack => array_obj_ref_2639_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2639_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp180_2636, dout => simple_obj_ref_2638_resized, req => array_obj_ref_2639_index_0_resize_req_0, ack => array_obj_ref_2639_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2639_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2638_scaled, dout => array_obj_ref_2639_final_offset, req => array_obj_ref_2639_offset_inst_req_0, ack => array_obj_ref_2639_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2657_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => array_obj_ref_2657_resized_base_address, req => array_obj_ref_2657_base_resize_req_0, ack => array_obj_ref_2657_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2657_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2657_root_address, dout => tmp185_2658, req => array_obj_ref_2657_final_reg_req_0, ack => array_obj_ref_2657_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2657_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp149_2492, dout => simple_obj_ref_2656_resized, req => array_obj_ref_2657_index_0_resize_req_0, ack => array_obj_ref_2657_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2657_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2656_scaled, dout => array_obj_ref_2657_final_offset, req => array_obj_ref_2657_offset_inst_req_0, ack => array_obj_ref_2657_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2273_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp128_2270, dout => ptr_deref_2273_resized_base_address, req => ptr_deref_2273_base_resize_req_0, ack => ptr_deref_2273_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2286_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp130_2283, dout => ptr_deref_2286_resized_base_address, req => ptr_deref_2286_base_resize_req_0, ack => ptr_deref_2286_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2305_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp132_2302, dout => ptr_deref_2305_resized_base_address, req => ptr_deref_2305_base_resize_req_0, ack => ptr_deref_2305_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2324_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp134_2321, dout => ptr_deref_2324_resized_base_address, req => ptr_deref_2324_base_resize_req_0, ack => ptr_deref_2324_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2343_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp136_2340, dout => ptr_deref_2343_resized_base_address, req => ptr_deref_2343_base_resize_req_0, ack => ptr_deref_2343_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2362_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp138_2359, dout => ptr_deref_2362_resized_base_address, req => ptr_deref_2362_base_resize_req_0, ack => ptr_deref_2362_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2376_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_2247, dout => ptr_deref_2376_resized_base_address, req => ptr_deref_2376_base_resize_req_0, ack => ptr_deref_2376_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2395_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp141_2392, dout => ptr_deref_2395_resized_base_address, req => ptr_deref_2395_base_resize_req_0, ack => ptr_deref_2395_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2505_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp151_2502, dout => ptr_deref_2505_resized_base_address, req => ptr_deref_2505_base_resize_req_0, ack => ptr_deref_2505_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2523_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp156_2520, dout => ptr_deref_2523_resized_base_address, req => ptr_deref_2523_base_resize_req_0, ack => ptr_deref_2523_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2547_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp161_2544, dout => ptr_deref_2547_resized_base_address, req => ptr_deref_2547_base_resize_req_0, ack => ptr_deref_2547_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2571_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp166_2568, dout => ptr_deref_2571_resized_base_address, req => ptr_deref_2571_base_resize_req_0, ack => ptr_deref_2571_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2595_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp171_2592, dout => ptr_deref_2595_resized_base_address, req => ptr_deref_2595_base_resize_req_0, ack => ptr_deref_2595_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2619_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp176_2616, dout => ptr_deref_2619_resized_base_address, req => ptr_deref_2619_base_resize_req_0, ack => ptr_deref_2619_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2643_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp181_2640, dout => ptr_deref_2643_resized_base_address, req => ptr_deref_2643_base_resize_req_0, ack => ptr_deref_2643_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2661_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp185_2658, dout => ptr_deref_2661_resized_base_address, req => ptr_deref_2661_base_resize_req_0, ack => ptr_deref_2661_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2246_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp124_2243, dout => tmp125_2247, req => type_cast_2246_inst_req_0, ack => type_cast_2246_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2277_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp129_2274, dout => tmp3_2278, req => type_cast_2277_inst_req_0, ack => type_cast_2277_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2290_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp131_2287, dout => tmp5_2291, req => type_cast_2290_inst_req_0, ack => type_cast_2290_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2309_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp133_2306, dout => tmp10_2310, req => type_cast_2309_inst_req_0, ack => type_cast_2309_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2328_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp135_2325, dout => tmp15_2329, req => type_cast_2328_inst_req_0, ack => type_cast_2328_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2347_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp137_2344, dout => tmp20_2348, req => type_cast_2347_inst_req_0, ack => type_cast_2347_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2366_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp139_2363, dout => tmp25_2367, req => type_cast_2366_inst_req_0, ack => type_cast_2366_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2380_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp140_2377, dout => tmp30_2381, req => type_cast_2380_inst_req_0, ack => type_cast_2380_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2399_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp142_2396, dout => tmp35_2400, req => type_cast_2399_inst_req_0, ack => type_cast_2399_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2473_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => phitmp_2739, dout => type_cast_2473_wire, req => type_cast_2473_inst_req_0, ack => type_cast_2473_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2480_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => indvar_2469, dout => tmp144_2481, req => type_cast_2480_inst_req_0, ack => type_cast_2480_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2509_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp152_2506, dout => tmp40_2510, req => type_cast_2509_inst_req_0, ack => type_cast_2509_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2527_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp157_2524, dout => tmp44_2528, req => type_cast_2527_inst_req_0, ack => type_cast_2527_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2551_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp162_2548, dout => tmp49_2552, req => type_cast_2551_inst_req_0, ack => type_cast_2551_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2575_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp167_2572, dout => tmp54_2576, req => type_cast_2575_inst_req_0, ack => type_cast_2575_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2599_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp172_2596, dout => tmp59_2600, req => type_cast_2599_inst_req_0, ack => type_cast_2599_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2623_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp177_2620, dout => tmp64_2624, req => type_cast_2623_inst_req_0, ack => type_cast_2623_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2647_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp182_2644, dout => tmp69_2648, req => type_cast_2647_inst_req_0, ack => type_cast_2647_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2665_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp186_2662, dout => tmp74_2666, req => type_cast_2665_inst_req_0, ack => type_cast_2665_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2501_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2501_index_0_rename_ack_0 <= array_obj_ref_2501_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2500_resized;
      simple_obj_ref_2500_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2519_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2519_index_0_rename_ack_0 <= array_obj_ref_2519_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2518_resized;
      simple_obj_ref_2518_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2543_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2543_index_0_rename_ack_0 <= array_obj_ref_2543_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2542_resized;
      simple_obj_ref_2542_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2567_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2567_index_0_rename_ack_0 <= array_obj_ref_2567_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2566_resized;
      simple_obj_ref_2566_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2591_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2591_index_0_rename_ack_0 <= array_obj_ref_2591_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2590_resized;
      simple_obj_ref_2590_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2615_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2615_index_0_rename_ack_0 <= array_obj_ref_2615_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2614_resized;
      simple_obj_ref_2614_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2639_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2639_index_0_rename_ack_0 <= array_obj_ref_2639_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2638_resized;
      simple_obj_ref_2638_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2657_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2657_index_0_rename_ack_0 <= array_obj_ref_2657_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2656_resized;
      simple_obj_ref_2656_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2273_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2273_addr_0_ack_0 <= ptr_deref_2273_addr_0_req_0;
      aggregated_sig <= ptr_deref_2273_root_address;
      ptr_deref_2273_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2273_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2273_gather_scatter_ack_0 <= ptr_deref_2273_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2273_data_0;
      tmp129_2274 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2273_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2273_root_address_inst_ack_0 <= ptr_deref_2273_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2273_resized_base_address;
      ptr_deref_2273_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2286_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2286_addr_0_ack_0 <= ptr_deref_2286_addr_0_req_0;
      aggregated_sig <= ptr_deref_2286_root_address;
      ptr_deref_2286_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2286_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2286_gather_scatter_ack_0 <= ptr_deref_2286_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2286_data_0;
      tmp131_2287 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2286_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2286_root_address_inst_ack_0 <= ptr_deref_2286_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2286_resized_base_address;
      ptr_deref_2286_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2305_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2305_addr_0_ack_0 <= ptr_deref_2305_addr_0_req_0;
      aggregated_sig <= ptr_deref_2305_root_address;
      ptr_deref_2305_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2305_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2305_gather_scatter_ack_0 <= ptr_deref_2305_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2305_data_0;
      tmp133_2306 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2305_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2305_root_address_inst_ack_0 <= ptr_deref_2305_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2305_resized_base_address;
      ptr_deref_2305_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2324_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2324_addr_0_ack_0 <= ptr_deref_2324_addr_0_req_0;
      aggregated_sig <= ptr_deref_2324_root_address;
      ptr_deref_2324_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2324_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2324_gather_scatter_ack_0 <= ptr_deref_2324_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2324_data_0;
      tmp135_2325 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2324_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2324_root_address_inst_ack_0 <= ptr_deref_2324_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2324_resized_base_address;
      ptr_deref_2324_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2343_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2343_addr_0_ack_0 <= ptr_deref_2343_addr_0_req_0;
      aggregated_sig <= ptr_deref_2343_root_address;
      ptr_deref_2343_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2343_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2343_gather_scatter_ack_0 <= ptr_deref_2343_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2343_data_0;
      tmp137_2344 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2343_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2343_root_address_inst_ack_0 <= ptr_deref_2343_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2343_resized_base_address;
      ptr_deref_2343_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2362_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2362_addr_0_ack_0 <= ptr_deref_2362_addr_0_req_0;
      aggregated_sig <= ptr_deref_2362_root_address;
      ptr_deref_2362_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2362_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2362_gather_scatter_ack_0 <= ptr_deref_2362_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2362_data_0;
      tmp139_2363 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2362_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2362_root_address_inst_ack_0 <= ptr_deref_2362_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2362_resized_base_address;
      ptr_deref_2362_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2376_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2376_addr_0_ack_0 <= ptr_deref_2376_addr_0_req_0;
      aggregated_sig <= ptr_deref_2376_root_address;
      ptr_deref_2376_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2376_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2376_gather_scatter_ack_0 <= ptr_deref_2376_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2376_data_0;
      tmp140_2377 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2376_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2376_root_address_inst_ack_0 <= ptr_deref_2376_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2376_resized_base_address;
      ptr_deref_2376_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2395_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2395_addr_0_ack_0 <= ptr_deref_2395_addr_0_req_0;
      aggregated_sig <= ptr_deref_2395_root_address;
      ptr_deref_2395_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2395_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2395_gather_scatter_ack_0 <= ptr_deref_2395_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2395_data_0;
      tmp142_2396 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2395_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2395_root_address_inst_ack_0 <= ptr_deref_2395_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2395_resized_base_address;
      ptr_deref_2395_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2505_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2505_addr_0_ack_0 <= ptr_deref_2505_addr_0_req_0;
      aggregated_sig <= ptr_deref_2505_root_address;
      ptr_deref_2505_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2505_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2505_gather_scatter_ack_0 <= ptr_deref_2505_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2505_data_0;
      tmp152_2506 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2505_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2505_root_address_inst_ack_0 <= ptr_deref_2505_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2505_resized_base_address;
      ptr_deref_2505_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2523_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2523_addr_0_ack_0 <= ptr_deref_2523_addr_0_req_0;
      aggregated_sig <= ptr_deref_2523_root_address;
      ptr_deref_2523_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2523_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2523_gather_scatter_ack_0 <= ptr_deref_2523_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2523_data_0;
      tmp157_2524 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2523_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2523_root_address_inst_ack_0 <= ptr_deref_2523_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2523_resized_base_address;
      ptr_deref_2523_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2547_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2547_addr_0_ack_0 <= ptr_deref_2547_addr_0_req_0;
      aggregated_sig <= ptr_deref_2547_root_address;
      ptr_deref_2547_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2547_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2547_gather_scatter_ack_0 <= ptr_deref_2547_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2547_data_0;
      tmp162_2548 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2547_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2547_root_address_inst_ack_0 <= ptr_deref_2547_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2547_resized_base_address;
      ptr_deref_2547_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2571_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2571_addr_0_ack_0 <= ptr_deref_2571_addr_0_req_0;
      aggregated_sig <= ptr_deref_2571_root_address;
      ptr_deref_2571_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2571_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2571_gather_scatter_ack_0 <= ptr_deref_2571_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2571_data_0;
      tmp167_2572 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2571_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2571_root_address_inst_ack_0 <= ptr_deref_2571_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2571_resized_base_address;
      ptr_deref_2571_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2595_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2595_addr_0_ack_0 <= ptr_deref_2595_addr_0_req_0;
      aggregated_sig <= ptr_deref_2595_root_address;
      ptr_deref_2595_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2595_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2595_gather_scatter_ack_0 <= ptr_deref_2595_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2595_data_0;
      tmp172_2596 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2595_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2595_root_address_inst_ack_0 <= ptr_deref_2595_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2595_resized_base_address;
      ptr_deref_2595_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2619_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2619_addr_0_ack_0 <= ptr_deref_2619_addr_0_req_0;
      aggregated_sig <= ptr_deref_2619_root_address;
      ptr_deref_2619_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2619_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2619_gather_scatter_ack_0 <= ptr_deref_2619_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2619_data_0;
      tmp177_2620 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2619_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2619_root_address_inst_ack_0 <= ptr_deref_2619_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2619_resized_base_address;
      ptr_deref_2619_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2643_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2643_addr_0_ack_0 <= ptr_deref_2643_addr_0_req_0;
      aggregated_sig <= ptr_deref_2643_root_address;
      ptr_deref_2643_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2643_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2643_gather_scatter_ack_0 <= ptr_deref_2643_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2643_data_0;
      tmp182_2644 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2643_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2643_root_address_inst_ack_0 <= ptr_deref_2643_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2643_resized_base_address;
      ptr_deref_2643_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2661_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2661_addr_0_ack_0 <= ptr_deref_2661_addr_0_req_0;
      aggregated_sig <= ptr_deref_2661_root_address;
      ptr_deref_2661_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2661_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2661_gather_scatter_ack_0 <= ptr_deref_2661_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2661_data_0;
      tmp186_2662 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2661_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2661_root_address_inst_ack_0 <= ptr_deref_2661_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2661_resized_base_address;
      ptr_deref_2661_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_2714_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp146_2486;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2714_branch_req_0,
          ack0 => if_stmt_2714_branch_ack_0,
          ack1 => if_stmt_2714_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_2269_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2269_resized_base_address;
      array_obj_ref_2269_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000111",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2269_root_address_inst_req_0,
          ackL => array_obj_ref_2269_root_address_inst_ack_0,
          reqR => array_obj_ref_2269_root_address_inst_req_1,
          ackR => array_obj_ref_2269_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2282_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2282_resized_base_address;
      array_obj_ref_2282_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000110",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2282_root_address_inst_req_0,
          ackL => array_obj_ref_2282_root_address_inst_ack_0,
          reqR => array_obj_ref_2282_root_address_inst_req_1,
          ackR => array_obj_ref_2282_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_2301_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2301_resized_base_address;
      array_obj_ref_2301_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000101",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2301_root_address_inst_req_0,
          ackL => array_obj_ref_2301_root_address_inst_ack_0,
          reqR => array_obj_ref_2301_root_address_inst_req_1,
          ackR => array_obj_ref_2301_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_2320_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2320_resized_base_address;
      array_obj_ref_2320_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2320_root_address_inst_req_0,
          ackL => array_obj_ref_2320_root_address_inst_ack_0,
          reqR => array_obj_ref_2320_root_address_inst_req_1,
          ackR => array_obj_ref_2320_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_2339_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2339_resized_base_address;
      array_obj_ref_2339_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2339_root_address_inst_req_0,
          ackL => array_obj_ref_2339_root_address_inst_ack_0,
          reqR => array_obj_ref_2339_root_address_inst_req_1,
          ackR => array_obj_ref_2339_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_2358_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2358_resized_base_address;
      array_obj_ref_2358_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2358_root_address_inst_req_0,
          ackL => array_obj_ref_2358_root_address_inst_ack_0,
          reqR => array_obj_ref_2358_root_address_inst_req_1,
          ackR => array_obj_ref_2358_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_2391_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2391_resized_base_address;
      array_obj_ref_2391_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2391_root_address_inst_req_0,
          ackL => array_obj_ref_2391_root_address_inst_ack_0,
          reqR => array_obj_ref_2391_root_address_inst_req_1,
          ackR => array_obj_ref_2391_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_2501_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2501_final_offset & array_obj_ref_2501_resized_base_address;
      array_obj_ref_2501_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2501_root_address_inst_req_0,
          ackL => array_obj_ref_2501_root_address_inst_ack_0,
          reqR => array_obj_ref_2501_root_address_inst_req_1,
          ackR => array_obj_ref_2501_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_2519_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2519_final_offset & array_obj_ref_2519_resized_base_address;
      array_obj_ref_2519_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2519_root_address_inst_req_0,
          ackL => array_obj_ref_2519_root_address_inst_ack_0,
          reqR => array_obj_ref_2519_root_address_inst_req_1,
          ackR => array_obj_ref_2519_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_2543_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2543_final_offset & array_obj_ref_2543_resized_base_address;
      array_obj_ref_2543_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2543_root_address_inst_req_0,
          ackL => array_obj_ref_2543_root_address_inst_ack_0,
          reqR => array_obj_ref_2543_root_address_inst_req_1,
          ackR => array_obj_ref_2543_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_2567_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2567_final_offset & array_obj_ref_2567_resized_base_address;
      array_obj_ref_2567_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2567_root_address_inst_req_0,
          ackL => array_obj_ref_2567_root_address_inst_ack_0,
          reqR => array_obj_ref_2567_root_address_inst_req_1,
          ackR => array_obj_ref_2567_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_2591_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2591_final_offset & array_obj_ref_2591_resized_base_address;
      array_obj_ref_2591_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2591_root_address_inst_req_0,
          ackL => array_obj_ref_2591_root_address_inst_ack_0,
          reqR => array_obj_ref_2591_root_address_inst_req_1,
          ackR => array_obj_ref_2591_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_2615_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2615_final_offset & array_obj_ref_2615_resized_base_address;
      array_obj_ref_2615_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2615_root_address_inst_req_0,
          ackL => array_obj_ref_2615_root_address_inst_ack_0,
          reqR => array_obj_ref_2615_root_address_inst_req_1,
          ackR => array_obj_ref_2615_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_2639_root_address_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2639_final_offset & array_obj_ref_2639_resized_base_address;
      array_obj_ref_2639_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2639_root_address_inst_req_0,
          ackL => array_obj_ref_2639_root_address_inst_ack_0,
          reqR => array_obj_ref_2639_root_address_inst_req_1,
          ackR => array_obj_ref_2639_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_2657_root_address_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2657_final_offset & array_obj_ref_2657_resized_base_address;
      array_obj_ref_2657_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2657_root_address_inst_req_0,
          ackL => array_obj_ref_2657_root_address_inst_ack_0,
          reqR => array_obj_ref_2657_root_address_inst_req_1,
          ackR => array_obj_ref_2657_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_2296_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp5_2291;
      tmp6_2297 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2296_inst_req_0,
          ackL => binary_2296_inst_ack_0,
          reqR => binary_2296_inst_req_1,
          ackR => binary_2296_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_2315_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp10_2310;
      tmp11_2316 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2315_inst_req_0,
          ackL => binary_2315_inst_ack_0,
          reqR => binary_2315_inst_req_1,
          ackR => binary_2315_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_2334_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2329;
      tmp16_2335 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2334_inst_req_0,
          ackL => binary_2334_inst_ack_0,
          reqR => binary_2334_inst_req_1,
          ackR => binary_2334_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_2353_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_2348;
      tmp21_2354 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2353_inst_req_0,
          ackL => binary_2353_inst_ack_0,
          reqR => binary_2353_inst_req_1,
          ackR => binary_2353_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_2372_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp25_2367;
      tmp26_2373 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2372_inst_req_0,
          ackL => binary_2372_inst_ack_0,
          reqR => binary_2372_inst_req_1,
          ackR => binary_2372_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_2386_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_2381;
      tmp31_2387 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2386_inst_req_0,
          ackL => binary_2386_inst_ack_0,
          reqR => binary_2386_inst_req_1,
          ackR => binary_2386_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_2405_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp35_2400;
      tmp36_2406 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2405_inst_req_0,
          ackL => binary_2405_inst_ack_0,
          reqR => binary_2405_inst_req_1,
          ackR => binary_2405_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_2410_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_2297 & tmp3_2278;
      mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_2411 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2410_inst_req_0,
          ackL => binary_2410_inst_ack_0,
          reqR => binary_2410_inst_req_1,
          ackR => binary_2410_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_2415_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_2411 & tmp11_2316;
      mask17x_xmaskedx_xmaskedx_xmasked_2416 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2415_inst_req_0,
          ackL => binary_2415_inst_ack_0,
          reqR => binary_2415_inst_req_1,
          ackR => binary_2415_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_2420_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask17x_xmaskedx_xmaskedx_xmasked_2416 & tmp16_2335;
      mask22x_xmaskedx_xmaskedx_xmasked_2421 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2420_inst_req_0,
          ackL => binary_2420_inst_ack_0,
          reqR => binary_2420_inst_req_1,
          ackR => binary_2420_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_2425_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask22x_xmaskedx_xmaskedx_xmasked_2421 & tmp21_2354;
      mask27x_xmaskedx_xmasked_2426 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2425_inst_req_0,
          ackL => binary_2425_inst_ack_0,
          reqR => binary_2425_inst_req_1,
          ackR => binary_2425_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_2430_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask27x_xmaskedx_xmasked_2426 & tmp26_2373;
      mask32x_xmasked_2431 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2430_inst_req_0,
          ackL => binary_2430_inst_ack_0,
          reqR => binary_2430_inst_req_1,
          ackR => binary_2430_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_2435_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask32x_xmasked_2431 & tmp31_2387;
      mask37_2436 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2435_inst_req_0,
          ackL => binary_2435_inst_ack_0,
          reqR => binary_2435_inst_req_1,
          ackR => binary_2435_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_2440_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask37_2436 & tmp36_2406;
      ins38_2441 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2440_inst_req_0,
          ackL => binary_2440_inst_ack_0,
          reqR => binary_2440_inst_req_1,
          ackR => binary_2440_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_2465_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp126_2256;
      tmp145_2466 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2465_inst_req_0,
          ackL => binary_2465_inst_ack_0,
          reqR => binary_2465_inst_req_1,
          ackR => binary_2465_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_2485_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp144_2481 & tmp145_2466;
      tmp146_2486 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2485_inst_req_0,
          ackL => binary_2485_inst_ack_0,
          reqR => binary_2485_inst_req_1,
          ackR => binary_2485_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_2491_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp144_2481;
      tmp149_2492 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2491_inst_req_0,
          ackL => binary_2491_inst_ack_0,
          reqR => binary_2491_inst_req_1,
          ackR => binary_2491_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_2497_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp150_2498 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2497_inst_req_0,
          ackL => binary_2497_inst_ack_0,
          reqR => binary_2497_inst_req_1,
          ackR => binary_2497_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_2515_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp155_2516 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2515_inst_req_0,
          ackL => binary_2515_inst_ack_0,
          reqR => binary_2515_inst_req_1,
          ackR => binary_2515_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_2533_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp44_2528;
      tmp45_2534 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2533_inst_req_0,
          ackL => binary_2533_inst_ack_0,
          reqR => binary_2533_inst_req_1,
          ackR => binary_2533_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_2539_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp160_2540 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2539_inst_req_0,
          ackL => binary_2539_inst_ack_0,
          reqR => binary_2539_inst_req_1,
          ackR => binary_2539_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_2557_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp49_2552;
      tmp50_2558 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2557_inst_req_0,
          ackL => binary_2557_inst_ack_0,
          reqR => binary_2557_inst_req_1,
          ackR => binary_2557_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_2563_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp165_2564 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2563_inst_req_0,
          ackL => binary_2563_inst_ack_0,
          reqR => binary_2563_inst_req_1,
          ackR => binary_2563_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_2581_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp54_2576;
      tmp55_2582 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2581_inst_req_0,
          ackL => binary_2581_inst_ack_0,
          reqR => binary_2581_inst_req_1,
          ackR => binary_2581_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_2587_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp170_2588 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2587_inst_req_0,
          ackL => binary_2587_inst_ack_0,
          reqR => binary_2587_inst_req_1,
          ackR => binary_2587_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_2605_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp59_2600;
      tmp60_2606 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2605_inst_req_0,
          ackL => binary_2605_inst_ack_0,
          reqR => binary_2605_inst_req_1,
          ackR => binary_2605_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_2611_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp175_2612 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2611_inst_req_0,
          ackL => binary_2611_inst_ack_0,
          reqR => binary_2611_inst_req_1,
          ackR => binary_2611_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_2629_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp64_2624;
      tmp65_2630 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2629_inst_req_0,
          ackL => binary_2629_inst_ack_0,
          reqR => binary_2629_inst_req_1,
          ackR => binary_2629_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_2635_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp149_2492;
      tmp180_2636 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2635_inst_req_0,
          ackL => binary_2635_inst_ack_0,
          reqR => binary_2635_inst_req_1,
          ackR => binary_2635_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_2653_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp69_2648;
      tmp70_2654 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2653_inst_req_0,
          ackL => binary_2653_inst_ack_0,
          reqR => binary_2653_inst_req_1,
          ackR => binary_2653_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_2671_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_2666;
      tmp75_2672 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2671_inst_req_0,
          ackL => binary_2671_inst_ack_0,
          reqR => binary_2671_inst_req_1,
          ackR => binary_2671_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_2676_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp45_2534 & tmp40_2510;
      mask51_2677 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2676_inst_req_0,
          ackL => binary_2676_inst_ack_0,
          reqR => binary_2676_inst_req_1,
          ackR => binary_2676_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_2681_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask51_2677 & tmp50_2558;
      mask56_2682 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2681_inst_req_0,
          ackL => binary_2681_inst_ack_0,
          reqR => binary_2681_inst_req_1,
          ackR => binary_2681_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_2686_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask56_2682 & tmp55_2582;
      mask61x_xmaskedx_xmasked_2687 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2686_inst_req_0,
          ackL => binary_2686_inst_ack_0,
          reqR => binary_2686_inst_req_1,
          ackR => binary_2686_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_2691_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask61x_xmaskedx_xmasked_2687 & tmp60_2606;
      mask66x_xmaskedx_xmasked_2692 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2691_inst_req_0,
          ackL => binary_2691_inst_ack_0,
          reqR => binary_2691_inst_req_1,
          ackR => binary_2691_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_2696_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask66x_xmaskedx_xmasked_2692 & tmp65_2630;
      mask71x_xmasked_2697 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2696_inst_req_0,
          ackL => binary_2696_inst_ack_0,
          reqR => binary_2696_inst_req_1,
          ackR => binary_2696_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_2701_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask71x_xmasked_2697 & tmp70_2654;
      mask76_2702 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2701_inst_req_0,
          ackL => binary_2701_inst_ack_0,
          reqR => binary_2701_inst_req_1,
          ackR => binary_2701_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_2706_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask76_2702 & tmp75_2672;
      ins77_2707 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2706_inst_req_0,
          ackL => binary_2706_inst_ack_0,
          reqR => binary_2706_inst_req_1,
          ackR => binary_2706_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_2738_inst 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_2469;
      phitmp_2739 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2738_inst_req_0,
          ackL => binary_2738_inst_ack_0,
          reqR => binary_2738_inst_req_1,
          ackR => binary_2738_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared load operator group (0) : ptr_deref_2273_load_0 ptr_deref_2505_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2273_load_0_req_0;
      reqL(0) <= ptr_deref_2505_load_0_req_0;
      ptr_deref_2273_load_0_ack_0 <= ackL(1);
      ptr_deref_2505_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2273_load_0_req_1;
      reqR(0) <= ptr_deref_2505_load_0_req_1;
      ptr_deref_2273_load_0_ack_1 <= ackR(1);
      ptr_deref_2505_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2273_word_address_0 & ptr_deref_2505_word_address_0;
      ptr_deref_2273_data_0 <= data_out(15 downto 8);
      ptr_deref_2505_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(7),
          mack => memory_space_3_lr_ack(7),
          maddr => memory_space_3_lr_addr(87 downto 77),
          mtag => memory_space_3_lr_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(7),
          mack => memory_space_3_lc_ack(7),
          mdata => memory_space_3_lc_data(63 downto 56),
          mtag => memory_space_3_lc_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2286_load_0 ptr_deref_2523_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2286_load_0_req_0;
      reqL(0) <= ptr_deref_2523_load_0_req_0;
      ptr_deref_2286_load_0_ack_0 <= ackL(1);
      ptr_deref_2523_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2286_load_0_req_1;
      reqR(0) <= ptr_deref_2523_load_0_req_1;
      ptr_deref_2286_load_0_ack_1 <= ackR(1);
      ptr_deref_2523_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2286_word_address_0 & ptr_deref_2523_word_address_0;
      ptr_deref_2286_data_0 <= data_out(15 downto 8);
      ptr_deref_2523_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(6),
          mack => memory_space_3_lr_ack(6),
          maddr => memory_space_3_lr_addr(76 downto 66),
          mtag => memory_space_3_lr_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(6),
          mack => memory_space_3_lc_ack(6),
          mdata => memory_space_3_lc_data(55 downto 48),
          mtag => memory_space_3_lc_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2305_load_0 ptr_deref_2547_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2305_load_0_req_0;
      reqL(0) <= ptr_deref_2547_load_0_req_0;
      ptr_deref_2305_load_0_ack_0 <= ackL(1);
      ptr_deref_2547_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2305_load_0_req_1;
      reqR(0) <= ptr_deref_2547_load_0_req_1;
      ptr_deref_2305_load_0_ack_1 <= ackR(1);
      ptr_deref_2547_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2305_word_address_0 & ptr_deref_2547_word_address_0;
      ptr_deref_2305_data_0 <= data_out(15 downto 8);
      ptr_deref_2547_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(5),
          mack => memory_space_3_lr_ack(5),
          maddr => memory_space_3_lr_addr(65 downto 55),
          mtag => memory_space_3_lr_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(5),
          mack => memory_space_3_lc_ack(5),
          mdata => memory_space_3_lc_data(47 downto 40),
          mtag => memory_space_3_lc_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2324_load_0 ptr_deref_2571_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2324_load_0_req_0;
      reqL(0) <= ptr_deref_2571_load_0_req_0;
      ptr_deref_2324_load_0_ack_0 <= ackL(1);
      ptr_deref_2571_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2324_load_0_req_1;
      reqR(0) <= ptr_deref_2571_load_0_req_1;
      ptr_deref_2324_load_0_ack_1 <= ackR(1);
      ptr_deref_2571_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2324_word_address_0 & ptr_deref_2571_word_address_0;
      ptr_deref_2324_data_0 <= data_out(15 downto 8);
      ptr_deref_2571_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(4),
          mack => memory_space_3_lr_ack(4),
          maddr => memory_space_3_lr_addr(54 downto 44),
          mtag => memory_space_3_lr_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(4),
          mack => memory_space_3_lc_ack(4),
          mdata => memory_space_3_lc_data(39 downto 32),
          mtag => memory_space_3_lc_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2343_load_0 ptr_deref_2595_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2343_load_0_req_0;
      reqL(0) <= ptr_deref_2595_load_0_req_0;
      ptr_deref_2343_load_0_ack_0 <= ackL(1);
      ptr_deref_2595_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2343_load_0_req_1;
      reqR(0) <= ptr_deref_2595_load_0_req_1;
      ptr_deref_2343_load_0_ack_1 <= ackR(1);
      ptr_deref_2595_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2343_word_address_0 & ptr_deref_2595_word_address_0;
      ptr_deref_2343_data_0 <= data_out(15 downto 8);
      ptr_deref_2595_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(3),
          mack => memory_space_3_lr_ack(3),
          maddr => memory_space_3_lr_addr(43 downto 33),
          mtag => memory_space_3_lr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(3),
          mack => memory_space_3_lc_ack(3),
          mdata => memory_space_3_lc_data(31 downto 24),
          mtag => memory_space_3_lc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2362_load_0 ptr_deref_2619_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2362_load_0_req_0;
      reqL(0) <= ptr_deref_2619_load_0_req_0;
      ptr_deref_2362_load_0_ack_0 <= ackL(1);
      ptr_deref_2619_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2362_load_0_req_1;
      reqR(0) <= ptr_deref_2619_load_0_req_1;
      ptr_deref_2362_load_0_ack_1 <= ackR(1);
      ptr_deref_2619_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2362_word_address_0 & ptr_deref_2619_word_address_0;
      ptr_deref_2362_data_0 <= data_out(15 downto 8);
      ptr_deref_2619_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(2),
          mack => memory_space_3_lr_ack(2),
          maddr => memory_space_3_lr_addr(32 downto 22),
          mtag => memory_space_3_lr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(2),
          mack => memory_space_3_lc_ack(2),
          mdata => memory_space_3_lc_data(23 downto 16),
          mtag => memory_space_3_lc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_2376_load_0 ptr_deref_2643_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2376_load_0_req_0;
      reqL(0) <= ptr_deref_2643_load_0_req_0;
      ptr_deref_2376_load_0_ack_0 <= ackL(1);
      ptr_deref_2643_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2376_load_0_req_1;
      reqR(0) <= ptr_deref_2643_load_0_req_1;
      ptr_deref_2376_load_0_ack_1 <= ackR(1);
      ptr_deref_2643_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2376_word_address_0 & ptr_deref_2643_word_address_0;
      ptr_deref_2376_data_0 <= data_out(15 downto 8);
      ptr_deref_2643_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(1),
          mack => memory_space_3_lr_ack(1),
          maddr => memory_space_3_lr_addr(21 downto 11),
          mtag => memory_space_3_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(1),
          mack => memory_space_3_lc_ack(1),
          mdata => memory_space_3_lc_data(15 downto 8),
          mtag => memory_space_3_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_2395_load_0 ptr_deref_2661_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2395_load_0_req_0;
      reqL(0) <= ptr_deref_2661_load_0_req_0;
      ptr_deref_2395_load_0_ack_0 <= ackL(1);
      ptr_deref_2661_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2395_load_0_req_1;
      reqR(0) <= ptr_deref_2661_load_0_req_1;
      ptr_deref_2395_load_0_ack_1 <= ackR(1);
      ptr_deref_2661_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2395_word_address_0 & ptr_deref_2661_word_address_0;
      ptr_deref_2395_data_0 <= data_out(15 downto 8);
      ptr_deref_2661_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(10 downto 0),
          mtag => memory_space_3_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared inport operator group (0) : simple_obj_ref_2231_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2231_inst_req_0;
      simple_obj_ref_2231_inst_ack_0 <= ack(0);
      tmp_2232 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => start_wrapper_output_pipe_read_req(0),
          oack => start_wrapper_output_pipe_read_ack(0),
          odata => start_wrapper_output_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_2242_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2242_inst_req_0;
      simple_obj_ref_2242_inst_ack_0 <= ack(0);
      tmp124_2243 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => midpipe_pipe_read_req(0),
          oack => midpipe_pipe_read_ack(0),
          odata => midpipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_2255_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2255_inst_req_0;
      simple_obj_ref_2255_inst_ack_0 <= ack(0);
      tmp126_2256 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => pkt_length_pipe_read_req(0),
          oack => pkt_length_pipe_read_ack(0),
          odata => pkt_length_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_2264_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2264_inst_req_0;
      simple_obj_ref_2264_inst_ack_0 <= ack(0);
      tmp127_2265 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => last_ctrl_pipe_read_req(0),
          oack => last_ctrl_pipe_read_ack(0),
          odata => last_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : simple_obj_ref_2448_inst simple_obj_ref_2721_inst simple_obj_ref_2742_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_2448_inst_req_0;
      req(1) <= simple_obj_ref_2721_inst_req_0;
      req(0) <= simple_obj_ref_2742_inst_req_0;
      simple_obj_ref_2448_inst_ack_0 <= ack(2);
      simple_obj_ref_2721_inst_ack_0 <= ack(1);
      simple_obj_ref_2742_inst_ack_0 <= ack(0);
      data_in <= type_cast_2450_wire_constant & type_cast_2723_wire_constant & tmp127_2265;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 3,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => op_lut_ctrl_pipe_write_req(0),
          oack => op_lut_ctrl_pipe_write_ack(0),
          odata => op_lut_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_2458_inst simple_obj_ref_2731_inst simple_obj_ref_2751_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_2458_inst_req_0;
      req(1) <= simple_obj_ref_2731_inst_req_0;
      req(0) <= simple_obj_ref_2751_inst_req_0;
      simple_obj_ref_2458_inst_ack_0 <= ack(2);
      simple_obj_ref_2731_inst_ack_0 <= ack(1);
      simple_obj_ref_2751_inst_ack_0 <= ack(0);
      data_in <= ins38_2441 & ins77_2707 & ins77_2707;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 3,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => op_lut_data_pipe_write_req(0),
          oack => op_lut_data_pipe_write_ack(0),
          odata => op_lut_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_2760_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2760_inst_req_0;
      simple_obj_ref_2760_inst_ack_0 <= ack(0);
      data_in <= type_cast_2762_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : simple_obj_ref_2770_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2770_inst_req_0;
      simple_obj_ref_2770_inst_ack_0 <= ack(0);
      data_in <= tmp124_2243;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_put_pipe_write_req(0),
          oack => free_queue_put_pipe_write_ack(0),
          odata => free_queue_put_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
    in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
    in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
    out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_10
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_11
  signal memory_space_11_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_11_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_11_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_11_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_12
  signal memory_space_12_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_12_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_12_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_12_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_13
  signal memory_space_13_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_13_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_13_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_13_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_14
  signal memory_space_14_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_14_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_14_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_14_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_14_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_14_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_14_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_15
  signal memory_space_15_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_15_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_15_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_15_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_15_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_15_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_15_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_16
  signal memory_space_16_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_16_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_16_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_16_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_17
  signal memory_space_17_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_17_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_17_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_17_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_18
  signal memory_space_18_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_18_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_18_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_18_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_18_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_18_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_18_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_18_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_19
  signal memory_space_19_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_19_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_19_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_19_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_19_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_19_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_19_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_19_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(14 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(39 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(9 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(9 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(7 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(7 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(87 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(15 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(15 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(8 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(8 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(98 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(71 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(8 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(8 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(17 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_9
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module default_initializer_foo
  component default_initializer_foo is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_foo
  signal default_initializer_foo_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_foo_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_foo_start_req : std_logic;
  signal default_initializer_foo_start_ack : std_logic;
  signal default_initializer_foo_fin_req   : std_logic;
  signal default_initializer_foo_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_foo
  signal default_initializer_foo_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_foo_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_foo_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_foo_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_foo_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_foo_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_free_queue
  component default_initializer_free_queue is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_free_queue
  signal default_initializer_free_queue_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_free_queue_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_start_req : std_logic;
  signal default_initializer_free_queue_start_ack : std_logic;
  signal default_initializer_free_queue_fin_req   : std_logic;
  signal default_initializer_free_queue_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_free_queue
  signal default_initializer_free_queue_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_free_queue_ram
  component default_initializer_free_queue_ram is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_free_queue_ram
  signal default_initializer_free_queue_ram_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_free_queue_ram_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_start_req : std_logic;
  signal default_initializer_free_queue_ram_start_ack : std_logic;
  signal default_initializer_free_queue_ram_fin_req   : std_logic;
  signal default_initializer_free_queue_ram_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_free_queue_ram
  signal default_initializer_free_queue_ram_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr
  component default_initializer_xx_xstr is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr
  signal default_initializer_xx_xstr_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_start_req : std_logic;
  signal default_initializer_xx_xstr_start_ack : std_logic;
  signal default_initializer_xx_xstr_fin_req   : std_logic;
  signal default_initializer_xx_xstr_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr
  signal default_initializer_xx_xstr_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr1
  component default_initializer_xx_xstr1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr1
  signal default_initializer_xx_xstr1_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr1_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_start_req : std_logic;
  signal default_initializer_xx_xstr1_start_ack : std_logic;
  signal default_initializer_xx_xstr1_fin_req   : std_logic;
  signal default_initializer_xx_xstr1_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr1
  signal default_initializer_xx_xstr1_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr10
  component default_initializer_xx_xstr10 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr10
  signal default_initializer_xx_xstr10_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr10_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr10_start_req : std_logic;
  signal default_initializer_xx_xstr10_start_ack : std_logic;
  signal default_initializer_xx_xstr10_fin_req   : std_logic;
  signal default_initializer_xx_xstr10_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr10
  signal default_initializer_xx_xstr10_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr10_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr10_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr10_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr10_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr10_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr11
  component default_initializer_xx_xstr11 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr11
  signal default_initializer_xx_xstr11_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr11_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr11_start_req : std_logic;
  signal default_initializer_xx_xstr11_start_ack : std_logic;
  signal default_initializer_xx_xstr11_fin_req   : std_logic;
  signal default_initializer_xx_xstr11_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr11
  signal default_initializer_xx_xstr11_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr11_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr11_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr11_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr11_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr11_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr12
  component default_initializer_xx_xstr12 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr12
  signal default_initializer_xx_xstr12_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr12_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr12_start_req : std_logic;
  signal default_initializer_xx_xstr12_start_ack : std_logic;
  signal default_initializer_xx_xstr12_fin_req   : std_logic;
  signal default_initializer_xx_xstr12_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr12
  signal default_initializer_xx_xstr12_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr12_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr12_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr12_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr12_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr12_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr13
  component default_initializer_xx_xstr13 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_9_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr13
  signal default_initializer_xx_xstr13_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr13_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr13_start_req : std_logic;
  signal default_initializer_xx_xstr13_start_ack : std_logic;
  signal default_initializer_xx_xstr13_fin_req   : std_logic;
  signal default_initializer_xx_xstr13_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr13
  signal default_initializer_xx_xstr13_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr13_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr13_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr13_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr13_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr13_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr14
  component default_initializer_xx_xstr14 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_10_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr14
  signal default_initializer_xx_xstr14_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr14_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr14_start_req : std_logic;
  signal default_initializer_xx_xstr14_start_ack : std_logic;
  signal default_initializer_xx_xstr14_fin_req   : std_logic;
  signal default_initializer_xx_xstr14_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr14
  signal default_initializer_xx_xstr14_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr14_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr14_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr14_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr14_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr14_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr15
  component default_initializer_xx_xstr15 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_11_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_11_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr15
  signal default_initializer_xx_xstr15_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr15_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr15_start_req : std_logic;
  signal default_initializer_xx_xstr15_start_ack : std_logic;
  signal default_initializer_xx_xstr15_fin_req   : std_logic;
  signal default_initializer_xx_xstr15_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr15
  signal default_initializer_xx_xstr15_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr15_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr15_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr15_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr15_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr15_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr2
  component default_initializer_xx_xstr2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_12_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_12_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_12_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_12_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_12_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_12_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr2
  signal default_initializer_xx_xstr2_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr2_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_start_req : std_logic;
  signal default_initializer_xx_xstr2_start_ack : std_logic;
  signal default_initializer_xx_xstr2_fin_req   : std_logic;
  signal default_initializer_xx_xstr2_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr2
  signal default_initializer_xx_xstr2_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr3
  component default_initializer_xx_xstr3 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_13_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_13_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_13_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_13_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_13_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_13_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr3
  signal default_initializer_xx_xstr3_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr3_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_start_req : std_logic;
  signal default_initializer_xx_xstr3_start_ack : std_logic;
  signal default_initializer_xx_xstr3_fin_req   : std_logic;
  signal default_initializer_xx_xstr3_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr3
  signal default_initializer_xx_xstr3_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr4
  component default_initializer_xx_xstr4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_14_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_14_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_14_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_14_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_14_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_14_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_14_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_14_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr4
  signal default_initializer_xx_xstr4_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr4_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_start_req : std_logic;
  signal default_initializer_xx_xstr4_start_ack : std_logic;
  signal default_initializer_xx_xstr4_fin_req   : std_logic;
  signal default_initializer_xx_xstr4_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr4
  signal default_initializer_xx_xstr4_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr5
  component default_initializer_xx_xstr5 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_15_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_15_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_15_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_15_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_15_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_15_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_15_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_15_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr5
  signal default_initializer_xx_xstr5_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr5_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_start_req : std_logic;
  signal default_initializer_xx_xstr5_start_ack : std_logic;
  signal default_initializer_xx_xstr5_fin_req   : std_logic;
  signal default_initializer_xx_xstr5_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr5
  signal default_initializer_xx_xstr5_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr6
  component default_initializer_xx_xstr6 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_16_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_16_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_16_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_16_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_16_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_16_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_16_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_16_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr6
  signal default_initializer_xx_xstr6_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr6_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_start_req : std_logic;
  signal default_initializer_xx_xstr6_start_ack : std_logic;
  signal default_initializer_xx_xstr6_fin_req   : std_logic;
  signal default_initializer_xx_xstr6_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr6
  signal default_initializer_xx_xstr6_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr7
  component default_initializer_xx_xstr7 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_17_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_17_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_17_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_17_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_17_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_17_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_17_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_17_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr7
  signal default_initializer_xx_xstr7_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr7_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_start_req : std_logic;
  signal default_initializer_xx_xstr7_start_ack : std_logic;
  signal default_initializer_xx_xstr7_fin_req   : std_logic;
  signal default_initializer_xx_xstr7_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr7
  signal default_initializer_xx_xstr7_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr8
  component default_initializer_xx_xstr8 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_18_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_18_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_18_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_18_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_18_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_18_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_18_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_18_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr8
  signal default_initializer_xx_xstr8_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr8_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_start_req : std_logic;
  signal default_initializer_xx_xstr8_start_ack : std_logic;
  signal default_initializer_xx_xstr8_fin_req   : std_logic;
  signal default_initializer_xx_xstr8_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr8
  signal default_initializer_xx_xstr8_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr9
  component default_initializer_xx_xstr9 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_19_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_19_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_19_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_19_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_19_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_19_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_19_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_19_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr9
  signal default_initializer_xx_xstr9_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr9_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr9_start_req : std_logic;
  signal default_initializer_xx_xstr9_start_ack : std_logic;
  signal default_initializer_xx_xstr9_fin_req   : std_logic;
  signal default_initializer_xx_xstr9_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr9
  signal default_initializer_xx_xstr9_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr9_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr9_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr9_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr9_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr9_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module free_queue_manager
  component free_queue_manager is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(3 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(3 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(3 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(7 downto 0);
      free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_ack_pipe_write_data : out  std_logic_vector(7 downto 0);
      free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
      start_output_port_lookup_pipe_write_req : out  std_logic_vector(0 downto 0);
      start_output_port_lookup_pipe_write_ack : in   std_logic_vector(0 downto 0);
      start_output_port_lookup_pipe_write_data : out  std_logic_vector(7 downto 0);
      start_wrapper_input_pipe_write_req : out  std_logic_vector(0 downto 0);
      start_wrapper_input_pipe_write_ack : in   std_logic_vector(0 downto 0);
      start_wrapper_input_pipe_write_data : out  std_logic_vector(7 downto 0);
      start_wrapper_output_pipe_write_req : out  std_logic_vector(0 downto 0);
      start_wrapper_output_pipe_write_ack : in   std_logic_vector(0 downto 0);
      start_wrapper_output_pipe_write_data : out  std_logic_vector(7 downto 0);
      global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_manager
  signal free_queue_manager_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal free_queue_manager_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_manager_start_req : std_logic;
  signal free_queue_manager_start_ack : std_logic;
  signal free_queue_manager_fin_req   : std_logic;
  signal free_queue_manager_fin_ack : std_logic;
  -- declarations related to module global_storage_initializer_x
  component global_storage_initializer_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      default_initializer_foo_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_foo_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_foo_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_foo_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_foo_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_foo_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr12_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr12_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr12_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr12_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr12_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr12_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr13_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr13_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr13_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr13_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr13_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr13_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr10_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr10_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr10_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr10_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr10_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr10_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr11_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr11_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr11_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr11_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr11_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr11_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr14_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr14_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr14_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr14_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr14_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr14_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr15_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr15_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr15_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr15_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr15_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr15_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr9_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr9_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr9_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr9_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr9_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr9_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module global_storage_initializer_x
  signal global_storage_initializer_x_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal global_storage_initializer_x_tag_out   : std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_start_req : std_logic;
  signal global_storage_initializer_x_start_ack : std_logic;
  signal global_storage_initializer_x_fin_req   : std_logic;
  signal global_storage_initializer_x_fin_ack : std_logic;
  -- caller side aggregated signals for module global_storage_initializer_x
  signal global_storage_initializer_x_call_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_tag: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module output_port_lookup
  component output_port_lookup is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      op_lut_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      op_lut_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      op_lut_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      op_lut_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      start_output_port_lookup_pipe_read_req : out  std_logic_vector(0 downto 0);
      start_output_port_lookup_pipe_read_ack : in   std_logic_vector(0 downto 0);
      start_output_port_lookup_pipe_read_data : in   std_logic_vector(7 downto 0);
      out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module output_port_lookup
  signal output_port_lookup_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal output_port_lookup_tag_out   : std_logic_vector(0 downto 0);
  signal output_port_lookup_start_req : std_logic;
  signal output_port_lookup_start_ack : std_logic;
  signal output_port_lookup_fin_req   : std_logic;
  signal output_port_lookup_fin_ack : std_logic;
  -- declarations related to module wrapper_input
  component wrapper_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(87 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(15 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(7 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(15 downto 0);
      free_queue_ack_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
      in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      start_wrapper_input_pipe_read_req : out  std_logic_vector(0 downto 0);
      start_wrapper_input_pipe_read_ack : in   std_logic_vector(0 downto 0);
      start_wrapper_input_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      midpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      midpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      midpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      last_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      last_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      last_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      pkt_length_pipe_write_req : out  std_logic_vector(0 downto 0);
      pkt_length_pipe_write_ack : in   std_logic_vector(0 downto 0);
      pkt_length_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_input
  signal wrapper_input_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_input_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic;
  signal wrapper_input_start_ack : std_logic;
  signal wrapper_input_fin_req   : std_logic;
  signal wrapper_input_fin_ack : std_logic;
  -- declarations related to module wrapper_output
  component wrapper_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_3_lr_req : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(87 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(15 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(7 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(15 downto 0);
      midpipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      midpipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      midpipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      last_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      last_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      last_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      pkt_length_pipe_read_req : out  std_logic_vector(0 downto 0);
      pkt_length_pipe_read_ack : in   std_logic_vector(0 downto 0);
      pkt_length_pipe_read_data : in   std_logic_vector(31 downto 0);
      start_wrapper_output_pipe_read_req : out  std_logic_vector(0 downto 0);
      start_wrapper_output_pipe_read_ack : in   std_logic_vector(0 downto 0);
      start_wrapper_output_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
      op_lut_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      op_lut_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      op_lut_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      op_lut_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_output
  signal wrapper_output_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_output_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic;
  signal wrapper_output_start_ack : std_logic;
  signal wrapper_output_fin_req   : std_logic;
  signal wrapper_output_fin_ack : std_logic;
  -- aggregate signals for write to pipe free_queue_ack
  signal free_queue_ack_pipe_write_data: std_logic_vector(7 downto 0);
  signal free_queue_ack_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_ack_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_ack
  signal free_queue_ack_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_ack_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_ack_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_get
  signal free_queue_get_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_get
  signal free_queue_get_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_put
  signal free_queue_put_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_put
  signal free_queue_put_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_request
  signal free_queue_request_pipe_write_data: std_logic_vector(15 downto 0);
  signal free_queue_request_pipe_write_req: std_logic_vector(1 downto 0);
  signal free_queue_request_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe free_queue_request
  signal free_queue_request_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_ctrl
  signal in_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe last_ctrl
  signal last_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal last_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal last_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe last_ctrl
  signal last_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal last_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal last_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe midpipe
  signal midpipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal midpipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal midpipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe midpipe
  signal midpipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal midpipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal midpipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe op_lut_ctrl
  signal op_lut_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal op_lut_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal op_lut_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe op_lut_ctrl
  signal op_lut_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal op_lut_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal op_lut_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe op_lut_data
  signal op_lut_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal op_lut_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal op_lut_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe op_lut_data
  signal op_lut_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal op_lut_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal op_lut_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_ctrl
  signal out_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe pkt_length
  signal pkt_length_pipe_write_data: std_logic_vector(31 downto 0);
  signal pkt_length_pipe_write_req: std_logic_vector(0 downto 0);
  signal pkt_length_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe pkt_length
  signal pkt_length_pipe_read_data: std_logic_vector(31 downto 0);
  signal pkt_length_pipe_read_req: std_logic_vector(0 downto 0);
  signal pkt_length_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe start_output_port_lookup
  signal start_output_port_lookup_pipe_write_data: std_logic_vector(7 downto 0);
  signal start_output_port_lookup_pipe_write_req: std_logic_vector(0 downto 0);
  signal start_output_port_lookup_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe start_output_port_lookup
  signal start_output_port_lookup_pipe_read_data: std_logic_vector(7 downto 0);
  signal start_output_port_lookup_pipe_read_req: std_logic_vector(0 downto 0);
  signal start_output_port_lookup_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe start_wrapper_input
  signal start_wrapper_input_pipe_write_data: std_logic_vector(7 downto 0);
  signal start_wrapper_input_pipe_write_req: std_logic_vector(0 downto 0);
  signal start_wrapper_input_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe start_wrapper_input
  signal start_wrapper_input_pipe_read_data: std_logic_vector(7 downto 0);
  signal start_wrapper_input_pipe_read_req: std_logic_vector(0 downto 0);
  signal start_wrapper_input_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe start_wrapper_output
  signal start_wrapper_output_pipe_write_data: std_logic_vector(7 downto 0);
  signal start_wrapper_output_pipe_write_req: std_logic_vector(0 downto 0);
  signal start_wrapper_output_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe start_wrapper_output
  signal start_wrapper_output_pipe_read_data: std_logic_vector(7 downto 0);
  signal start_wrapper_output_pipe_read_req: std_logic_vector(0 downto 0);
  signal start_wrapper_output_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module default_initializer_foo
  -- call arbiter for module default_initializer_foo
  default_initializer_foo_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_foo_call_reqs,
      call_acks => default_initializer_foo_call_acks,
      return_reqs => default_initializer_foo_return_reqs,
      return_acks => default_initializer_foo_return_acks,
      call_tag  => default_initializer_foo_call_tag,
      return_tag  => default_initializer_foo_return_tag,
      call_mtag => default_initializer_foo_tag_in,
      return_mtag => default_initializer_foo_tag_out,
      call_mreq => default_initializer_foo_start_req,
      call_mack => default_initializer_foo_start_ack,
      return_mreq => default_initializer_foo_fin_req,
      return_mack => default_initializer_foo_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_foo_instance:default_initializer_foo-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_foo_start_req,
      start_ack => default_initializer_foo_start_ack,
      fin_req => default_initializer_foo_fin_req,
      fin_ack => default_initializer_foo_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(1 downto 1),
      memory_space_1_sr_ack => memory_space_1_sr_ack(1 downto 1),
      memory_space_1_sr_addr => memory_space_1_sr_addr(7 downto 4),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 8),
      memory_space_1_sr_tag => memory_space_1_sr_tag(1 downto 1),
      memory_space_1_sc_req => memory_space_1_sc_req(1 downto 1),
      memory_space_1_sc_ack => memory_space_1_sc_ack(1 downto 1),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 1),
      tag_in => default_initializer_foo_tag_in,
      tag_out => default_initializer_foo_tag_out-- 
    ); -- 
  -- module default_initializer_free_queue
  -- call arbiter for module default_initializer_free_queue
  default_initializer_free_queue_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_free_queue_call_reqs,
      call_acks => default_initializer_free_queue_call_acks,
      return_reqs => default_initializer_free_queue_return_reqs,
      return_acks => default_initializer_free_queue_return_acks,
      call_tag  => default_initializer_free_queue_call_tag,
      return_tag  => default_initializer_free_queue_return_tag,
      call_mtag => default_initializer_free_queue_tag_in,
      return_mtag => default_initializer_free_queue_tag_out,
      call_mreq => default_initializer_free_queue_start_req,
      call_mack => default_initializer_free_queue_start_ack,
      return_mreq => default_initializer_free_queue_fin_req,
      return_mack => default_initializer_free_queue_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_free_queue_instance:default_initializer_free_queue-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_free_queue_start_req,
      start_ack => default_initializer_free_queue_start_ack,
      fin_req => default_initializer_free_queue_fin_req,
      fin_ack => default_initializer_free_queue_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(14 downto 12),
      memory_space_2_sr_data => memory_space_2_sr_data(39 downto 32),
      memory_space_2_sr_tag => memory_space_2_sr_tag(9 downto 8),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(9 downto 8),
      tag_in => default_initializer_free_queue_tag_in,
      tag_out => default_initializer_free_queue_tag_out-- 
    ); -- 
  -- module default_initializer_free_queue_ram
  -- call arbiter for module default_initializer_free_queue_ram
  default_initializer_free_queue_ram_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_free_queue_ram_call_reqs,
      call_acks => default_initializer_free_queue_ram_call_acks,
      return_reqs => default_initializer_free_queue_ram_return_reqs,
      return_acks => default_initializer_free_queue_ram_return_acks,
      call_tag  => default_initializer_free_queue_ram_call_tag,
      return_tag  => default_initializer_free_queue_ram_return_tag,
      call_mtag => default_initializer_free_queue_ram_tag_in,
      return_mtag => default_initializer_free_queue_ram_tag_out,
      call_mreq => default_initializer_free_queue_ram_start_req,
      call_mack => default_initializer_free_queue_ram_start_ack,
      return_mreq => default_initializer_free_queue_ram_fin_req,
      return_mack => default_initializer_free_queue_ram_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_free_queue_ram_instance:default_initializer_free_queue_ram-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_free_queue_ram_start_req,
      start_ack => default_initializer_free_queue_ram_start_ack,
      fin_req => default_initializer_free_queue_ram_fin_req,
      fin_ack => default_initializer_free_queue_ram_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_sr_req => memory_space_3_sr_req(8 downto 8),
      memory_space_3_sr_ack => memory_space_3_sr_ack(8 downto 8),
      memory_space_3_sr_addr => memory_space_3_sr_addr(98 downto 88),
      memory_space_3_sr_data => memory_space_3_sr_data(71 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(17 downto 16),
      memory_space_3_sc_req => memory_space_3_sc_req(8 downto 8),
      memory_space_3_sc_ack => memory_space_3_sc_ack(8 downto 8),
      memory_space_3_sc_tag => memory_space_3_sc_tag(17 downto 16),
      tag_in => default_initializer_free_queue_ram_tag_in,
      tag_out => default_initializer_free_queue_ram_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr
  -- call arbiter for module default_initializer_xx_xstr
  default_initializer_xx_xstr_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr_call_reqs,
      call_acks => default_initializer_xx_xstr_call_acks,
      return_reqs => default_initializer_xx_xstr_return_reqs,
      return_acks => default_initializer_xx_xstr_return_acks,
      call_tag  => default_initializer_xx_xstr_call_tag,
      return_tag  => default_initializer_xx_xstr_return_tag,
      call_mtag => default_initializer_xx_xstr_tag_in,
      return_mtag => default_initializer_xx_xstr_tag_out,
      call_mreq => default_initializer_xx_xstr_start_req,
      call_mack => default_initializer_xx_xstr_start_ack,
      return_mreq => default_initializer_xx_xstr_fin_req,
      return_mack => default_initializer_xx_xstr_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr_instance:default_initializer_xx_xstr-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr_start_req,
      start_ack => default_initializer_xx_xstr_start_ack,
      fin_req => default_initializer_xx_xstr_fin_req,
      fin_ack => default_initializer_xx_xstr_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(4 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(4 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(4 downto 0),
      tag_in => default_initializer_xx_xstr_tag_in,
      tag_out => default_initializer_xx_xstr_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr1
  -- call arbiter for module default_initializer_xx_xstr1
  default_initializer_xx_xstr1_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr1_call_reqs,
      call_acks => default_initializer_xx_xstr1_call_acks,
      return_reqs => default_initializer_xx_xstr1_return_reqs,
      return_acks => default_initializer_xx_xstr1_return_acks,
      call_tag  => default_initializer_xx_xstr1_call_tag,
      return_tag  => default_initializer_xx_xstr1_return_tag,
      call_mtag => default_initializer_xx_xstr1_tag_in,
      return_mtag => default_initializer_xx_xstr1_tag_out,
      call_mreq => default_initializer_xx_xstr1_start_req,
      call_mack => default_initializer_xx_xstr1_start_ack,
      return_mreq => default_initializer_xx_xstr1_fin_req,
      return_mack => default_initializer_xx_xstr1_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr1_instance:default_initializer_xx_xstr1-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr1_start_req,
      start_ack => default_initializer_xx_xstr1_start_ack,
      fin_req => default_initializer_xx_xstr1_fin_req,
      fin_ack => default_initializer_xx_xstr1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(3 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(7 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(3 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr1_tag_in,
      tag_out => default_initializer_xx_xstr1_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr10
  -- call arbiter for module default_initializer_xx_xstr10
  default_initializer_xx_xstr10_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr10_call_reqs,
      call_acks => default_initializer_xx_xstr10_call_acks,
      return_reqs => default_initializer_xx_xstr10_return_reqs,
      return_acks => default_initializer_xx_xstr10_return_acks,
      call_tag  => default_initializer_xx_xstr10_call_tag,
      return_tag  => default_initializer_xx_xstr10_return_tag,
      call_mtag => default_initializer_xx_xstr10_tag_in,
      return_mtag => default_initializer_xx_xstr10_tag_out,
      call_mreq => default_initializer_xx_xstr10_start_req,
      call_mack => default_initializer_xx_xstr10_start_ack,
      return_mreq => default_initializer_xx_xstr10_fin_req,
      return_mack => default_initializer_xx_xstr10_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr10_instance:default_initializer_xx_xstr10-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr10_start_req,
      start_ack => default_initializer_xx_xstr10_start_ack,
      fin_req => default_initializer_xx_xstr10_fin_req,
      fin_ack => default_initializer_xx_xstr10_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(4 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(7 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(4 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 0),
      tag_in => default_initializer_xx_xstr10_tag_in,
      tag_out => default_initializer_xx_xstr10_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr11
  -- call arbiter for module default_initializer_xx_xstr11
  default_initializer_xx_xstr11_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr11_call_reqs,
      call_acks => default_initializer_xx_xstr11_call_acks,
      return_reqs => default_initializer_xx_xstr11_return_reqs,
      return_acks => default_initializer_xx_xstr11_return_acks,
      call_tag  => default_initializer_xx_xstr11_call_tag,
      return_tag  => default_initializer_xx_xstr11_return_tag,
      call_mtag => default_initializer_xx_xstr11_tag_in,
      return_mtag => default_initializer_xx_xstr11_tag_out,
      call_mreq => default_initializer_xx_xstr11_start_req,
      call_mack => default_initializer_xx_xstr11_start_ack,
      return_mreq => default_initializer_xx_xstr11_fin_req,
      return_mack => default_initializer_xx_xstr11_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr11_instance:default_initializer_xx_xstr11-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr11_start_req,
      start_ack => default_initializer_xx_xstr11_start_ack,
      fin_req => default_initializer_xx_xstr11_fin_req,
      fin_ack => default_initializer_xx_xstr11_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(3 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(7 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(3 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr11_tag_in,
      tag_out => default_initializer_xx_xstr11_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr12
  -- call arbiter for module default_initializer_xx_xstr12
  default_initializer_xx_xstr12_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr12_call_reqs,
      call_acks => default_initializer_xx_xstr12_call_acks,
      return_reqs => default_initializer_xx_xstr12_return_reqs,
      return_acks => default_initializer_xx_xstr12_return_acks,
      call_tag  => default_initializer_xx_xstr12_call_tag,
      return_tag  => default_initializer_xx_xstr12_return_tag,
      call_mtag => default_initializer_xx_xstr12_tag_in,
      return_mtag => default_initializer_xx_xstr12_tag_out,
      call_mreq => default_initializer_xx_xstr12_start_req,
      call_mack => default_initializer_xx_xstr12_start_ack,
      return_mreq => default_initializer_xx_xstr12_fin_req,
      return_mack => default_initializer_xx_xstr12_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr12_instance:default_initializer_xx_xstr12-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr12_start_req,
      start_ack => default_initializer_xx_xstr12_start_ack,
      fin_req => default_initializer_xx_xstr12_fin_req,
      fin_ack => default_initializer_xx_xstr12_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(3 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(7 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(3 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr12_tag_in,
      tag_out => default_initializer_xx_xstr12_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr13
  -- call arbiter for module default_initializer_xx_xstr13
  default_initializer_xx_xstr13_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr13_call_reqs,
      call_acks => default_initializer_xx_xstr13_call_acks,
      return_reqs => default_initializer_xx_xstr13_return_reqs,
      return_acks => default_initializer_xx_xstr13_return_acks,
      call_tag  => default_initializer_xx_xstr13_call_tag,
      return_tag  => default_initializer_xx_xstr13_return_tag,
      call_mtag => default_initializer_xx_xstr13_tag_in,
      return_mtag => default_initializer_xx_xstr13_tag_out,
      call_mreq => default_initializer_xx_xstr13_start_req,
      call_mack => default_initializer_xx_xstr13_start_ack,
      return_mreq => default_initializer_xx_xstr13_fin_req,
      return_mack => default_initializer_xx_xstr13_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr13_instance:default_initializer_xx_xstr13-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr13_start_req,
      start_ack => default_initializer_xx_xstr13_start_ack,
      fin_req => default_initializer_xx_xstr13_fin_req,
      fin_ack => default_initializer_xx_xstr13_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_9_sr_req => memory_space_9_sr_req(0 downto 0),
      memory_space_9_sr_ack => memory_space_9_sr_ack(0 downto 0),
      memory_space_9_sr_addr => memory_space_9_sr_addr(3 downto 0),
      memory_space_9_sr_data => memory_space_9_sr_data(7 downto 0),
      memory_space_9_sr_tag => memory_space_9_sr_tag(3 downto 0),
      memory_space_9_sc_req => memory_space_9_sc_req(0 downto 0),
      memory_space_9_sc_ack => memory_space_9_sc_ack(0 downto 0),
      memory_space_9_sc_tag => memory_space_9_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr13_tag_in,
      tag_out => default_initializer_xx_xstr13_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr14
  -- call arbiter for module default_initializer_xx_xstr14
  default_initializer_xx_xstr14_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr14_call_reqs,
      call_acks => default_initializer_xx_xstr14_call_acks,
      return_reqs => default_initializer_xx_xstr14_return_reqs,
      return_acks => default_initializer_xx_xstr14_return_acks,
      call_tag  => default_initializer_xx_xstr14_call_tag,
      return_tag  => default_initializer_xx_xstr14_return_tag,
      call_mtag => default_initializer_xx_xstr14_tag_in,
      return_mtag => default_initializer_xx_xstr14_tag_out,
      call_mreq => default_initializer_xx_xstr14_start_req,
      call_mack => default_initializer_xx_xstr14_start_ack,
      return_mreq => default_initializer_xx_xstr14_fin_req,
      return_mack => default_initializer_xx_xstr14_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr14_instance:default_initializer_xx_xstr14-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr14_start_req,
      start_ack => default_initializer_xx_xstr14_start_ack,
      fin_req => default_initializer_xx_xstr14_fin_req,
      fin_ack => default_initializer_xx_xstr14_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_10_sr_req => memory_space_10_sr_req(0 downto 0),
      memory_space_10_sr_ack => memory_space_10_sr_ack(0 downto 0),
      memory_space_10_sr_addr => memory_space_10_sr_addr(3 downto 0),
      memory_space_10_sr_data => memory_space_10_sr_data(7 downto 0),
      memory_space_10_sr_tag => memory_space_10_sr_tag(3 downto 0),
      memory_space_10_sc_req => memory_space_10_sc_req(0 downto 0),
      memory_space_10_sc_ack => memory_space_10_sc_ack(0 downto 0),
      memory_space_10_sc_tag => memory_space_10_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr14_tag_in,
      tag_out => default_initializer_xx_xstr14_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr15
  -- call arbiter for module default_initializer_xx_xstr15
  default_initializer_xx_xstr15_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr15_call_reqs,
      call_acks => default_initializer_xx_xstr15_call_acks,
      return_reqs => default_initializer_xx_xstr15_return_reqs,
      return_acks => default_initializer_xx_xstr15_return_acks,
      call_tag  => default_initializer_xx_xstr15_call_tag,
      return_tag  => default_initializer_xx_xstr15_return_tag,
      call_mtag => default_initializer_xx_xstr15_tag_in,
      return_mtag => default_initializer_xx_xstr15_tag_out,
      call_mreq => default_initializer_xx_xstr15_start_req,
      call_mack => default_initializer_xx_xstr15_start_ack,
      return_mreq => default_initializer_xx_xstr15_fin_req,
      return_mack => default_initializer_xx_xstr15_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr15_instance:default_initializer_xx_xstr15-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr15_start_req,
      start_ack => default_initializer_xx_xstr15_start_ack,
      fin_req => default_initializer_xx_xstr15_fin_req,
      fin_ack => default_initializer_xx_xstr15_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_11_sr_req => memory_space_11_sr_req(0 downto 0),
      memory_space_11_sr_ack => memory_space_11_sr_ack(0 downto 0),
      memory_space_11_sr_addr => memory_space_11_sr_addr(3 downto 0),
      memory_space_11_sr_data => memory_space_11_sr_data(7 downto 0),
      memory_space_11_sr_tag => memory_space_11_sr_tag(3 downto 0),
      memory_space_11_sc_req => memory_space_11_sc_req(0 downto 0),
      memory_space_11_sc_ack => memory_space_11_sc_ack(0 downto 0),
      memory_space_11_sc_tag => memory_space_11_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr15_tag_in,
      tag_out => default_initializer_xx_xstr15_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr2
  -- call arbiter for module default_initializer_xx_xstr2
  default_initializer_xx_xstr2_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr2_call_reqs,
      call_acks => default_initializer_xx_xstr2_call_acks,
      return_reqs => default_initializer_xx_xstr2_return_reqs,
      return_acks => default_initializer_xx_xstr2_return_acks,
      call_tag  => default_initializer_xx_xstr2_call_tag,
      return_tag  => default_initializer_xx_xstr2_return_tag,
      call_mtag => default_initializer_xx_xstr2_tag_in,
      return_mtag => default_initializer_xx_xstr2_tag_out,
      call_mreq => default_initializer_xx_xstr2_start_req,
      call_mack => default_initializer_xx_xstr2_start_ack,
      return_mreq => default_initializer_xx_xstr2_fin_req,
      return_mack => default_initializer_xx_xstr2_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr2_instance:default_initializer_xx_xstr2-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr2_start_req,
      start_ack => default_initializer_xx_xstr2_start_ack,
      fin_req => default_initializer_xx_xstr2_fin_req,
      fin_ack => default_initializer_xx_xstr2_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_12_sr_req => memory_space_12_sr_req(0 downto 0),
      memory_space_12_sr_ack => memory_space_12_sr_ack(0 downto 0),
      memory_space_12_sr_addr => memory_space_12_sr_addr(3 downto 0),
      memory_space_12_sr_data => memory_space_12_sr_data(7 downto 0),
      memory_space_12_sr_tag => memory_space_12_sr_tag(3 downto 0),
      memory_space_12_sc_req => memory_space_12_sc_req(0 downto 0),
      memory_space_12_sc_ack => memory_space_12_sc_ack(0 downto 0),
      memory_space_12_sc_tag => memory_space_12_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr2_tag_in,
      tag_out => default_initializer_xx_xstr2_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr3
  -- call arbiter for module default_initializer_xx_xstr3
  default_initializer_xx_xstr3_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr3_call_reqs,
      call_acks => default_initializer_xx_xstr3_call_acks,
      return_reqs => default_initializer_xx_xstr3_return_reqs,
      return_acks => default_initializer_xx_xstr3_return_acks,
      call_tag  => default_initializer_xx_xstr3_call_tag,
      return_tag  => default_initializer_xx_xstr3_return_tag,
      call_mtag => default_initializer_xx_xstr3_tag_in,
      return_mtag => default_initializer_xx_xstr3_tag_out,
      call_mreq => default_initializer_xx_xstr3_start_req,
      call_mack => default_initializer_xx_xstr3_start_ack,
      return_mreq => default_initializer_xx_xstr3_fin_req,
      return_mack => default_initializer_xx_xstr3_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr3_instance:default_initializer_xx_xstr3-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr3_start_req,
      start_ack => default_initializer_xx_xstr3_start_ack,
      fin_req => default_initializer_xx_xstr3_fin_req,
      fin_ack => default_initializer_xx_xstr3_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_13_sr_req => memory_space_13_sr_req(0 downto 0),
      memory_space_13_sr_ack => memory_space_13_sr_ack(0 downto 0),
      memory_space_13_sr_addr => memory_space_13_sr_addr(3 downto 0),
      memory_space_13_sr_data => memory_space_13_sr_data(7 downto 0),
      memory_space_13_sr_tag => memory_space_13_sr_tag(3 downto 0),
      memory_space_13_sc_req => memory_space_13_sc_req(0 downto 0),
      memory_space_13_sc_ack => memory_space_13_sc_ack(0 downto 0),
      memory_space_13_sc_tag => memory_space_13_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr3_tag_in,
      tag_out => default_initializer_xx_xstr3_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr4
  -- call arbiter for module default_initializer_xx_xstr4
  default_initializer_xx_xstr4_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr4_call_reqs,
      call_acks => default_initializer_xx_xstr4_call_acks,
      return_reqs => default_initializer_xx_xstr4_return_reqs,
      return_acks => default_initializer_xx_xstr4_return_acks,
      call_tag  => default_initializer_xx_xstr4_call_tag,
      return_tag  => default_initializer_xx_xstr4_return_tag,
      call_mtag => default_initializer_xx_xstr4_tag_in,
      return_mtag => default_initializer_xx_xstr4_tag_out,
      call_mreq => default_initializer_xx_xstr4_start_req,
      call_mack => default_initializer_xx_xstr4_start_ack,
      return_mreq => default_initializer_xx_xstr4_fin_req,
      return_mack => default_initializer_xx_xstr4_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr4_instance:default_initializer_xx_xstr4-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr4_start_req,
      start_ack => default_initializer_xx_xstr4_start_ack,
      fin_req => default_initializer_xx_xstr4_fin_req,
      fin_ack => default_initializer_xx_xstr4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_14_sr_req => memory_space_14_sr_req(0 downto 0),
      memory_space_14_sr_ack => memory_space_14_sr_ack(0 downto 0),
      memory_space_14_sr_addr => memory_space_14_sr_addr(3 downto 0),
      memory_space_14_sr_data => memory_space_14_sr_data(7 downto 0),
      memory_space_14_sr_tag => memory_space_14_sr_tag(3 downto 0),
      memory_space_14_sc_req => memory_space_14_sc_req(0 downto 0),
      memory_space_14_sc_ack => memory_space_14_sc_ack(0 downto 0),
      memory_space_14_sc_tag => memory_space_14_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr4_tag_in,
      tag_out => default_initializer_xx_xstr4_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr5
  -- call arbiter for module default_initializer_xx_xstr5
  default_initializer_xx_xstr5_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr5_call_reqs,
      call_acks => default_initializer_xx_xstr5_call_acks,
      return_reqs => default_initializer_xx_xstr5_return_reqs,
      return_acks => default_initializer_xx_xstr5_return_acks,
      call_tag  => default_initializer_xx_xstr5_call_tag,
      return_tag  => default_initializer_xx_xstr5_return_tag,
      call_mtag => default_initializer_xx_xstr5_tag_in,
      return_mtag => default_initializer_xx_xstr5_tag_out,
      call_mreq => default_initializer_xx_xstr5_start_req,
      call_mack => default_initializer_xx_xstr5_start_ack,
      return_mreq => default_initializer_xx_xstr5_fin_req,
      return_mack => default_initializer_xx_xstr5_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr5_instance:default_initializer_xx_xstr5-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr5_start_req,
      start_ack => default_initializer_xx_xstr5_start_ack,
      fin_req => default_initializer_xx_xstr5_fin_req,
      fin_ack => default_initializer_xx_xstr5_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_15_sr_req => memory_space_15_sr_req(0 downto 0),
      memory_space_15_sr_ack => memory_space_15_sr_ack(0 downto 0),
      memory_space_15_sr_addr => memory_space_15_sr_addr(4 downto 0),
      memory_space_15_sr_data => memory_space_15_sr_data(7 downto 0),
      memory_space_15_sr_tag => memory_space_15_sr_tag(4 downto 0),
      memory_space_15_sc_req => memory_space_15_sc_req(0 downto 0),
      memory_space_15_sc_ack => memory_space_15_sc_ack(0 downto 0),
      memory_space_15_sc_tag => memory_space_15_sc_tag(4 downto 0),
      tag_in => default_initializer_xx_xstr5_tag_in,
      tag_out => default_initializer_xx_xstr5_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr6
  -- call arbiter for module default_initializer_xx_xstr6
  default_initializer_xx_xstr6_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr6_call_reqs,
      call_acks => default_initializer_xx_xstr6_call_acks,
      return_reqs => default_initializer_xx_xstr6_return_reqs,
      return_acks => default_initializer_xx_xstr6_return_acks,
      call_tag  => default_initializer_xx_xstr6_call_tag,
      return_tag  => default_initializer_xx_xstr6_return_tag,
      call_mtag => default_initializer_xx_xstr6_tag_in,
      return_mtag => default_initializer_xx_xstr6_tag_out,
      call_mreq => default_initializer_xx_xstr6_start_req,
      call_mack => default_initializer_xx_xstr6_start_ack,
      return_mreq => default_initializer_xx_xstr6_fin_req,
      return_mack => default_initializer_xx_xstr6_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr6_instance:default_initializer_xx_xstr6-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr6_start_req,
      start_ack => default_initializer_xx_xstr6_start_ack,
      fin_req => default_initializer_xx_xstr6_fin_req,
      fin_ack => default_initializer_xx_xstr6_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_16_sr_req => memory_space_16_sr_req(0 downto 0),
      memory_space_16_sr_ack => memory_space_16_sr_ack(0 downto 0),
      memory_space_16_sr_addr => memory_space_16_sr_addr(3 downto 0),
      memory_space_16_sr_data => memory_space_16_sr_data(7 downto 0),
      memory_space_16_sr_tag => memory_space_16_sr_tag(3 downto 0),
      memory_space_16_sc_req => memory_space_16_sc_req(0 downto 0),
      memory_space_16_sc_ack => memory_space_16_sc_ack(0 downto 0),
      memory_space_16_sc_tag => memory_space_16_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr6_tag_in,
      tag_out => default_initializer_xx_xstr6_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr7
  -- call arbiter for module default_initializer_xx_xstr7
  default_initializer_xx_xstr7_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr7_call_reqs,
      call_acks => default_initializer_xx_xstr7_call_acks,
      return_reqs => default_initializer_xx_xstr7_return_reqs,
      return_acks => default_initializer_xx_xstr7_return_acks,
      call_tag  => default_initializer_xx_xstr7_call_tag,
      return_tag  => default_initializer_xx_xstr7_return_tag,
      call_mtag => default_initializer_xx_xstr7_tag_in,
      return_mtag => default_initializer_xx_xstr7_tag_out,
      call_mreq => default_initializer_xx_xstr7_start_req,
      call_mack => default_initializer_xx_xstr7_start_ack,
      return_mreq => default_initializer_xx_xstr7_fin_req,
      return_mack => default_initializer_xx_xstr7_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr7_instance:default_initializer_xx_xstr7-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr7_start_req,
      start_ack => default_initializer_xx_xstr7_start_ack,
      fin_req => default_initializer_xx_xstr7_fin_req,
      fin_ack => default_initializer_xx_xstr7_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_17_sr_req => memory_space_17_sr_req(0 downto 0),
      memory_space_17_sr_ack => memory_space_17_sr_ack(0 downto 0),
      memory_space_17_sr_addr => memory_space_17_sr_addr(3 downto 0),
      memory_space_17_sr_data => memory_space_17_sr_data(7 downto 0),
      memory_space_17_sr_tag => memory_space_17_sr_tag(3 downto 0),
      memory_space_17_sc_req => memory_space_17_sc_req(0 downto 0),
      memory_space_17_sc_ack => memory_space_17_sc_ack(0 downto 0),
      memory_space_17_sc_tag => memory_space_17_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr7_tag_in,
      tag_out => default_initializer_xx_xstr7_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr8
  -- call arbiter for module default_initializer_xx_xstr8
  default_initializer_xx_xstr8_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr8_call_reqs,
      call_acks => default_initializer_xx_xstr8_call_acks,
      return_reqs => default_initializer_xx_xstr8_return_reqs,
      return_acks => default_initializer_xx_xstr8_return_acks,
      call_tag  => default_initializer_xx_xstr8_call_tag,
      return_tag  => default_initializer_xx_xstr8_return_tag,
      call_mtag => default_initializer_xx_xstr8_tag_in,
      return_mtag => default_initializer_xx_xstr8_tag_out,
      call_mreq => default_initializer_xx_xstr8_start_req,
      call_mack => default_initializer_xx_xstr8_start_ack,
      return_mreq => default_initializer_xx_xstr8_fin_req,
      return_mack => default_initializer_xx_xstr8_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr8_instance:default_initializer_xx_xstr8-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr8_start_req,
      start_ack => default_initializer_xx_xstr8_start_ack,
      fin_req => default_initializer_xx_xstr8_fin_req,
      fin_ack => default_initializer_xx_xstr8_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_18_sr_req => memory_space_18_sr_req(0 downto 0),
      memory_space_18_sr_ack => memory_space_18_sr_ack(0 downto 0),
      memory_space_18_sr_addr => memory_space_18_sr_addr(3 downto 0),
      memory_space_18_sr_data => memory_space_18_sr_data(7 downto 0),
      memory_space_18_sr_tag => memory_space_18_sr_tag(3 downto 0),
      memory_space_18_sc_req => memory_space_18_sc_req(0 downto 0),
      memory_space_18_sc_ack => memory_space_18_sc_ack(0 downto 0),
      memory_space_18_sc_tag => memory_space_18_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr8_tag_in,
      tag_out => default_initializer_xx_xstr8_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr9
  -- call arbiter for module default_initializer_xx_xstr9
  default_initializer_xx_xstr9_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr9_call_reqs,
      call_acks => default_initializer_xx_xstr9_call_acks,
      return_reqs => default_initializer_xx_xstr9_return_reqs,
      return_acks => default_initializer_xx_xstr9_return_acks,
      call_tag  => default_initializer_xx_xstr9_call_tag,
      return_tag  => default_initializer_xx_xstr9_return_tag,
      call_mtag => default_initializer_xx_xstr9_tag_in,
      return_mtag => default_initializer_xx_xstr9_tag_out,
      call_mreq => default_initializer_xx_xstr9_start_req,
      call_mack => default_initializer_xx_xstr9_start_ack,
      return_mreq => default_initializer_xx_xstr9_fin_req,
      return_mack => default_initializer_xx_xstr9_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr9_instance:default_initializer_xx_xstr9-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr9_start_req,
      start_ack => default_initializer_xx_xstr9_start_ack,
      fin_req => default_initializer_xx_xstr9_fin_req,
      fin_ack => default_initializer_xx_xstr9_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_19_sr_req => memory_space_19_sr_req(0 downto 0),
      memory_space_19_sr_ack => memory_space_19_sr_ack(0 downto 0),
      memory_space_19_sr_addr => memory_space_19_sr_addr(4 downto 0),
      memory_space_19_sr_data => memory_space_19_sr_data(7 downto 0),
      memory_space_19_sr_tag => memory_space_19_sr_tag(4 downto 0),
      memory_space_19_sc_req => memory_space_19_sc_req(0 downto 0),
      memory_space_19_sc_ack => memory_space_19_sc_ack(0 downto 0),
      memory_space_19_sc_tag => memory_space_19_sc_tag(4 downto 0),
      tag_in => default_initializer_xx_xstr9_tag_in,
      tag_out => default_initializer_xx_xstr9_tag_out-- 
    ); -- 
  -- module free_queue_manager
  free_queue_manager_instance:free_queue_manager-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => free_queue_manager_start_req,
      start_ack => free_queue_manager_start_ack,
      fin_req => free_queue_manager_fin_req,
      fin_ack => free_queue_manager_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(2 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(1 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(11 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(7 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(7 downto 0),
      free_queue_request_pipe_read_req => free_queue_request_pipe_read_req(0 downto 0),
      free_queue_request_pipe_read_ack => free_queue_request_pipe_read_ack(0 downto 0),
      free_queue_request_pipe_read_data => free_queue_request_pipe_read_data(7 downto 0),
      free_queue_put_pipe_read_req => free_queue_put_pipe_read_req(0 downto 0),
      free_queue_put_pipe_read_ack => free_queue_put_pipe_read_ack(0 downto 0),
      free_queue_put_pipe_read_data => free_queue_put_pipe_read_data(31 downto 0),
      free_queue_ack_pipe_write_req => free_queue_ack_pipe_write_req(0 downto 0),
      free_queue_ack_pipe_write_ack => free_queue_ack_pipe_write_ack(0 downto 0),
      free_queue_ack_pipe_write_data => free_queue_ack_pipe_write_data(7 downto 0),
      free_queue_get_pipe_write_req => free_queue_get_pipe_write_req(0 downto 0),
      free_queue_get_pipe_write_ack => free_queue_get_pipe_write_ack(0 downto 0),
      free_queue_get_pipe_write_data => free_queue_get_pipe_write_data(31 downto 0),
      start_output_port_lookup_pipe_write_req => start_output_port_lookup_pipe_write_req(0 downto 0),
      start_output_port_lookup_pipe_write_ack => start_output_port_lookup_pipe_write_ack(0 downto 0),
      start_output_port_lookup_pipe_write_data => start_output_port_lookup_pipe_write_data(7 downto 0),
      start_wrapper_input_pipe_write_req => start_wrapper_input_pipe_write_req(0 downto 0),
      start_wrapper_input_pipe_write_ack => start_wrapper_input_pipe_write_ack(0 downto 0),
      start_wrapper_input_pipe_write_data => start_wrapper_input_pipe_write_data(7 downto 0),
      start_wrapper_output_pipe_write_req => start_wrapper_output_pipe_write_req(0 downto 0),
      start_wrapper_output_pipe_write_ack => start_wrapper_output_pipe_write_ack(0 downto 0),
      start_wrapper_output_pipe_write_data => start_wrapper_output_pipe_write_data(7 downto 0),
      global_storage_initializer_x_call_reqs => global_storage_initializer_x_call_reqs(0 downto 0),
      global_storage_initializer_x_call_acks => global_storage_initializer_x_call_acks(0 downto 0),
      global_storage_initializer_x_call_tag => global_storage_initializer_x_call_tag(0 downto 0),
      global_storage_initializer_x_return_reqs => global_storage_initializer_x_return_reqs(0 downto 0),
      global_storage_initializer_x_return_acks => global_storage_initializer_x_return_acks(0 downto 0),
      global_storage_initializer_x_return_tag => global_storage_initializer_x_return_tag(0 downto 0),
      tag_in => free_queue_manager_tag_in,
      tag_out => free_queue_manager_tag_out-- 
    ); -- 
  -- module will be run forever 
  free_queue_manager_tag_in <= (others => '0');
  free_queue_manager_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => free_queue_manager_start_req, start_ack => free_queue_manager_start_ack,  fin_req => free_queue_manager_fin_req,  fin_ack => free_queue_manager_fin_ack);
  -- module global_storage_initializer_x
  -- call arbiter for module global_storage_initializer_x
  global_storage_initializer_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => global_storage_initializer_x_call_reqs,
      call_acks => global_storage_initializer_x_call_acks,
      return_reqs => global_storage_initializer_x_return_reqs,
      return_acks => global_storage_initializer_x_return_acks,
      call_tag  => global_storage_initializer_x_call_tag,
      return_tag  => global_storage_initializer_x_return_tag,
      call_mtag => global_storage_initializer_x_tag_in,
      return_mtag => global_storage_initializer_x_tag_out,
      call_mreq => global_storage_initializer_x_start_req,
      call_mack => global_storage_initializer_x_start_ack,
      return_mreq => global_storage_initializer_x_fin_req,
      return_mack => global_storage_initializer_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  global_storage_initializer_x_instance:global_storage_initializer_x-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => global_storage_initializer_x_start_req,
      start_ack => global_storage_initializer_x_start_ack,
      fin_req => global_storage_initializer_x_fin_req,
      fin_ack => global_storage_initializer_x_fin_ack,
      clk => clk,
      reset => reset,
      default_initializer_foo_call_reqs => default_initializer_foo_call_reqs(0 downto 0),
      default_initializer_foo_call_acks => default_initializer_foo_call_acks(0 downto 0),
      default_initializer_foo_call_tag => default_initializer_foo_call_tag(0 downto 0),
      default_initializer_foo_return_reqs => default_initializer_foo_return_reqs(0 downto 0),
      default_initializer_foo_return_acks => default_initializer_foo_return_acks(0 downto 0),
      default_initializer_foo_return_tag => default_initializer_foo_return_tag(0 downto 0),
      default_initializer_free_queue_call_reqs => default_initializer_free_queue_call_reqs(0 downto 0),
      default_initializer_free_queue_call_acks => default_initializer_free_queue_call_acks(0 downto 0),
      default_initializer_free_queue_call_tag => default_initializer_free_queue_call_tag(0 downto 0),
      default_initializer_free_queue_return_reqs => default_initializer_free_queue_return_reqs(0 downto 0),
      default_initializer_free_queue_return_acks => default_initializer_free_queue_return_acks(0 downto 0),
      default_initializer_free_queue_return_tag => default_initializer_free_queue_return_tag(0 downto 0),
      default_initializer_free_queue_ram_call_reqs => default_initializer_free_queue_ram_call_reqs(0 downto 0),
      default_initializer_free_queue_ram_call_acks => default_initializer_free_queue_ram_call_acks(0 downto 0),
      default_initializer_free_queue_ram_call_tag => default_initializer_free_queue_ram_call_tag(0 downto 0),
      default_initializer_free_queue_ram_return_reqs => default_initializer_free_queue_ram_return_reqs(0 downto 0),
      default_initializer_free_queue_ram_return_acks => default_initializer_free_queue_ram_return_acks(0 downto 0),
      default_initializer_free_queue_ram_return_tag => default_initializer_free_queue_ram_return_tag(0 downto 0),
      default_initializer_xx_xstr_call_reqs => default_initializer_xx_xstr_call_reqs(0 downto 0),
      default_initializer_xx_xstr_call_acks => default_initializer_xx_xstr_call_acks(0 downto 0),
      default_initializer_xx_xstr_call_tag => default_initializer_xx_xstr_call_tag(0 downto 0),
      default_initializer_xx_xstr_return_reqs => default_initializer_xx_xstr_return_reqs(0 downto 0),
      default_initializer_xx_xstr_return_acks => default_initializer_xx_xstr_return_acks(0 downto 0),
      default_initializer_xx_xstr_return_tag => default_initializer_xx_xstr_return_tag(0 downto 0),
      default_initializer_xx_xstr1_call_reqs => default_initializer_xx_xstr1_call_reqs(0 downto 0),
      default_initializer_xx_xstr1_call_acks => default_initializer_xx_xstr1_call_acks(0 downto 0),
      default_initializer_xx_xstr1_call_tag => default_initializer_xx_xstr1_call_tag(0 downto 0),
      default_initializer_xx_xstr1_return_reqs => default_initializer_xx_xstr1_return_reqs(0 downto 0),
      default_initializer_xx_xstr1_return_acks => default_initializer_xx_xstr1_return_acks(0 downto 0),
      default_initializer_xx_xstr1_return_tag => default_initializer_xx_xstr1_return_tag(0 downto 0),
      default_initializer_xx_xstr10_call_reqs => default_initializer_xx_xstr10_call_reqs(0 downto 0),
      default_initializer_xx_xstr10_call_acks => default_initializer_xx_xstr10_call_acks(0 downto 0),
      default_initializer_xx_xstr10_call_tag => default_initializer_xx_xstr10_call_tag(0 downto 0),
      default_initializer_xx_xstr10_return_reqs => default_initializer_xx_xstr10_return_reqs(0 downto 0),
      default_initializer_xx_xstr10_return_acks => default_initializer_xx_xstr10_return_acks(0 downto 0),
      default_initializer_xx_xstr10_return_tag => default_initializer_xx_xstr10_return_tag(0 downto 0),
      default_initializer_xx_xstr11_call_reqs => default_initializer_xx_xstr11_call_reqs(0 downto 0),
      default_initializer_xx_xstr11_call_acks => default_initializer_xx_xstr11_call_acks(0 downto 0),
      default_initializer_xx_xstr11_call_tag => default_initializer_xx_xstr11_call_tag(0 downto 0),
      default_initializer_xx_xstr11_return_reqs => default_initializer_xx_xstr11_return_reqs(0 downto 0),
      default_initializer_xx_xstr11_return_acks => default_initializer_xx_xstr11_return_acks(0 downto 0),
      default_initializer_xx_xstr11_return_tag => default_initializer_xx_xstr11_return_tag(0 downto 0),
      default_initializer_xx_xstr12_call_reqs => default_initializer_xx_xstr12_call_reqs(0 downto 0),
      default_initializer_xx_xstr12_call_acks => default_initializer_xx_xstr12_call_acks(0 downto 0),
      default_initializer_xx_xstr12_call_tag => default_initializer_xx_xstr12_call_tag(0 downto 0),
      default_initializer_xx_xstr12_return_reqs => default_initializer_xx_xstr12_return_reqs(0 downto 0),
      default_initializer_xx_xstr12_return_acks => default_initializer_xx_xstr12_return_acks(0 downto 0),
      default_initializer_xx_xstr12_return_tag => default_initializer_xx_xstr12_return_tag(0 downto 0),
      default_initializer_xx_xstr13_call_reqs => default_initializer_xx_xstr13_call_reqs(0 downto 0),
      default_initializer_xx_xstr13_call_acks => default_initializer_xx_xstr13_call_acks(0 downto 0),
      default_initializer_xx_xstr13_call_tag => default_initializer_xx_xstr13_call_tag(0 downto 0),
      default_initializer_xx_xstr13_return_reqs => default_initializer_xx_xstr13_return_reqs(0 downto 0),
      default_initializer_xx_xstr13_return_acks => default_initializer_xx_xstr13_return_acks(0 downto 0),
      default_initializer_xx_xstr13_return_tag => default_initializer_xx_xstr13_return_tag(0 downto 0),
      default_initializer_xx_xstr14_call_reqs => default_initializer_xx_xstr14_call_reqs(0 downto 0),
      default_initializer_xx_xstr14_call_acks => default_initializer_xx_xstr14_call_acks(0 downto 0),
      default_initializer_xx_xstr14_call_tag => default_initializer_xx_xstr14_call_tag(0 downto 0),
      default_initializer_xx_xstr14_return_reqs => default_initializer_xx_xstr14_return_reqs(0 downto 0),
      default_initializer_xx_xstr14_return_acks => default_initializer_xx_xstr14_return_acks(0 downto 0),
      default_initializer_xx_xstr14_return_tag => default_initializer_xx_xstr14_return_tag(0 downto 0),
      default_initializer_xx_xstr15_call_reqs => default_initializer_xx_xstr15_call_reqs(0 downto 0),
      default_initializer_xx_xstr15_call_acks => default_initializer_xx_xstr15_call_acks(0 downto 0),
      default_initializer_xx_xstr15_call_tag => default_initializer_xx_xstr15_call_tag(0 downto 0),
      default_initializer_xx_xstr15_return_reqs => default_initializer_xx_xstr15_return_reqs(0 downto 0),
      default_initializer_xx_xstr15_return_acks => default_initializer_xx_xstr15_return_acks(0 downto 0),
      default_initializer_xx_xstr15_return_tag => default_initializer_xx_xstr15_return_tag(0 downto 0),
      default_initializer_xx_xstr2_call_reqs => default_initializer_xx_xstr2_call_reqs(0 downto 0),
      default_initializer_xx_xstr2_call_acks => default_initializer_xx_xstr2_call_acks(0 downto 0),
      default_initializer_xx_xstr2_call_tag => default_initializer_xx_xstr2_call_tag(0 downto 0),
      default_initializer_xx_xstr2_return_reqs => default_initializer_xx_xstr2_return_reqs(0 downto 0),
      default_initializer_xx_xstr2_return_acks => default_initializer_xx_xstr2_return_acks(0 downto 0),
      default_initializer_xx_xstr2_return_tag => default_initializer_xx_xstr2_return_tag(0 downto 0),
      default_initializer_xx_xstr3_call_reqs => default_initializer_xx_xstr3_call_reqs(0 downto 0),
      default_initializer_xx_xstr3_call_acks => default_initializer_xx_xstr3_call_acks(0 downto 0),
      default_initializer_xx_xstr3_call_tag => default_initializer_xx_xstr3_call_tag(0 downto 0),
      default_initializer_xx_xstr3_return_reqs => default_initializer_xx_xstr3_return_reqs(0 downto 0),
      default_initializer_xx_xstr3_return_acks => default_initializer_xx_xstr3_return_acks(0 downto 0),
      default_initializer_xx_xstr3_return_tag => default_initializer_xx_xstr3_return_tag(0 downto 0),
      default_initializer_xx_xstr4_call_reqs => default_initializer_xx_xstr4_call_reqs(0 downto 0),
      default_initializer_xx_xstr4_call_acks => default_initializer_xx_xstr4_call_acks(0 downto 0),
      default_initializer_xx_xstr4_call_tag => default_initializer_xx_xstr4_call_tag(0 downto 0),
      default_initializer_xx_xstr4_return_reqs => default_initializer_xx_xstr4_return_reqs(0 downto 0),
      default_initializer_xx_xstr4_return_acks => default_initializer_xx_xstr4_return_acks(0 downto 0),
      default_initializer_xx_xstr4_return_tag => default_initializer_xx_xstr4_return_tag(0 downto 0),
      default_initializer_xx_xstr5_call_reqs => default_initializer_xx_xstr5_call_reqs(0 downto 0),
      default_initializer_xx_xstr5_call_acks => default_initializer_xx_xstr5_call_acks(0 downto 0),
      default_initializer_xx_xstr5_call_tag => default_initializer_xx_xstr5_call_tag(0 downto 0),
      default_initializer_xx_xstr5_return_reqs => default_initializer_xx_xstr5_return_reqs(0 downto 0),
      default_initializer_xx_xstr5_return_acks => default_initializer_xx_xstr5_return_acks(0 downto 0),
      default_initializer_xx_xstr5_return_tag => default_initializer_xx_xstr5_return_tag(0 downto 0),
      default_initializer_xx_xstr6_call_reqs => default_initializer_xx_xstr6_call_reqs(0 downto 0),
      default_initializer_xx_xstr6_call_acks => default_initializer_xx_xstr6_call_acks(0 downto 0),
      default_initializer_xx_xstr6_call_tag => default_initializer_xx_xstr6_call_tag(0 downto 0),
      default_initializer_xx_xstr6_return_reqs => default_initializer_xx_xstr6_return_reqs(0 downto 0),
      default_initializer_xx_xstr6_return_acks => default_initializer_xx_xstr6_return_acks(0 downto 0),
      default_initializer_xx_xstr6_return_tag => default_initializer_xx_xstr6_return_tag(0 downto 0),
      default_initializer_xx_xstr7_call_reqs => default_initializer_xx_xstr7_call_reqs(0 downto 0),
      default_initializer_xx_xstr7_call_acks => default_initializer_xx_xstr7_call_acks(0 downto 0),
      default_initializer_xx_xstr7_call_tag => default_initializer_xx_xstr7_call_tag(0 downto 0),
      default_initializer_xx_xstr7_return_reqs => default_initializer_xx_xstr7_return_reqs(0 downto 0),
      default_initializer_xx_xstr7_return_acks => default_initializer_xx_xstr7_return_acks(0 downto 0),
      default_initializer_xx_xstr7_return_tag => default_initializer_xx_xstr7_return_tag(0 downto 0),
      default_initializer_xx_xstr8_call_reqs => default_initializer_xx_xstr8_call_reqs(0 downto 0),
      default_initializer_xx_xstr8_call_acks => default_initializer_xx_xstr8_call_acks(0 downto 0),
      default_initializer_xx_xstr8_call_tag => default_initializer_xx_xstr8_call_tag(0 downto 0),
      default_initializer_xx_xstr8_return_reqs => default_initializer_xx_xstr8_return_reqs(0 downto 0),
      default_initializer_xx_xstr8_return_acks => default_initializer_xx_xstr8_return_acks(0 downto 0),
      default_initializer_xx_xstr8_return_tag => default_initializer_xx_xstr8_return_tag(0 downto 0),
      default_initializer_xx_xstr9_call_reqs => default_initializer_xx_xstr9_call_reqs(0 downto 0),
      default_initializer_xx_xstr9_call_acks => default_initializer_xx_xstr9_call_acks(0 downto 0),
      default_initializer_xx_xstr9_call_tag => default_initializer_xx_xstr9_call_tag(0 downto 0),
      default_initializer_xx_xstr9_return_reqs => default_initializer_xx_xstr9_return_reqs(0 downto 0),
      default_initializer_xx_xstr9_return_acks => default_initializer_xx_xstr9_return_acks(0 downto 0),
      default_initializer_xx_xstr9_return_tag => default_initializer_xx_xstr9_return_tag(0 downto 0),
      tag_in => global_storage_initializer_x_tag_in,
      tag_out => global_storage_initializer_x_tag_out-- 
    ); -- 
  -- module output_port_lookup
  output_port_lookup_instance:output_port_lookup-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => output_port_lookup_start_req,
      start_ack => output_port_lookup_start_ack,
      fin_req => output_port_lookup_fin_req,
      fin_ack => output_port_lookup_fin_ack,
      clk => clk,
      reset => reset,
      op_lut_ctrl_pipe_read_req => op_lut_ctrl_pipe_read_req(0 downto 0),
      op_lut_ctrl_pipe_read_ack => op_lut_ctrl_pipe_read_ack(0 downto 0),
      op_lut_ctrl_pipe_read_data => op_lut_ctrl_pipe_read_data(7 downto 0),
      op_lut_data_pipe_read_req => op_lut_data_pipe_read_req(0 downto 0),
      op_lut_data_pipe_read_ack => op_lut_data_pipe_read_ack(0 downto 0),
      op_lut_data_pipe_read_data => op_lut_data_pipe_read_data(63 downto 0),
      start_output_port_lookup_pipe_read_req => start_output_port_lookup_pipe_read_req(0 downto 0),
      start_output_port_lookup_pipe_read_ack => start_output_port_lookup_pipe_read_ack(0 downto 0),
      start_output_port_lookup_pipe_read_data => start_output_port_lookup_pipe_read_data(7 downto 0),
      out_ctrl_pipe_write_req => out_ctrl_pipe_write_req(0 downto 0),
      out_ctrl_pipe_write_ack => out_ctrl_pipe_write_ack(0 downto 0),
      out_ctrl_pipe_write_data => out_ctrl_pipe_write_data(7 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      tag_in => output_port_lookup_tag_in,
      tag_out => output_port_lookup_tag_out-- 
    ); -- 
  -- module will be run forever 
  output_port_lookup_tag_in <= (others => '0');
  output_port_lookup_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => output_port_lookup_start_req, start_ack => output_port_lookup_start_ack,  fin_req => output_port_lookup_fin_req,  fin_ack => output_port_lookup_fin_ack);
  -- module wrapper_input
  wrapper_input_instance:wrapper_input-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_input_start_req,
      start_ack => wrapper_input_start_ack,
      fin_req => wrapper_input_fin_req,
      fin_ack => wrapper_input_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(3 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(7 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(7 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(7 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(87 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(15 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(7 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(7 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(15 downto 0),
      free_queue_ack_pipe_read_req => free_queue_ack_pipe_read_req(0 downto 0),
      free_queue_ack_pipe_read_ack => free_queue_ack_pipe_read_ack(0 downto 0),
      free_queue_ack_pipe_read_data => free_queue_ack_pipe_read_data(7 downto 0),
      free_queue_get_pipe_read_req => free_queue_get_pipe_read_req(0 downto 0),
      free_queue_get_pipe_read_ack => free_queue_get_pipe_read_ack(0 downto 0),
      free_queue_get_pipe_read_data => free_queue_get_pipe_read_data(31 downto 0),
      in_ctrl_pipe_read_req => in_ctrl_pipe_read_req(0 downto 0),
      in_ctrl_pipe_read_ack => in_ctrl_pipe_read_ack(0 downto 0),
      in_ctrl_pipe_read_data => in_ctrl_pipe_read_data(7 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      start_wrapper_input_pipe_read_req => start_wrapper_input_pipe_read_req(0 downto 0),
      start_wrapper_input_pipe_read_ack => start_wrapper_input_pipe_read_ack(0 downto 0),
      start_wrapper_input_pipe_read_data => start_wrapper_input_pipe_read_data(7 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(1 downto 1),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(1 downto 1),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(15 downto 8),
      midpipe_pipe_write_req => midpipe_pipe_write_req(0 downto 0),
      midpipe_pipe_write_ack => midpipe_pipe_write_ack(0 downto 0),
      midpipe_pipe_write_data => midpipe_pipe_write_data(31 downto 0),
      last_ctrl_pipe_write_req => last_ctrl_pipe_write_req(0 downto 0),
      last_ctrl_pipe_write_ack => last_ctrl_pipe_write_ack(0 downto 0),
      last_ctrl_pipe_write_data => last_ctrl_pipe_write_data(7 downto 0),
      pkt_length_pipe_write_req => pkt_length_pipe_write_req(0 downto 0),
      pkt_length_pipe_write_ack => pkt_length_pipe_write_ack(0 downto 0),
      pkt_length_pipe_write_data => pkt_length_pipe_write_data(31 downto 0),
      tag_in => wrapper_input_tag_in,
      tag_out => wrapper_input_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_input_tag_in <= (others => '0');
  wrapper_input_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_input_start_req, start_ack => wrapper_input_start_ack,  fin_req => wrapper_input_fin_req,  fin_ack => wrapper_input_fin_ack);
  -- module wrapper_output
  wrapper_output_instance:wrapper_output-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_output_start_req,
      start_ack => wrapper_output_start_ack,
      fin_req => wrapper_output_fin_req,
      fin_ack => wrapper_output_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(7 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(7 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(87 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(15 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(7 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(7 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(15 downto 0),
      midpipe_pipe_read_req => midpipe_pipe_read_req(0 downto 0),
      midpipe_pipe_read_ack => midpipe_pipe_read_ack(0 downto 0),
      midpipe_pipe_read_data => midpipe_pipe_read_data(31 downto 0),
      last_ctrl_pipe_read_req => last_ctrl_pipe_read_req(0 downto 0),
      last_ctrl_pipe_read_ack => last_ctrl_pipe_read_ack(0 downto 0),
      last_ctrl_pipe_read_data => last_ctrl_pipe_read_data(7 downto 0),
      pkt_length_pipe_read_req => pkt_length_pipe_read_req(0 downto 0),
      pkt_length_pipe_read_ack => pkt_length_pipe_read_ack(0 downto 0),
      pkt_length_pipe_read_data => pkt_length_pipe_read_data(31 downto 0),
      start_wrapper_output_pipe_read_req => start_wrapper_output_pipe_read_req(0 downto 0),
      start_wrapper_output_pipe_read_ack => start_wrapper_output_pipe_read_ack(0 downto 0),
      start_wrapper_output_pipe_read_data => start_wrapper_output_pipe_read_data(7 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(0 downto 0),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(0 downto 0),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(7 downto 0),
      free_queue_put_pipe_write_req => free_queue_put_pipe_write_req(0 downto 0),
      free_queue_put_pipe_write_ack => free_queue_put_pipe_write_ack(0 downto 0),
      free_queue_put_pipe_write_data => free_queue_put_pipe_write_data(31 downto 0),
      op_lut_ctrl_pipe_write_req => op_lut_ctrl_pipe_write_req(0 downto 0),
      op_lut_ctrl_pipe_write_ack => op_lut_ctrl_pipe_write_ack(0 downto 0),
      op_lut_ctrl_pipe_write_data => op_lut_ctrl_pipe_write_data(7 downto 0),
      op_lut_data_pipe_write_req => op_lut_data_pipe_write_req(0 downto 0),
      op_lut_data_pipe_write_ack => op_lut_data_pipe_write_ack(0 downto 0),
      op_lut_data_pipe_write_data => op_lut_data_pipe_write_data(63 downto 0),
      tag_in => wrapper_output_tag_in,
      tag_out => wrapper_output_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_output_tag_in <= (others => '0');
  wrapper_output_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_output_start_req, start_ack => wrapper_output_start_ack,  fin_req => wrapper_output_fin_req,  fin_ack => wrapper_output_fin_ack);
  free_queue_ack_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_ack_pipe_read_req,
      read_ack => free_queue_ack_pipe_read_ack,
      read_data => free_queue_ack_pipe_read_data,
      write_req => free_queue_ack_pipe_write_req,
      write_ack => free_queue_ack_pipe_write_ack,
      write_data => free_queue_ack_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_get_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_get_pipe_read_req,
      read_ack => free_queue_get_pipe_read_ack,
      read_data => free_queue_get_pipe_read_data,
      write_req => free_queue_get_pipe_write_req,
      write_ack => free_queue_get_pipe_write_ack,
      write_data => free_queue_get_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_put_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_put_pipe_read_req,
      read_ack => free_queue_put_pipe_read_ack,
      read_data => free_queue_put_pipe_read_data,
      write_req => free_queue_put_pipe_write_req,
      write_ack => free_queue_put_pipe_write_ack,
      write_data => free_queue_put_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_request_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_request_pipe_read_req,
      read_ack => free_queue_request_pipe_read_ack,
      read_data => free_queue_request_pipe_read_data,
      write_req => free_queue_request_pipe_write_req,
      write_ack => free_queue_request_pipe_write_ack,
      write_data => free_queue_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => in_ctrl_pipe_read_req,
      read_ack => in_ctrl_pipe_read_ack,
      read_data => in_ctrl_pipe_read_data,
      write_req => in_ctrl_pipe_write_req,
      write_ack => in_ctrl_pipe_write_ack,
      write_data => in_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  last_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => last_ctrl_pipe_read_req,
      read_ack => last_ctrl_pipe_read_ack,
      read_data => last_ctrl_pipe_read_data,
      write_req => last_ctrl_pipe_write_req,
      write_ack => last_ctrl_pipe_write_ack,
      write_data => last_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  midpipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => midpipe_pipe_read_req,
      read_ack => midpipe_pipe_read_ack,
      read_data => midpipe_pipe_read_data,
      write_req => midpipe_pipe_write_req,
      write_ack => midpipe_pipe_write_ack,
      write_data => midpipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  op_lut_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => op_lut_ctrl_pipe_read_req,
      read_ack => op_lut_ctrl_pipe_read_ack,
      read_data => op_lut_ctrl_pipe_read_data,
      write_req => op_lut_ctrl_pipe_write_req,
      write_ack => op_lut_ctrl_pipe_write_ack,
      write_data => op_lut_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  op_lut_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => op_lut_data_pipe_read_req,
      read_ack => op_lut_data_pipe_read_ack,
      read_data => op_lut_data_pipe_read_data,
      write_req => op_lut_data_pipe_write_req,
      write_ack => op_lut_data_pipe_write_ack,
      write_data => op_lut_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => out_ctrl_pipe_read_req,
      read_ack => out_ctrl_pipe_read_ack,
      read_data => out_ctrl_pipe_read_data,
      write_req => out_ctrl_pipe_write_req,
      write_ack => out_ctrl_pipe_write_ack,
      write_data => out_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  pkt_length_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => pkt_length_pipe_read_req,
      read_ack => pkt_length_pipe_read_ack,
      read_data => pkt_length_pipe_read_data,
      write_req => pkt_length_pipe_write_req,
      write_ack => pkt_length_pipe_write_ack,
      write_data => pkt_length_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  start_output_port_lookup_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => start_output_port_lookup_pipe_read_req,
      read_ack => start_output_port_lookup_pipe_read_ack,
      read_data => start_output_port_lookup_pipe_read_data,
      write_req => start_output_port_lookup_pipe_write_req,
      write_ack => start_output_port_lookup_pipe_write_ack,
      write_data => start_output_port_lookup_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  start_wrapper_input_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => start_wrapper_input_pipe_read_req,
      read_ack => start_wrapper_input_pipe_read_ack,
      read_data => start_wrapper_input_pipe_read_data,
      write_req => start_wrapper_input_pipe_write_req,
      write_ack => start_wrapper_input_pipe_write_ack,
      write_data => start_wrapper_input_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  start_wrapper_output_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => start_wrapper_output_pipe_read_req,
      read_ack => start_wrapper_output_pipe_read_ack,
      read_data => start_wrapper_output_pipe_read_data,
      write_req => start_wrapper_output_pipe_write_req,
      write_ack => start_wrapper_output_pipe_write_ack,
      write_data => start_wrapper_output_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 2,
      addr_width => 4,
      data_width => 8,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_10: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_11: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_11_sr_addr,
      sr_data_in => memory_space_11_sr_data,
      sr_req_in => memory_space_11_sr_req,
      sr_ack_out => memory_space_11_sr_ack,
      sr_tag_in => memory_space_11_sr_tag,
      sc_req_in=> memory_space_11_sc_req,
      sc_ack_out => memory_space_11_sc_ack,
      sc_tag_out => memory_space_11_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_12: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_12_sr_addr,
      sr_data_in => memory_space_12_sr_data,
      sr_req_in => memory_space_12_sr_req,
      sr_ack_out => memory_space_12_sr_ack,
      sr_tag_in => memory_space_12_sr_tag,
      sc_req_in=> memory_space_12_sc_req,
      sc_ack_out => memory_space_12_sc_ack,
      sc_tag_out => memory_space_12_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_13: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_13_sr_addr,
      sr_data_in => memory_space_13_sr_data,
      sr_req_in => memory_space_13_sr_req,
      sr_ack_out => memory_space_13_sr_ack,
      sr_tag_in => memory_space_13_sr_tag,
      sc_req_in=> memory_space_13_sc_req,
      sc_ack_out => memory_space_13_sc_ack,
      sc_tag_out => memory_space_13_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_14: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_14_sr_addr,
      sr_data_in => memory_space_14_sr_data,
      sr_req_in => memory_space_14_sr_req,
      sr_ack_out => memory_space_14_sr_ack,
      sr_tag_in => memory_space_14_sr_tag,
      sc_req_in=> memory_space_14_sc_req,
      sc_ack_out => memory_space_14_sc_ack,
      sc_tag_out => memory_space_14_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_15: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 5,
      data_width => 8,
      tag_width => 5
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_15_sr_addr,
      sr_data_in => memory_space_15_sr_data,
      sr_req_in => memory_space_15_sr_req,
      sr_ack_out => memory_space_15_sr_ack,
      sr_tag_in => memory_space_15_sr_tag,
      sc_req_in=> memory_space_15_sc_req,
      sc_ack_out => memory_space_15_sc_ack,
      sc_tag_out => memory_space_15_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_16: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_16_sr_addr,
      sr_data_in => memory_space_16_sr_data,
      sr_req_in => memory_space_16_sr_req,
      sr_ack_out => memory_space_16_sr_ack,
      sr_tag_in => memory_space_16_sr_tag,
      sc_req_in=> memory_space_16_sc_req,
      sc_ack_out => memory_space_16_sc_ack,
      sc_tag_out => memory_space_16_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_17: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_17_sr_addr,
      sr_data_in => memory_space_17_sr_data,
      sr_req_in => memory_space_17_sr_req,
      sr_ack_out => memory_space_17_sr_ack,
      sr_tag_in => memory_space_17_sr_tag,
      sc_req_in=> memory_space_17_sc_req,
      sc_ack_out => memory_space_17_sc_ack,
      sc_tag_out => memory_space_17_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_18: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_18_sr_addr,
      sr_data_in => memory_space_18_sr_data,
      sr_req_in => memory_space_18_sr_req,
      sr_ack_out => memory_space_18_sr_ack,
      sr_tag_in => memory_space_18_sr_tag,
      sc_req_in=> memory_space_18_sc_req,
      sc_ack_out => memory_space_18_sc_ack,
      sc_tag_out => memory_space_18_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_19: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 5,
      data_width => 8,
      tag_width => 5
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_19_sr_addr,
      sr_data_in => memory_space_19_sr_data,
      sr_req_in => memory_space_19_sr_req,
      sr_ack_out => memory_space_19_sr_ack,
      sr_tag_in => memory_space_19_sr_tag,
      sc_req_in=> memory_space_19_sc_req,
      sc_ack_out => memory_space_19_sc_ack,
      sc_tag_out => memory_space_19_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_2: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 5,
      addr_width => 3,
      data_width => 8,
      tag_width => 2,
      num_registers => 4) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: memory_subsystem -- 
    generic map(-- 
      num_loads => 8,
      num_stores => 9,
      addr_width => 11,
      data_width => 8,
      tag_width => 2,
      number_of_banks => 4,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_4: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 5,
      data_width => 8,
      tag_width => 5
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_6: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 5,
      data_width => 8,
      tag_width => 5
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_7: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_8: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_9: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
