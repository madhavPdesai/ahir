-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity maxOfTwo is -- 
  generic (tag_length : integer); 
  port ( -- 
    a : in  std_logic_vector(31 downto 0);
    b : in  std_logic_vector(31 downto 0);
    ret_val_x_x : out  std_logic_vector(31 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity maxOfTwo;
architecture Default of maxOfTwo is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal a_buffer :  std_logic_vector(31 downto 0);
  signal a_update_enable: Boolean;
  signal b_buffer :  std_logic_vector(31 downto 0);
  signal b_update_enable: Boolean;
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(31 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal maxOfTwo_CP_0_start: Boolean;
  signal maxOfTwo_CP_0_symbol: Boolean;
  -- links between control-path and data-path
  signal UGT_u32_u1_9_inst_req_0 : boolean;
  signal UGT_u32_u1_9_inst_ack_0 : boolean;
  signal MUX_16_inst_req_0 : boolean;
  signal MUX_16_inst_ack_0 : boolean;
  signal UGT_u32_u1_9_inst_req_1 : boolean;
  signal UGT_u32_u1_9_inst_ack_1 : boolean;
  signal MUX_16_inst_req_1 : boolean;
  signal MUX_16_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxOfTwo_input_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= a;
  a_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= b;
  b_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxOfTwo_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxOfTwo_out_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 32, 
      kill_counter_range => 1) -- 
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      kill => default_zero_sig,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxOfTwo_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxOfTwo_CP_0_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxOfTwo_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxOfTwo_CP_0: Block -- control-path 
    signal maxOfTwo_CP_0_elements: BooleanArray(13 downto 0);
    -- 
  begin -- 
    maxOfTwo_CP_0_elements(0) <= maxOfTwo_CP_0_start;
    maxOfTwo_CP_0_symbol <= maxOfTwo_CP_0_elements(13);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 1 
    -- members (4) 
      -- 	branch_block_stmt_5/$entry
      -- 	$entry
      -- 	branch_block_stmt_5/branch_block_stmt_5__entry__
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17__entry__
      -- 
    -- CP-element group 1 fork  transition  bypass 
    -- predecessors 0 
    -- successors 3 4 5 9 10 11 
    -- members (1) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/$entry
      -- 
    maxOfTwo_CP_0_elements(1) <= maxOfTwo_CP_0_elements(0);
    -- CP-element group 2 join  transition  output  bypass 
    -- predecessors 4 5 
    -- successors 6 
    -- members (3) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_sample_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Sample/$entry
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Sample/rr
      -- 
    cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 18) := "cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxOfTwo_CP_0_elements(4) & maxOfTwo_CP_0_elements(5);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxOfTwo_CP_0_elements(2), clk => clk, reset => reset); --
    end block;
    rr_30_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => maxOfTwo_CP_0_elements(2), ack => UGT_u32_u1_9_inst_req_0); -- 
    -- CP-element group 3 transition  output  bypass 
    -- predecessors 1 
    -- successors 7 
    -- members (3) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Update/$entry
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Update/cr
      -- 
    maxOfTwo_CP_0_elements(3) <= maxOfTwo_CP_0_elements(1);
    cr_35_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => maxOfTwo_CP_0_elements(3), ack => UGT_u32_u1_9_inst_req_1); -- 
    -- CP-element group 4 transition  bypass 
    -- predecessors 1 
    -- successors 2 
    -- members (4) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_7_sample_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_7_sample_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_7_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_7_update_completed_
      -- 
    maxOfTwo_CP_0_elements(4) <= maxOfTwo_CP_0_elements(1);
    -- CP-element group 5 transition  bypass 
    -- predecessors 1 
    -- successors 2 
    -- members (4) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_8_sample_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_8_sample_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_8_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_8_update_completed_
      -- 
    maxOfTwo_CP_0_elements(5) <= maxOfTwo_CP_0_elements(1);
    -- CP-element group 6 transition  input  bypass 
    -- predecessors 2 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_sample_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Sample/$exit
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Sample/ra
      -- 
    ra_31_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_9_inst_ack_0, ack => maxOfTwo_CP_0_elements(6)); -- 
    -- CP-element group 7 transition  input  bypass 
    -- predecessors 3 
    -- successors 8 
    -- members (7) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_update_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Update/$exit
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/UGT_u32_u1_9_Update/ca
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_iNsTr_0_13_sample_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_iNsTr_0_13_sample_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_iNsTr_0_13_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_iNsTr_0_13_update_completed_
      -- 
    ca_36_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_9_inst_ack_1, ack => maxOfTwo_CP_0_elements(7)); -- 
    -- CP-element group 8 join  transition  output  bypass 
    -- predecessors 7 10 11 
    -- successors 12 
    -- members (3) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_start/$entry
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_start/req
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_sample_start_
      -- 
    cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 18) := "cp_element_group_8"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxOfTwo_CP_0_elements(7) & maxOfTwo_CP_0_elements(10) & maxOfTwo_CP_0_elements(11);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxOfTwo_CP_0_elements(8), clk => clk, reset => reset); --
    end block;
    req_56_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => maxOfTwo_CP_0_elements(8), ack => MUX_16_inst_req_0); -- 
    -- CP-element group 9 transition  output  bypass 
    -- predecessors 1 
    -- successors 13 
    -- members (3) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_complete/$entry
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_complete/req
      -- 
    maxOfTwo_CP_0_elements(9) <= maxOfTwo_CP_0_elements(1);
    req_61_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => maxOfTwo_CP_0_elements(9), ack => MUX_16_inst_req_1); -- 
    -- CP-element group 10 transition  bypass 
    -- predecessors 1 
    -- successors 8 
    -- members (4) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_14_sample_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_14_sample_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_14_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_a_14_update_completed_
      -- 
    maxOfTwo_CP_0_elements(10) <= maxOfTwo_CP_0_elements(1);
    -- CP-element group 11 transition  bypass 
    -- predecessors 1 
    -- successors 8 
    -- members (4) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_15_sample_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_15_sample_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_15_update_start_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/R_b_15_update_completed_
      -- 
    maxOfTwo_CP_0_elements(11) <= maxOfTwo_CP_0_elements(1);
    -- CP-element group 12 transition  input  bypass 
    -- predecessors 8 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_start/$exit
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_start/ack
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_sample_completed_
      -- 
    ack_57_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_16_inst_ack_0, ack => maxOfTwo_CP_0_elements(12)); -- 
    -- CP-element group 13 transition  place  input  bypass 
    -- predecessors 9 
    -- successors 
    -- members (16) 
      -- 	branch_block_stmt_5/$exit
      -- 	$exit
      -- 	branch_block_stmt_5/merge_stmt_19__exit__
      -- 	branch_block_stmt_5/branch_block_stmt_5__exit__
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17__exit__
      -- 	branch_block_stmt_5/return__
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/$exit
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_update_completed_
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_complete/$exit
      -- 	branch_block_stmt_5/assign_stmt_11_to_assign_stmt_17/MUX_16_complete/ack
      -- 	branch_block_stmt_5/return___PhiReq/$entry
      -- 	branch_block_stmt_5/return___PhiReq/$exit
      -- 	branch_block_stmt_5/merge_stmt_19_PhiReqMerge
      -- 	branch_block_stmt_5/merge_stmt_19_PhiAck/$entry
      -- 	branch_block_stmt_5/merge_stmt_19_PhiAck/$exit
      -- 	branch_block_stmt_5/merge_stmt_19_PhiAck/dummy
      -- 
    ack_62_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_16_inst_ack_1, ack => maxOfTwo_CP_0_elements(13)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal iNsTr_0_11 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    MUX_16_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_16_inst_req_0;
      MUX_16_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_16_inst_req_1;
      MUX_16_inst_ack_1<= update_ack(0);
      MUX_16_inst: SelectSplitProtocol generic map(name => "MUX_16_inst", data_width => 32, buffering => 1, flow_through => false) -- 
        port map( x => a_buffer, y => b_buffer, sel => iNsTr_0_11, z => ret_val_x_x_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared split operator group (0) : UGT_u32_u1_9_inst 
    ApIntUgt_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= a_buffer & b_buffer;
      iNsTr_0_11 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_9_inst_req_0;
      UGT_u32_u1_9_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_9_inst_req_1;
      UGT_u32_u1_9_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    maxOfTwo_a : in  std_logic_vector(31 downto 0);
    maxOfTwo_b : in  std_logic_vector(31 downto 0);
    maxOfTwo_ret_val_x_x : out  std_logic_vector(31 downto 0);
    maxOfTwo_tag_in: in std_logic_vector(1 downto 0);
    maxOfTwo_tag_out: out std_logic_vector(1 downto 0);
    maxOfTwo_start_req : in std_logic;
    maxOfTwo_start_ack : out std_logic;
    maxOfTwo_fin_req   : in std_logic;
    maxOfTwo_fin_ack   : out std_logic;
    clk : in std_logic;
    reset : in std_logic); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- declarations related to module maxOfTwo
  component maxOfTwo is -- 
    generic (tag_length : integer); 
    port ( -- 
      a : in  std_logic_vector(31 downto 0);
      b : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- 
begin -- 
  -- module maxOfTwo
  maxOfTwo_instance:maxOfTwo-- 
    generic map(tag_length => 2)
    port map(-- 
      a => maxOfTwo_a,
      b => maxOfTwo_b,
      ret_val_x_x => maxOfTwo_ret_val_x_x,
      start_req => maxOfTwo_start_req,
      start_ack => maxOfTwo_start_ack,
      fin_req => maxOfTwo_fin_req,
      fin_ack => maxOfTwo_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => maxOfTwo_tag_in,
      tag_out => maxOfTwo_tag_out-- 
    ); -- 
  -- 
end Default;
