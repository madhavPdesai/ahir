-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant free_list_base_address : std_logic_vector(5 downto 0) := "000000";
  constant head_base_address : std_logic_vector(0 downto 0) := "0";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  constant xx_xstr1_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr2_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr3_base_address : std_logic_vector(2 downto 0) := "000";
  constant xx_xstr4_base_address : std_logic_vector(2 downto 0) := "000";
  constant xx_xstr5_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr6_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr_base_address : std_logic_vector(4 downto 0) := "00000";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity foo is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(15 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(15 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(95 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(47 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(15 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(127 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(47 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(47 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(23 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(7 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(23 downto 0);
    foo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    foo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    foo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    foo_out_pipe_write_req : out  std_logic_vector(0 downto 0);
    foo_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
    foo_out_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity foo;
architecture Default of foo is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_84_load_0_req_0 : boolean;
  signal ptr_deref_84_load_0_ack_0 : boolean;
  signal ptr_deref_84_load_1_req_0 : boolean;
  signal ptr_deref_84_load_1_ack_0 : boolean;
  signal simple_obj_ref_71_inst_req_0 : boolean;
  signal simple_obj_ref_71_inst_ack_0 : boolean;
  signal type_cast_72_inst_req_0 : boolean;
  signal type_cast_72_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal ptr_deref_79_gather_scatter_req_0 : boolean;
  signal ptr_deref_79_gather_scatter_ack_0 : boolean;
  signal ptr_deref_79_store_0_req_0 : boolean;
  signal ptr_deref_79_store_0_ack_0 : boolean;
  signal ptr_deref_79_store_1_req_0 : boolean;
  signal ptr_deref_79_store_1_ack_0 : boolean;
  signal ptr_deref_79_store_2_req_0 : boolean;
  signal ptr_deref_79_store_2_ack_0 : boolean;
  signal ptr_deref_79_store_3_req_0 : boolean;
  signal ptr_deref_79_store_3_ack_0 : boolean;
  signal ptr_deref_79_store_0_req_1 : boolean;
  signal ptr_deref_79_store_0_ack_1 : boolean;
  signal ptr_deref_79_store_1_req_1 : boolean;
  signal ptr_deref_79_store_1_ack_1 : boolean;
  signal ptr_deref_79_store_2_req_1 : boolean;
  signal ptr_deref_79_store_2_ack_1 : boolean;
  signal ptr_deref_79_store_3_req_1 : boolean;
  signal ptr_deref_79_store_3_ack_1 : boolean;
  signal array_obj_ref_107_root_address_inst_req_0 : boolean;
  signal array_obj_ref_107_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_107_root_address_inst_req_1 : boolean;
  signal array_obj_ref_107_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_107_final_reg_req_0 : boolean;
  signal array_obj_ref_107_final_reg_ack_0 : boolean;
  signal ptr_deref_84_load_2_req_0 : boolean;
  signal ptr_deref_84_load_2_ack_0 : boolean;
  signal ptr_deref_84_load_3_req_0 : boolean;
  signal ptr_deref_84_load_3_ack_0 : boolean;
  signal ptr_deref_84_load_0_req_1 : boolean;
  signal ptr_deref_84_load_0_ack_1 : boolean;
  signal ptr_deref_84_load_1_req_1 : boolean;
  signal ptr_deref_84_load_1_ack_1 : boolean;
  signal ptr_deref_84_load_2_req_1 : boolean;
  signal ptr_deref_84_load_2_ack_1 : boolean;
  signal ptr_deref_84_load_3_req_1 : boolean;
  signal ptr_deref_84_load_3_ack_1 : boolean;
  signal ptr_deref_84_gather_scatter_req_0 : boolean;
  signal ptr_deref_84_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_89_base_resize_req_0 : boolean;
  signal array_obj_ref_89_base_resize_ack_0 : boolean;
  signal array_obj_ref_89_root_address_inst_req_0 : boolean;
  signal array_obj_ref_89_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_89_root_address_inst_req_1 : boolean;
  signal array_obj_ref_89_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_89_final_reg_req_0 : boolean;
  signal array_obj_ref_89_final_reg_ack_0 : boolean;
  signal ptr_deref_93_base_resize_req_0 : boolean;
  signal ptr_deref_93_base_resize_ack_0 : boolean;
  signal ptr_deref_93_root_address_inst_req_0 : boolean;
  signal ptr_deref_93_root_address_inst_ack_0 : boolean;
  signal ptr_deref_93_addr_0_req_0 : boolean;
  signal ptr_deref_93_addr_0_ack_0 : boolean;
  signal ptr_deref_93_addr_0_req_1 : boolean;
  signal ptr_deref_93_addr_0_ack_1 : boolean;
  signal ptr_deref_93_addr_1_req_0 : boolean;
  signal ptr_deref_93_addr_1_ack_0 : boolean;
  signal ptr_deref_93_addr_1_req_1 : boolean;
  signal ptr_deref_93_addr_1_ack_1 : boolean;
  signal ptr_deref_93_addr_2_req_0 : boolean;
  signal ptr_deref_93_addr_2_ack_0 : boolean;
  signal ptr_deref_93_addr_2_req_1 : boolean;
  signal ptr_deref_93_addr_2_ack_1 : boolean;
  signal ptr_deref_93_addr_3_req_0 : boolean;
  signal ptr_deref_93_addr_3_ack_0 : boolean;
  signal ptr_deref_93_addr_3_req_1 : boolean;
  signal ptr_deref_93_addr_3_ack_1 : boolean;
  signal ptr_deref_93_load_0_req_0 : boolean;
  signal ptr_deref_93_load_0_ack_0 : boolean;
  signal ptr_deref_93_load_1_req_0 : boolean;
  signal ptr_deref_93_load_1_ack_0 : boolean;
  signal ptr_deref_93_load_2_req_0 : boolean;
  signal ptr_deref_93_load_2_ack_0 : boolean;
  signal ptr_deref_93_load_3_req_0 : boolean;
  signal ptr_deref_93_load_3_ack_0 : boolean;
  signal ptr_deref_93_load_0_req_1 : boolean;
  signal ptr_deref_93_load_0_ack_1 : boolean;
  signal ptr_deref_93_load_1_req_1 : boolean;
  signal ptr_deref_93_load_1_ack_1 : boolean;
  signal ptr_deref_93_load_2_req_1 : boolean;
  signal ptr_deref_93_load_2_ack_1 : boolean;
  signal ptr_deref_93_load_3_req_1 : boolean;
  signal ptr_deref_93_load_3_ack_1 : boolean;
  signal ptr_deref_93_gather_scatter_req_0 : boolean;
  signal ptr_deref_93_gather_scatter_ack_0 : boolean;
  signal binary_98_inst_req_0 : boolean;
  signal binary_98_inst_ack_0 : boolean;
  signal binary_98_inst_req_1 : boolean;
  signal binary_98_inst_ack_1 : boolean;
  signal ptr_deref_102_load_0_req_0 : boolean;
  signal ptr_deref_102_load_0_ack_0 : boolean;
  signal ptr_deref_102_load_1_req_0 : boolean;
  signal ptr_deref_102_load_1_ack_0 : boolean;
  signal ptr_deref_102_load_2_req_0 : boolean;
  signal ptr_deref_102_load_2_ack_0 : boolean;
  signal ptr_deref_102_load_3_req_0 : boolean;
  signal ptr_deref_102_load_3_ack_0 : boolean;
  signal ptr_deref_102_load_0_req_1 : boolean;
  signal ptr_deref_102_load_0_ack_1 : boolean;
  signal ptr_deref_102_load_1_req_1 : boolean;
  signal ptr_deref_102_load_1_ack_1 : boolean;
  signal ptr_deref_102_load_2_req_1 : boolean;
  signal ptr_deref_102_load_2_ack_1 : boolean;
  signal ptr_deref_102_load_3_req_1 : boolean;
  signal ptr_deref_102_load_3_ack_1 : boolean;
  signal ptr_deref_102_gather_scatter_req_0 : boolean;
  signal ptr_deref_102_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_107_base_resize_req_0 : boolean;
  signal array_obj_ref_107_base_resize_ack_0 : boolean;
  signal ptr_deref_110_base_resize_req_0 : boolean;
  signal ptr_deref_110_base_resize_ack_0 : boolean;
  signal ptr_deref_110_root_address_inst_req_0 : boolean;
  signal ptr_deref_110_root_address_inst_ack_0 : boolean;
  signal ptr_deref_110_addr_0_req_0 : boolean;
  signal ptr_deref_110_addr_0_ack_0 : boolean;
  signal ptr_deref_110_addr_0_req_1 : boolean;
  signal ptr_deref_110_addr_0_ack_1 : boolean;
  signal ptr_deref_110_addr_1_req_0 : boolean;
  signal ptr_deref_110_addr_1_ack_0 : boolean;
  signal ptr_deref_110_addr_1_req_1 : boolean;
  signal ptr_deref_110_addr_1_ack_1 : boolean;
  signal ptr_deref_110_addr_2_req_0 : boolean;
  signal ptr_deref_110_addr_2_ack_0 : boolean;
  signal ptr_deref_110_addr_2_req_1 : boolean;
  signal ptr_deref_110_addr_2_ack_1 : boolean;
  signal ptr_deref_110_addr_3_req_0 : boolean;
  signal ptr_deref_110_addr_3_ack_0 : boolean;
  signal ptr_deref_110_addr_3_req_1 : boolean;
  signal ptr_deref_110_addr_3_ack_1 : boolean;
  signal ptr_deref_110_gather_scatter_req_0 : boolean;
  signal ptr_deref_110_gather_scatter_ack_0 : boolean;
  signal ptr_deref_110_store_0_req_0 : boolean;
  signal ptr_deref_110_store_0_ack_0 : boolean;
  signal ptr_deref_110_store_1_req_0 : boolean;
  signal ptr_deref_110_store_1_ack_0 : boolean;
  signal ptr_deref_110_store_2_req_0 : boolean;
  signal ptr_deref_110_store_2_ack_0 : boolean;
  signal ptr_deref_110_store_3_req_0 : boolean;
  signal ptr_deref_110_store_3_ack_0 : boolean;
  signal ptr_deref_110_store_0_req_1 : boolean;
  signal ptr_deref_110_store_0_ack_1 : boolean;
  signal ptr_deref_110_store_1_req_1 : boolean;
  signal ptr_deref_110_store_1_ack_1 : boolean;
  signal ptr_deref_110_store_2_req_1 : boolean;
  signal ptr_deref_110_store_2_ack_1 : boolean;
  signal ptr_deref_110_store_3_req_1 : boolean;
  signal ptr_deref_110_store_3_ack_1 : boolean;
  signal ptr_deref_115_load_0_req_0 : boolean;
  signal ptr_deref_115_load_0_ack_0 : boolean;
  signal ptr_deref_115_load_1_req_0 : boolean;
  signal ptr_deref_115_load_1_ack_0 : boolean;
  signal ptr_deref_115_load_2_req_0 : boolean;
  signal ptr_deref_115_load_2_ack_0 : boolean;
  signal ptr_deref_115_load_3_req_0 : boolean;
  signal ptr_deref_115_load_3_ack_0 : boolean;
  signal ptr_deref_115_load_0_req_1 : boolean;
  signal ptr_deref_115_load_0_ack_1 : boolean;
  signal ptr_deref_115_load_1_req_1 : boolean;
  signal ptr_deref_115_load_1_ack_1 : boolean;
  signal ptr_deref_115_load_2_req_1 : boolean;
  signal ptr_deref_115_load_2_ack_1 : boolean;
  signal ptr_deref_115_load_3_req_1 : boolean;
  signal ptr_deref_115_load_3_ack_1 : boolean;
  signal ptr_deref_115_gather_scatter_req_0 : boolean;
  signal ptr_deref_115_gather_scatter_ack_0 : boolean;
  signal type_cast_119_inst_req_0 : boolean;
  signal type_cast_119_inst_ack_0 : boolean;
  signal type_cast_128_inst_req_0 : boolean;
  signal type_cast_128_inst_ack_0 : boolean;
  signal simple_obj_ref_126_inst_req_0 : boolean;
  signal simple_obj_ref_126_inst_ack_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  foo_CP_0: Block -- control-path 
    signal foo_CP_0_start: Boolean;
    signal Xentry_1_symbol: Boolean;
    signal Xexit_2_symbol: Boolean;
    signal branch_block_stmt_56_3_symbol : Boolean;
    -- 
  begin -- 
    foo_CP_0_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_1_symbol  <= foo_CP_0_start; -- transition $entry
    branch_block_stmt_56_3: Block -- branch_block_stmt_56 
      signal branch_block_stmt_56_3_start: Boolean;
      signal Xentry_4_symbol: Boolean;
      signal Xexit_5_symbol: Boolean;
      signal branch_block_stmt_56_x_xentry_x_xx_x6_symbol : Boolean;
      signal branch_block_stmt_56_x_xexit_x_xx_x7_symbol : Boolean;
      signal assign_stmt_61_x_xentry_x_xx_x8_symbol : Boolean;
      signal assign_stmt_61_x_xexit_x_xx_x9_symbol : Boolean;
      signal bb_0_bb_1_10_symbol : Boolean;
      signal merge_stmt_63_x_xexit_x_xx_x11_symbol : Boolean;
      signal assign_stmt_68_x_xentry_x_xx_x12_symbol : Boolean;
      signal assign_stmt_68_x_xexit_x_xx_x13_symbol : Boolean;
      signal assign_stmt_73_x_xentry_x_xx_x14_symbol : Boolean;
      signal assign_stmt_73_x_xexit_x_xx_x15_symbol : Boolean;
      signal assign_stmt_77_to_assign_stmt_125_x_xentry_x_xx_x16_symbol : Boolean;
      signal assign_stmt_77_to_assign_stmt_125_x_xexit_x_xx_x17_symbol : Boolean;
      signal assign_stmt_129_x_xentry_x_xx_x18_symbol : Boolean;
      signal assign_stmt_129_x_xexit_x_xx_x19_symbol : Boolean;
      signal bb_1_bb_1_20_symbol : Boolean;
      signal assign_stmt_61_21_symbol : Boolean;
      signal assign_stmt_68_24_symbol : Boolean;
      signal assign_stmt_73_27_symbol : Boolean;
      signal assign_stmt_77_to_assign_stmt_125_45_symbol : Boolean;
      signal assign_stmt_129_584_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_603_symbol : Boolean;
      signal bb_1_bb_1_PhiReq_606_symbol : Boolean;
      signal merge_stmt_63_PhiReqMerge_609_symbol : Boolean;
      signal merge_stmt_63_PhiAck_610_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_56_3_start <= Xentry_1_symbol; -- control passed to block
      Xentry_4_symbol  <= branch_block_stmt_56_3_start; -- transition branch_block_stmt_56/$entry
      branch_block_stmt_56_x_xentry_x_xx_x6_symbol  <=  Xentry_4_symbol; -- place branch_block_stmt_56/branch_block_stmt_56__entry__ (optimized away) 
      branch_block_stmt_56_x_xexit_x_xx_x7_symbol  <=   false ; -- place branch_block_stmt_56/branch_block_stmt_56__exit__ (optimized away) 
      assign_stmt_61_x_xentry_x_xx_x8_symbol  <=  branch_block_stmt_56_x_xentry_x_xx_x6_symbol; -- place branch_block_stmt_56/assign_stmt_61__entry__ (optimized away) 
      assign_stmt_61_x_xexit_x_xx_x9_symbol  <=  assign_stmt_61_21_symbol; -- place branch_block_stmt_56/assign_stmt_61__exit__ (optimized away) 
      bb_0_bb_1_10_symbol  <=  assign_stmt_61_x_xexit_x_xx_x9_symbol; -- place branch_block_stmt_56/bb_0_bb_1 (optimized away) 
      merge_stmt_63_x_xexit_x_xx_x11_symbol  <=  merge_stmt_63_PhiAck_610_symbol; -- place branch_block_stmt_56/merge_stmt_63__exit__ (optimized away) 
      assign_stmt_68_x_xentry_x_xx_x12_symbol  <=  merge_stmt_63_x_xexit_x_xx_x11_symbol; -- place branch_block_stmt_56/assign_stmt_68__entry__ (optimized away) 
      assign_stmt_68_x_xexit_x_xx_x13_symbol  <=  assign_stmt_68_24_symbol; -- place branch_block_stmt_56/assign_stmt_68__exit__ (optimized away) 
      assign_stmt_73_x_xentry_x_xx_x14_symbol  <=  assign_stmt_68_x_xexit_x_xx_x13_symbol; -- place branch_block_stmt_56/assign_stmt_73__entry__ (optimized away) 
      assign_stmt_73_x_xexit_x_xx_x15_symbol  <=  assign_stmt_73_27_symbol; -- place branch_block_stmt_56/assign_stmt_73__exit__ (optimized away) 
      assign_stmt_77_to_assign_stmt_125_x_xentry_x_xx_x16_symbol  <=  assign_stmt_73_x_xexit_x_xx_x15_symbol; -- place branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125__entry__ (optimized away) 
      assign_stmt_77_to_assign_stmt_125_x_xexit_x_xx_x17_symbol  <=  assign_stmt_77_to_assign_stmt_125_45_symbol; -- place branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125__exit__ (optimized away) 
      assign_stmt_129_x_xentry_x_xx_x18_symbol  <=  assign_stmt_77_to_assign_stmt_125_x_xexit_x_xx_x17_symbol; -- place branch_block_stmt_56/assign_stmt_129__entry__ (optimized away) 
      assign_stmt_129_x_xexit_x_xx_x19_symbol  <=  assign_stmt_129_584_symbol; -- place branch_block_stmt_56/assign_stmt_129__exit__ (optimized away) 
      bb_1_bb_1_20_symbol  <=  assign_stmt_129_x_xexit_x_xx_x19_symbol; -- place branch_block_stmt_56/bb_1_bb_1 (optimized away) 
      assign_stmt_61_21: Block -- branch_block_stmt_56/assign_stmt_61 
        signal assign_stmt_61_21_start: Boolean;
        signal Xentry_22_symbol: Boolean;
        signal Xexit_23_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_61_21_start <= assign_stmt_61_x_xentry_x_xx_x8_symbol; -- control passed to block
        Xentry_22_symbol  <= assign_stmt_61_21_start; -- transition branch_block_stmt_56/assign_stmt_61/$entry
        Xexit_23_symbol <= Xentry_22_symbol; -- transition branch_block_stmt_56/assign_stmt_61/$exit
        assign_stmt_61_21_symbol <= Xexit_23_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_61
      assign_stmt_68_24: Block -- branch_block_stmt_56/assign_stmt_68 
        signal assign_stmt_68_24_start: Boolean;
        signal Xentry_25_symbol: Boolean;
        signal Xexit_26_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_68_24_start <= assign_stmt_68_x_xentry_x_xx_x12_symbol; -- control passed to block
        Xentry_25_symbol  <= assign_stmt_68_24_start; -- transition branch_block_stmt_56/assign_stmt_68/$entry
        Xexit_26_symbol <= Xentry_25_symbol; -- transition branch_block_stmt_56/assign_stmt_68/$exit
        assign_stmt_68_24_symbol <= Xexit_26_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_68
      assign_stmt_73_27: Block -- branch_block_stmt_56/assign_stmt_73 
        signal assign_stmt_73_27_start: Boolean;
        signal Xentry_28_symbol: Boolean;
        signal Xexit_29_symbol: Boolean;
        signal assign_stmt_73_active_x_x30_symbol : Boolean;
        signal assign_stmt_73_completed_x_x31_symbol : Boolean;
        signal type_cast_72_active_x_x32_symbol : Boolean;
        signal type_cast_72_trigger_x_x33_symbol : Boolean;
        signal simple_obj_ref_71_trigger_x_x34_symbol : Boolean;
        signal simple_obj_ref_71_complete_35_symbol : Boolean;
        signal type_cast_72_complete_40_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_73_27_start <= assign_stmt_73_x_xentry_x_xx_x14_symbol; -- control passed to block
        Xentry_28_symbol  <= assign_stmt_73_27_start; -- transition branch_block_stmt_56/assign_stmt_73/$entry
        assign_stmt_73_active_x_x30_symbol <= type_cast_72_complete_40_symbol; -- transition branch_block_stmt_56/assign_stmt_73/assign_stmt_73_active_
        assign_stmt_73_completed_x_x31_symbol <= assign_stmt_73_active_x_x30_symbol; -- transition branch_block_stmt_56/assign_stmt_73/assign_stmt_73_completed_
        type_cast_72_active_x_x32_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_73/type_cast_72_active_ 
          signal type_cast_72_active_x_x32_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_72_active_x_x32_predecessors(0) <= type_cast_72_trigger_x_x33_symbol;
          type_cast_72_active_x_x32_predecessors(1) <= simple_obj_ref_71_complete_35_symbol;
          type_cast_72_active_x_x32_join: join -- 
            port map( -- 
              preds => type_cast_72_active_x_x32_predecessors,
              symbol_out => type_cast_72_active_x_x32_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_73/type_cast_72_active_
        type_cast_72_trigger_x_x33_symbol <= Xentry_28_symbol; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_trigger_
        simple_obj_ref_71_trigger_x_x34_symbol <= Xentry_28_symbol; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_trigger_
        simple_obj_ref_71_complete_35: Block -- branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete 
          signal simple_obj_ref_71_complete_35_start: Boolean;
          signal Xentry_36_symbol: Boolean;
          signal Xexit_37_symbol: Boolean;
          signal req_38_symbol : Boolean;
          signal ack_39_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_71_complete_35_start <= simple_obj_ref_71_trigger_x_x34_symbol; -- control passed to block
          Xentry_36_symbol  <= simple_obj_ref_71_complete_35_start; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/$entry
          req_38_symbol <= Xentry_36_symbol; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/req
          simple_obj_ref_71_inst_req_0 <= req_38_symbol; -- link to DP
          ack_39_symbol <= simple_obj_ref_71_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/ack
          Xexit_37_symbol <= ack_39_symbol; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/$exit
          simple_obj_ref_71_complete_35_symbol <= Xexit_37_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete
        type_cast_72_complete_40: Block -- branch_block_stmt_56/assign_stmt_73/type_cast_72_complete 
          signal type_cast_72_complete_40_start: Boolean;
          signal Xentry_41_symbol: Boolean;
          signal Xexit_42_symbol: Boolean;
          signal req_43_symbol : Boolean;
          signal ack_44_symbol : Boolean;
          -- 
        begin -- 
          type_cast_72_complete_40_start <= type_cast_72_active_x_x32_symbol; -- control passed to block
          Xentry_41_symbol  <= type_cast_72_complete_40_start; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/$entry
          req_43_symbol <= Xentry_41_symbol; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/req
          type_cast_72_inst_req_0 <= req_43_symbol; -- link to DP
          ack_44_symbol <= type_cast_72_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/ack
          Xexit_42_symbol <= ack_44_symbol; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/$exit
          type_cast_72_complete_40_symbol <= Xexit_42_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_73/type_cast_72_complete
        Xexit_29_symbol <= assign_stmt_73_completed_x_x31_symbol; -- transition branch_block_stmt_56/assign_stmt_73/$exit
        assign_stmt_73_27_symbol <= Xexit_29_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_73
      assign_stmt_77_to_assign_stmt_125_45: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125 
        signal assign_stmt_77_to_assign_stmt_125_45_start: Boolean;
        signal Xentry_46_symbol: Boolean;
        signal Xexit_47_symbol: Boolean;
        signal assign_stmt_77_active_x_x48_symbol : Boolean;
        signal assign_stmt_77_completed_x_x49_symbol : Boolean;
        signal type_cast_76_active_x_x50_symbol : Boolean;
        signal type_cast_76_trigger_x_x51_symbol : Boolean;
        signal simple_obj_ref_75_complete_52_symbol : Boolean;
        signal type_cast_76_complete_53_symbol : Boolean;
        signal assign_stmt_81_active_x_x58_symbol : Boolean;
        signal assign_stmt_81_completed_x_x59_symbol : Boolean;
        signal simple_obj_ref_80_complete_60_symbol : Boolean;
        signal ptr_deref_79_trigger_x_x61_symbol : Boolean;
        signal ptr_deref_79_active_x_x62_symbol : Boolean;
        signal ptr_deref_79_base_address_calculated_63_symbol : Boolean;
        signal ptr_deref_79_root_address_calculated_64_symbol : Boolean;
        signal ptr_deref_79_word_address_calculated_65_symbol : Boolean;
        signal ptr_deref_79_request_66_symbol : Boolean;
        signal ptr_deref_79_complete_94_symbol : Boolean;
        signal assign_stmt_85_active_x_x120_symbol : Boolean;
        signal assign_stmt_85_completed_x_x121_symbol : Boolean;
        signal ptr_deref_84_trigger_x_x122_symbol : Boolean;
        signal ptr_deref_84_active_x_x123_symbol : Boolean;
        signal ptr_deref_84_base_address_calculated_124_symbol : Boolean;
        signal ptr_deref_84_root_address_calculated_125_symbol : Boolean;
        signal ptr_deref_84_word_address_calculated_126_symbol : Boolean;
        signal ptr_deref_84_request_127_symbol : Boolean;
        signal ptr_deref_84_complete_153_symbol : Boolean;
        signal assign_stmt_90_active_x_x181_symbol : Boolean;
        signal assign_stmt_90_completed_x_x182_symbol : Boolean;
        signal array_obj_ref_89_trigger_x_x183_symbol : Boolean;
        signal array_obj_ref_89_active_x_x184_symbol : Boolean;
        signal array_obj_ref_89_base_address_calculated_185_symbol : Boolean;
        signal array_obj_ref_89_root_address_calculated_186_symbol : Boolean;
        signal array_obj_ref_89_base_address_resized_187_symbol : Boolean;
        signal array_obj_ref_89_base_addr_resize_188_symbol : Boolean;
        signal array_obj_ref_89_base_plus_offset_trigger_193_symbol : Boolean;
        signal array_obj_ref_89_base_plus_offset_194_symbol : Boolean;
        signal array_obj_ref_89_complete_201_symbol : Boolean;
        signal assign_stmt_94_active_x_x206_symbol : Boolean;
        signal assign_stmt_94_completed_x_x207_symbol : Boolean;
        signal ptr_deref_93_trigger_x_x208_symbol : Boolean;
        signal ptr_deref_93_active_x_x209_symbol : Boolean;
        signal ptr_deref_93_base_address_calculated_210_symbol : Boolean;
        signal simple_obj_ref_92_complete_211_symbol : Boolean;
        signal ptr_deref_93_root_address_calculated_212_symbol : Boolean;
        signal ptr_deref_93_word_address_calculated_213_symbol : Boolean;
        signal ptr_deref_93_base_address_resized_214_symbol : Boolean;
        signal ptr_deref_93_base_addr_resize_215_symbol : Boolean;
        signal ptr_deref_93_base_plus_offset_220_symbol : Boolean;
        signal ptr_deref_93_word_addrgen_225_symbol : Boolean;
        signal ptr_deref_93_request_256_symbol : Boolean;
        signal ptr_deref_93_complete_282_symbol : Boolean;
        signal assign_stmt_99_active_x_x310_symbol : Boolean;
        signal assign_stmt_99_completed_x_x311_symbol : Boolean;
        signal binary_98_active_x_x312_symbol : Boolean;
        signal binary_98_trigger_x_x313_symbol : Boolean;
        signal simple_obj_ref_97_complete_314_symbol : Boolean;
        signal binary_98_complete_315_symbol : Boolean;
        signal assign_stmt_103_active_x_x322_symbol : Boolean;
        signal assign_stmt_103_completed_x_x323_symbol : Boolean;
        signal ptr_deref_102_trigger_x_x324_symbol : Boolean;
        signal ptr_deref_102_active_x_x325_symbol : Boolean;
        signal ptr_deref_102_base_address_calculated_326_symbol : Boolean;
        signal ptr_deref_102_root_address_calculated_327_symbol : Boolean;
        signal ptr_deref_102_word_address_calculated_328_symbol : Boolean;
        signal ptr_deref_102_request_329_symbol : Boolean;
        signal ptr_deref_102_complete_355_symbol : Boolean;
        signal assign_stmt_108_active_x_x383_symbol : Boolean;
        signal assign_stmt_108_completed_x_x384_symbol : Boolean;
        signal array_obj_ref_107_trigger_x_x385_symbol : Boolean;
        signal array_obj_ref_107_active_x_x386_symbol : Boolean;
        signal array_obj_ref_107_base_address_calculated_387_symbol : Boolean;
        signal array_obj_ref_107_root_address_calculated_388_symbol : Boolean;
        signal array_obj_ref_107_base_address_resized_389_symbol : Boolean;
        signal array_obj_ref_107_base_addr_resize_390_symbol : Boolean;
        signal array_obj_ref_107_base_plus_offset_trigger_395_symbol : Boolean;
        signal array_obj_ref_107_base_plus_offset_396_symbol : Boolean;
        signal array_obj_ref_107_complete_403_symbol : Boolean;
        signal assign_stmt_112_active_x_x408_symbol : Boolean;
        signal assign_stmt_112_completed_x_x409_symbol : Boolean;
        signal simple_obj_ref_111_complete_410_symbol : Boolean;
        signal ptr_deref_110_trigger_x_x411_symbol : Boolean;
        signal ptr_deref_110_active_x_x412_symbol : Boolean;
        signal ptr_deref_110_base_address_calculated_413_symbol : Boolean;
        signal simple_obj_ref_109_complete_414_symbol : Boolean;
        signal ptr_deref_110_root_address_calculated_415_symbol : Boolean;
        signal ptr_deref_110_word_address_calculated_416_symbol : Boolean;
        signal ptr_deref_110_base_address_resized_417_symbol : Boolean;
        signal ptr_deref_110_base_addr_resize_418_symbol : Boolean;
        signal ptr_deref_110_base_plus_offset_423_symbol : Boolean;
        signal ptr_deref_110_word_addrgen_428_symbol : Boolean;
        signal ptr_deref_110_request_459_symbol : Boolean;
        signal ptr_deref_110_complete_487_symbol : Boolean;
        signal assign_stmt_116_active_x_x513_symbol : Boolean;
        signal assign_stmt_116_completed_x_x514_symbol : Boolean;
        signal ptr_deref_115_trigger_x_x515_symbol : Boolean;
        signal ptr_deref_115_active_x_x516_symbol : Boolean;
        signal ptr_deref_115_base_address_calculated_517_symbol : Boolean;
        signal ptr_deref_115_root_address_calculated_518_symbol : Boolean;
        signal ptr_deref_115_word_address_calculated_519_symbol : Boolean;
        signal ptr_deref_115_request_520_symbol : Boolean;
        signal ptr_deref_115_complete_546_symbol : Boolean;
        signal assign_stmt_120_active_x_x574_symbol : Boolean;
        signal assign_stmt_120_completed_x_x575_symbol : Boolean;
        signal type_cast_119_active_x_x576_symbol : Boolean;
        signal type_cast_119_trigger_x_x577_symbol : Boolean;
        signal simple_obj_ref_118_complete_578_symbol : Boolean;
        signal type_cast_119_complete_579_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_77_to_assign_stmt_125_45_start <= assign_stmt_77_to_assign_stmt_125_x_xentry_x_xx_x16_symbol; -- control passed to block
        Xentry_46_symbol  <= assign_stmt_77_to_assign_stmt_125_45_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/$entry
        assign_stmt_77_active_x_x48_symbol <= type_cast_76_complete_53_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_77_active_
        assign_stmt_77_completed_x_x49_symbol <= assign_stmt_77_active_x_x48_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_77_completed_
        type_cast_76_active_x_x50_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_active_ 
          signal type_cast_76_active_x_x50_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_76_active_x_x50_predecessors(0) <= type_cast_76_trigger_x_x51_symbol;
          type_cast_76_active_x_x50_predecessors(1) <= simple_obj_ref_75_complete_52_symbol;
          type_cast_76_active_x_x50_join: join -- 
            port map( -- 
              preds => type_cast_76_active_x_x50_predecessors,
              symbol_out => type_cast_76_active_x_x50_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_active_
        type_cast_76_trigger_x_x51_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_trigger_
        simple_obj_ref_75_complete_52_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_75_complete
        type_cast_76_complete_53: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete 
          signal type_cast_76_complete_53_start: Boolean;
          signal Xentry_54_symbol: Boolean;
          signal Xexit_55_symbol: Boolean;
          signal req_56_symbol : Boolean;
          signal ack_57_symbol : Boolean;
          -- 
        begin -- 
          type_cast_76_complete_53_start <= type_cast_76_active_x_x50_symbol; -- control passed to block
          Xentry_54_symbol  <= type_cast_76_complete_53_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/$entry
          req_56_symbol <= Xentry_54_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/req
          type_cast_76_inst_req_0 <= req_56_symbol; -- link to DP
          ack_57_symbol <= type_cast_76_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/ack
          Xexit_55_symbol <= ack_57_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/$exit
          type_cast_76_complete_53_symbol <= Xexit_55_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete
        assign_stmt_81_active_x_x58_symbol <= simple_obj_ref_80_complete_60_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_81_active_
        assign_stmt_81_completed_x_x59_symbol <= ptr_deref_79_complete_94_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_81_completed_
        simple_obj_ref_80_complete_60_symbol <= assign_stmt_77_completed_x_x49_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_80_complete
        ptr_deref_79_trigger_x_x61_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_trigger_ 
          signal ptr_deref_79_trigger_x_x61_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_79_trigger_x_x61_predecessors(0) <= ptr_deref_79_word_address_calculated_65_symbol;
          ptr_deref_79_trigger_x_x61_predecessors(1) <= assign_stmt_81_active_x_x58_symbol;
          ptr_deref_79_trigger_x_x61_join: join -- 
            port map( -- 
              preds => ptr_deref_79_trigger_x_x61_predecessors,
              symbol_out => ptr_deref_79_trigger_x_x61_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_trigger_
        ptr_deref_79_active_x_x62_symbol <= ptr_deref_79_request_66_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_active_
        ptr_deref_79_base_address_calculated_63_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_base_address_calculated
        ptr_deref_79_root_address_calculated_64_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_root_address_calculated
        ptr_deref_79_word_address_calculated_65_symbol <= ptr_deref_79_root_address_calculated_64_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_word_address_calculated
        ptr_deref_79_request_66: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request 
          signal ptr_deref_79_request_66_start: Boolean;
          signal Xentry_67_symbol: Boolean;
          signal Xexit_68_symbol: Boolean;
          signal split_req_69_symbol : Boolean;
          signal split_ack_70_symbol : Boolean;
          signal word_access_71_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_79_request_66_start <= ptr_deref_79_trigger_x_x61_symbol; -- control passed to block
          Xentry_67_symbol  <= ptr_deref_79_request_66_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/$entry
          split_req_69_symbol <= Xentry_67_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/split_req
          ptr_deref_79_gather_scatter_req_0 <= split_req_69_symbol; -- link to DP
          split_ack_70_symbol <= ptr_deref_79_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/split_ack
          word_access_71: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access 
            signal word_access_71_start: Boolean;
            signal Xentry_72_symbol: Boolean;
            signal Xexit_73_symbol: Boolean;
            signal word_access_0_74_symbol : Boolean;
            signal word_access_1_79_symbol : Boolean;
            signal word_access_2_84_symbol : Boolean;
            signal word_access_3_89_symbol : Boolean;
            -- 
          begin -- 
            word_access_71_start <= split_ack_70_symbol; -- control passed to block
            Xentry_72_symbol  <= word_access_71_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/$entry
            word_access_0_74: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0 
              signal word_access_0_74_start: Boolean;
              signal Xentry_75_symbol: Boolean;
              signal Xexit_76_symbol: Boolean;
              signal rr_77_symbol : Boolean;
              signal ra_78_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_74_start <= Xentry_72_symbol; -- control passed to block
              Xentry_75_symbol  <= word_access_0_74_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/$entry
              rr_77_symbol <= Xentry_75_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/rr
              ptr_deref_79_store_0_req_0 <= rr_77_symbol; -- link to DP
              ra_78_symbol <= ptr_deref_79_store_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/ra
              Xexit_76_symbol <= ra_78_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/$exit
              word_access_0_74_symbol <= Xexit_76_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0
            word_access_1_79: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_1 
              signal word_access_1_79_start: Boolean;
              signal Xentry_80_symbol: Boolean;
              signal Xexit_81_symbol: Boolean;
              signal rr_82_symbol : Boolean;
              signal ra_83_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_79_start <= Xentry_72_symbol; -- control passed to block
              Xentry_80_symbol  <= word_access_1_79_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_1/$entry
              rr_82_symbol <= Xentry_80_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_1/rr
              ptr_deref_79_store_1_req_0 <= rr_82_symbol; -- link to DP
              ra_83_symbol <= ptr_deref_79_store_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_1/ra
              Xexit_81_symbol <= ra_83_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_1/$exit
              word_access_1_79_symbol <= Xexit_81_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_1
            word_access_2_84: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_2 
              signal word_access_2_84_start: Boolean;
              signal Xentry_85_symbol: Boolean;
              signal Xexit_86_symbol: Boolean;
              signal rr_87_symbol : Boolean;
              signal ra_88_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_84_start <= Xentry_72_symbol; -- control passed to block
              Xentry_85_symbol  <= word_access_2_84_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_2/$entry
              rr_87_symbol <= Xentry_85_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_2/rr
              ptr_deref_79_store_2_req_0 <= rr_87_symbol; -- link to DP
              ra_88_symbol <= ptr_deref_79_store_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_2/ra
              Xexit_86_symbol <= ra_88_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_2/$exit
              word_access_2_84_symbol <= Xexit_86_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_2
            word_access_3_89: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_3 
              signal word_access_3_89_start: Boolean;
              signal Xentry_90_symbol: Boolean;
              signal Xexit_91_symbol: Boolean;
              signal rr_92_symbol : Boolean;
              signal ra_93_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_89_start <= Xentry_72_symbol; -- control passed to block
              Xentry_90_symbol  <= word_access_3_89_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_3/$entry
              rr_92_symbol <= Xentry_90_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_3/rr
              ptr_deref_79_store_3_req_0 <= rr_92_symbol; -- link to DP
              ra_93_symbol <= ptr_deref_79_store_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_3/ra
              Xexit_91_symbol <= ra_93_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_3/$exit
              word_access_3_89_symbol <= Xexit_91_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_3
            Xexit_73_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/$exit 
              signal Xexit_73_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_73_predecessors(0) <= word_access_0_74_symbol;
              Xexit_73_predecessors(1) <= word_access_1_79_symbol;
              Xexit_73_predecessors(2) <= word_access_2_84_symbol;
              Xexit_73_predecessors(3) <= word_access_3_89_symbol;
              Xexit_73_join: join -- 
                port map( -- 
                  preds => Xexit_73_predecessors,
                  symbol_out => Xexit_73_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/$exit
            word_access_71_symbol <= Xexit_73_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access
          Xexit_68_symbol <= word_access_71_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/$exit
          ptr_deref_79_request_66_symbol <= Xexit_68_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request
        ptr_deref_79_complete_94: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete 
          signal ptr_deref_79_complete_94_start: Boolean;
          signal Xentry_95_symbol: Boolean;
          signal Xexit_96_symbol: Boolean;
          signal word_access_97_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_79_complete_94_start <= ptr_deref_79_active_x_x62_symbol; -- control passed to block
          Xentry_95_symbol  <= ptr_deref_79_complete_94_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/$entry
          word_access_97: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access 
            signal word_access_97_start: Boolean;
            signal Xentry_98_symbol: Boolean;
            signal Xexit_99_symbol: Boolean;
            signal word_access_0_100_symbol : Boolean;
            signal word_access_1_105_symbol : Boolean;
            signal word_access_2_110_symbol : Boolean;
            signal word_access_3_115_symbol : Boolean;
            -- 
          begin -- 
            word_access_97_start <= Xentry_95_symbol; -- control passed to block
            Xentry_98_symbol  <= word_access_97_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/$entry
            word_access_0_100: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0 
              signal word_access_0_100_start: Boolean;
              signal Xentry_101_symbol: Boolean;
              signal Xexit_102_symbol: Boolean;
              signal cr_103_symbol : Boolean;
              signal ca_104_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_100_start <= Xentry_98_symbol; -- control passed to block
              Xentry_101_symbol  <= word_access_0_100_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/$entry
              cr_103_symbol <= Xentry_101_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/cr
              ptr_deref_79_store_0_req_1 <= cr_103_symbol; -- link to DP
              ca_104_symbol <= ptr_deref_79_store_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/ca
              Xexit_102_symbol <= ca_104_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/$exit
              word_access_0_100_symbol <= Xexit_102_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0
            word_access_1_105: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_1 
              signal word_access_1_105_start: Boolean;
              signal Xentry_106_symbol: Boolean;
              signal Xexit_107_symbol: Boolean;
              signal cr_108_symbol : Boolean;
              signal ca_109_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_105_start <= Xentry_98_symbol; -- control passed to block
              Xentry_106_symbol  <= word_access_1_105_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_1/$entry
              cr_108_symbol <= Xentry_106_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_1/cr
              ptr_deref_79_store_1_req_1 <= cr_108_symbol; -- link to DP
              ca_109_symbol <= ptr_deref_79_store_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_1/ca
              Xexit_107_symbol <= ca_109_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_1/$exit
              word_access_1_105_symbol <= Xexit_107_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_1
            word_access_2_110: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_2 
              signal word_access_2_110_start: Boolean;
              signal Xentry_111_symbol: Boolean;
              signal Xexit_112_symbol: Boolean;
              signal cr_113_symbol : Boolean;
              signal ca_114_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_110_start <= Xentry_98_symbol; -- control passed to block
              Xentry_111_symbol  <= word_access_2_110_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_2/$entry
              cr_113_symbol <= Xentry_111_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_2/cr
              ptr_deref_79_store_2_req_1 <= cr_113_symbol; -- link to DP
              ca_114_symbol <= ptr_deref_79_store_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_2/ca
              Xexit_112_symbol <= ca_114_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_2/$exit
              word_access_2_110_symbol <= Xexit_112_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_2
            word_access_3_115: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_3 
              signal word_access_3_115_start: Boolean;
              signal Xentry_116_symbol: Boolean;
              signal Xexit_117_symbol: Boolean;
              signal cr_118_symbol : Boolean;
              signal ca_119_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_115_start <= Xentry_98_symbol; -- control passed to block
              Xentry_116_symbol  <= word_access_3_115_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_3/$entry
              cr_118_symbol <= Xentry_116_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_3/cr
              ptr_deref_79_store_3_req_1 <= cr_118_symbol; -- link to DP
              ca_119_symbol <= ptr_deref_79_store_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_3/ca
              Xexit_117_symbol <= ca_119_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_3/$exit
              word_access_3_115_symbol <= Xexit_117_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_3
            Xexit_99_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/$exit 
              signal Xexit_99_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_99_predecessors(0) <= word_access_0_100_symbol;
              Xexit_99_predecessors(1) <= word_access_1_105_symbol;
              Xexit_99_predecessors(2) <= word_access_2_110_symbol;
              Xexit_99_predecessors(3) <= word_access_3_115_symbol;
              Xexit_99_join: join -- 
                port map( -- 
                  preds => Xexit_99_predecessors,
                  symbol_out => Xexit_99_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/$exit
            word_access_97_symbol <= Xexit_99_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access
          Xexit_96_symbol <= word_access_97_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/$exit
          ptr_deref_79_complete_94_symbol <= Xexit_96_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete
        assign_stmt_85_active_x_x120_symbol <= ptr_deref_84_complete_153_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_85_active_
        assign_stmt_85_completed_x_x121_symbol <= assign_stmt_85_active_x_x120_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_85_completed_
        ptr_deref_84_trigger_x_x122_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_trigger_ 
          signal ptr_deref_84_trigger_x_x122_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_84_trigger_x_x122_predecessors(0) <= ptr_deref_84_word_address_calculated_126_symbol;
          ptr_deref_84_trigger_x_x122_predecessors(1) <= ptr_deref_79_active_x_x62_symbol;
          ptr_deref_84_trigger_x_x122_join: join -- 
            port map( -- 
              preds => ptr_deref_84_trigger_x_x122_predecessors,
              symbol_out => ptr_deref_84_trigger_x_x122_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_trigger_
        ptr_deref_84_active_x_x123_symbol <= ptr_deref_84_request_127_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_active_
        ptr_deref_84_base_address_calculated_124_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_base_address_calculated
        ptr_deref_84_root_address_calculated_125_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_root_address_calculated
        ptr_deref_84_word_address_calculated_126_symbol <= ptr_deref_84_root_address_calculated_125_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_word_address_calculated
        ptr_deref_84_request_127: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request 
          signal ptr_deref_84_request_127_start: Boolean;
          signal Xentry_128_symbol: Boolean;
          signal Xexit_129_symbol: Boolean;
          signal word_access_130_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_84_request_127_start <= ptr_deref_84_trigger_x_x122_symbol; -- control passed to block
          Xentry_128_symbol  <= ptr_deref_84_request_127_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/$entry
          word_access_130: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access 
            signal word_access_130_start: Boolean;
            signal Xentry_131_symbol: Boolean;
            signal Xexit_132_symbol: Boolean;
            signal word_access_0_133_symbol : Boolean;
            signal word_access_1_138_symbol : Boolean;
            signal word_access_2_143_symbol : Boolean;
            signal word_access_3_148_symbol : Boolean;
            -- 
          begin -- 
            word_access_130_start <= Xentry_128_symbol; -- control passed to block
            Xentry_131_symbol  <= word_access_130_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/$entry
            word_access_0_133: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0 
              signal word_access_0_133_start: Boolean;
              signal Xentry_134_symbol: Boolean;
              signal Xexit_135_symbol: Boolean;
              signal rr_136_symbol : Boolean;
              signal ra_137_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_133_start <= Xentry_131_symbol; -- control passed to block
              Xentry_134_symbol  <= word_access_0_133_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/$entry
              rr_136_symbol <= Xentry_134_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/rr
              ptr_deref_84_load_0_req_0 <= rr_136_symbol; -- link to DP
              ra_137_symbol <= ptr_deref_84_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/ra
              Xexit_135_symbol <= ra_137_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/$exit
              word_access_0_133_symbol <= Xexit_135_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0
            word_access_1_138: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_1 
              signal word_access_1_138_start: Boolean;
              signal Xentry_139_symbol: Boolean;
              signal Xexit_140_symbol: Boolean;
              signal rr_141_symbol : Boolean;
              signal ra_142_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_138_start <= Xentry_131_symbol; -- control passed to block
              Xentry_139_symbol  <= word_access_1_138_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_1/$entry
              rr_141_symbol <= Xentry_139_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_1/rr
              ptr_deref_84_load_1_req_0 <= rr_141_symbol; -- link to DP
              ra_142_symbol <= ptr_deref_84_load_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_1/ra
              Xexit_140_symbol <= ra_142_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_1/$exit
              word_access_1_138_symbol <= Xexit_140_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_1
            word_access_2_143: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_2 
              signal word_access_2_143_start: Boolean;
              signal Xentry_144_symbol: Boolean;
              signal Xexit_145_symbol: Boolean;
              signal rr_146_symbol : Boolean;
              signal ra_147_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_143_start <= Xentry_131_symbol; -- control passed to block
              Xentry_144_symbol  <= word_access_2_143_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_2/$entry
              rr_146_symbol <= Xentry_144_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_2/rr
              ptr_deref_84_load_2_req_0 <= rr_146_symbol; -- link to DP
              ra_147_symbol <= ptr_deref_84_load_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_2/ra
              Xexit_145_symbol <= ra_147_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_2/$exit
              word_access_2_143_symbol <= Xexit_145_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_2
            word_access_3_148: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_3 
              signal word_access_3_148_start: Boolean;
              signal Xentry_149_symbol: Boolean;
              signal Xexit_150_symbol: Boolean;
              signal rr_151_symbol : Boolean;
              signal ra_152_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_148_start <= Xentry_131_symbol; -- control passed to block
              Xentry_149_symbol  <= word_access_3_148_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_3/$entry
              rr_151_symbol <= Xentry_149_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_3/rr
              ptr_deref_84_load_3_req_0 <= rr_151_symbol; -- link to DP
              ra_152_symbol <= ptr_deref_84_load_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_3/ra
              Xexit_150_symbol <= ra_152_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_3/$exit
              word_access_3_148_symbol <= Xexit_150_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_3
            Xexit_132_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/$exit 
              signal Xexit_132_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_132_predecessors(0) <= word_access_0_133_symbol;
              Xexit_132_predecessors(1) <= word_access_1_138_symbol;
              Xexit_132_predecessors(2) <= word_access_2_143_symbol;
              Xexit_132_predecessors(3) <= word_access_3_148_symbol;
              Xexit_132_join: join -- 
                port map( -- 
                  preds => Xexit_132_predecessors,
                  symbol_out => Xexit_132_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/$exit
            word_access_130_symbol <= Xexit_132_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access
          Xexit_129_symbol <= word_access_130_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/$exit
          ptr_deref_84_request_127_symbol <= Xexit_129_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request
        ptr_deref_84_complete_153: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete 
          signal ptr_deref_84_complete_153_start: Boolean;
          signal Xentry_154_symbol: Boolean;
          signal Xexit_155_symbol: Boolean;
          signal word_access_156_symbol : Boolean;
          signal merge_req_179_symbol : Boolean;
          signal merge_ack_180_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_84_complete_153_start <= ptr_deref_84_active_x_x123_symbol; -- control passed to block
          Xentry_154_symbol  <= ptr_deref_84_complete_153_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/$entry
          word_access_156: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access 
            signal word_access_156_start: Boolean;
            signal Xentry_157_symbol: Boolean;
            signal Xexit_158_symbol: Boolean;
            signal word_access_0_159_symbol : Boolean;
            signal word_access_1_164_symbol : Boolean;
            signal word_access_2_169_symbol : Boolean;
            signal word_access_3_174_symbol : Boolean;
            -- 
          begin -- 
            word_access_156_start <= Xentry_154_symbol; -- control passed to block
            Xentry_157_symbol  <= word_access_156_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/$entry
            word_access_0_159: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0 
              signal word_access_0_159_start: Boolean;
              signal Xentry_160_symbol: Boolean;
              signal Xexit_161_symbol: Boolean;
              signal cr_162_symbol : Boolean;
              signal ca_163_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_159_start <= Xentry_157_symbol; -- control passed to block
              Xentry_160_symbol  <= word_access_0_159_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/$entry
              cr_162_symbol <= Xentry_160_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/cr
              ptr_deref_84_load_0_req_1 <= cr_162_symbol; -- link to DP
              ca_163_symbol <= ptr_deref_84_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/ca
              Xexit_161_symbol <= ca_163_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/$exit
              word_access_0_159_symbol <= Xexit_161_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0
            word_access_1_164: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_1 
              signal word_access_1_164_start: Boolean;
              signal Xentry_165_symbol: Boolean;
              signal Xexit_166_symbol: Boolean;
              signal cr_167_symbol : Boolean;
              signal ca_168_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_164_start <= Xentry_157_symbol; -- control passed to block
              Xentry_165_symbol  <= word_access_1_164_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_1/$entry
              cr_167_symbol <= Xentry_165_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_1/cr
              ptr_deref_84_load_1_req_1 <= cr_167_symbol; -- link to DP
              ca_168_symbol <= ptr_deref_84_load_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_1/ca
              Xexit_166_symbol <= ca_168_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_1/$exit
              word_access_1_164_symbol <= Xexit_166_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_1
            word_access_2_169: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_2 
              signal word_access_2_169_start: Boolean;
              signal Xentry_170_symbol: Boolean;
              signal Xexit_171_symbol: Boolean;
              signal cr_172_symbol : Boolean;
              signal ca_173_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_169_start <= Xentry_157_symbol; -- control passed to block
              Xentry_170_symbol  <= word_access_2_169_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_2/$entry
              cr_172_symbol <= Xentry_170_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_2/cr
              ptr_deref_84_load_2_req_1 <= cr_172_symbol; -- link to DP
              ca_173_symbol <= ptr_deref_84_load_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_2/ca
              Xexit_171_symbol <= ca_173_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_2/$exit
              word_access_2_169_symbol <= Xexit_171_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_2
            word_access_3_174: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_3 
              signal word_access_3_174_start: Boolean;
              signal Xentry_175_symbol: Boolean;
              signal Xexit_176_symbol: Boolean;
              signal cr_177_symbol : Boolean;
              signal ca_178_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_174_start <= Xentry_157_symbol; -- control passed to block
              Xentry_175_symbol  <= word_access_3_174_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_3/$entry
              cr_177_symbol <= Xentry_175_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_3/cr
              ptr_deref_84_load_3_req_1 <= cr_177_symbol; -- link to DP
              ca_178_symbol <= ptr_deref_84_load_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_3/ca
              Xexit_176_symbol <= ca_178_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_3/$exit
              word_access_3_174_symbol <= Xexit_176_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_3
            Xexit_158_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/$exit 
              signal Xexit_158_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_158_predecessors(0) <= word_access_0_159_symbol;
              Xexit_158_predecessors(1) <= word_access_1_164_symbol;
              Xexit_158_predecessors(2) <= word_access_2_169_symbol;
              Xexit_158_predecessors(3) <= word_access_3_174_symbol;
              Xexit_158_join: join -- 
                port map( -- 
                  preds => Xexit_158_predecessors,
                  symbol_out => Xexit_158_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/$exit
            word_access_156_symbol <= Xexit_158_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access
          merge_req_179_symbol <= word_access_156_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/merge_req
          ptr_deref_84_gather_scatter_req_0 <= merge_req_179_symbol; -- link to DP
          merge_ack_180_symbol <= ptr_deref_84_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/merge_ack
          Xexit_155_symbol <= merge_ack_180_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/$exit
          ptr_deref_84_complete_153_symbol <= Xexit_155_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete
        assign_stmt_90_active_x_x181_symbol <= array_obj_ref_89_complete_201_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_90_active_
        assign_stmt_90_completed_x_x182_symbol <= assign_stmt_90_active_x_x181_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_90_completed_
        array_obj_ref_89_trigger_x_x183_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_trigger_
        array_obj_ref_89_active_x_x184_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_active_ 
          signal array_obj_ref_89_active_x_x184_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_89_active_x_x184_predecessors(0) <= array_obj_ref_89_trigger_x_x183_symbol;
          array_obj_ref_89_active_x_x184_predecessors(1) <= array_obj_ref_89_root_address_calculated_186_symbol;
          array_obj_ref_89_active_x_x184_join: join -- 
            port map( -- 
              preds => array_obj_ref_89_active_x_x184_predecessors,
              symbol_out => array_obj_ref_89_active_x_x184_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_active_
        array_obj_ref_89_base_address_calculated_185_symbol <= assign_stmt_85_completed_x_x121_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_address_calculated
        array_obj_ref_89_root_address_calculated_186_symbol <= array_obj_ref_89_base_plus_offset_194_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_root_address_calculated
        array_obj_ref_89_base_address_resized_187_symbol <= array_obj_ref_89_base_addr_resize_188_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_address_resized
        array_obj_ref_89_base_addr_resize_188: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize 
          signal array_obj_ref_89_base_addr_resize_188_start: Boolean;
          signal Xentry_189_symbol: Boolean;
          signal Xexit_190_symbol: Boolean;
          signal base_resize_req_191_symbol : Boolean;
          signal base_resize_ack_192_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_89_base_addr_resize_188_start <= array_obj_ref_89_base_address_calculated_185_symbol; -- control passed to block
          Xentry_189_symbol  <= array_obj_ref_89_base_addr_resize_188_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/$entry
          base_resize_req_191_symbol <= Xentry_189_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/base_resize_req
          array_obj_ref_89_base_resize_req_0 <= base_resize_req_191_symbol; -- link to DP
          base_resize_ack_192_symbol <= array_obj_ref_89_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/base_resize_ack
          Xexit_190_symbol <= base_resize_ack_192_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/$exit
          array_obj_ref_89_base_addr_resize_188_symbol <= Xexit_190_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize
        array_obj_ref_89_base_plus_offset_trigger_193_symbol <= array_obj_ref_89_base_address_resized_187_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset_trigger
        array_obj_ref_89_base_plus_offset_194: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset 
          signal array_obj_ref_89_base_plus_offset_194_start: Boolean;
          signal Xentry_195_symbol: Boolean;
          signal Xexit_196_symbol: Boolean;
          signal plus_base_rr_197_symbol : Boolean;
          signal plus_base_ra_198_symbol : Boolean;
          signal plus_base_cr_199_symbol : Boolean;
          signal plus_base_ca_200_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_89_base_plus_offset_194_start <= array_obj_ref_89_base_plus_offset_trigger_193_symbol; -- control passed to block
          Xentry_195_symbol  <= array_obj_ref_89_base_plus_offset_194_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/$entry
          plus_base_rr_197_symbol <= Xentry_195_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_rr
          array_obj_ref_89_root_address_inst_req_0 <= plus_base_rr_197_symbol; -- link to DP
          plus_base_ra_198_symbol <= array_obj_ref_89_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_ra
          plus_base_cr_199_symbol <= plus_base_ra_198_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_cr
          array_obj_ref_89_root_address_inst_req_1 <= plus_base_cr_199_symbol; -- link to DP
          plus_base_ca_200_symbol <= array_obj_ref_89_root_address_inst_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_ca
          Xexit_196_symbol <= plus_base_ca_200_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/$exit
          array_obj_ref_89_base_plus_offset_194_symbol <= Xexit_196_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset
        array_obj_ref_89_complete_201: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete 
          signal array_obj_ref_89_complete_201_start: Boolean;
          signal Xentry_202_symbol: Boolean;
          signal Xexit_203_symbol: Boolean;
          signal final_reg_req_204_symbol : Boolean;
          signal final_reg_ack_205_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_89_complete_201_start <= array_obj_ref_89_active_x_x184_symbol; -- control passed to block
          Xentry_202_symbol  <= array_obj_ref_89_complete_201_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/$entry
          final_reg_req_204_symbol <= Xentry_202_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/final_reg_req
          array_obj_ref_89_final_reg_req_0 <= final_reg_req_204_symbol; -- link to DP
          final_reg_ack_205_symbol <= array_obj_ref_89_final_reg_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/final_reg_ack
          Xexit_203_symbol <= final_reg_ack_205_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/$exit
          array_obj_ref_89_complete_201_symbol <= Xexit_203_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete
        assign_stmt_94_active_x_x206_symbol <= ptr_deref_93_complete_282_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_94_active_
        assign_stmt_94_completed_x_x207_symbol <= assign_stmt_94_active_x_x206_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_94_completed_
        ptr_deref_93_trigger_x_x208_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_trigger_ 
          signal ptr_deref_93_trigger_x_x208_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          ptr_deref_93_trigger_x_x208_predecessors(0) <= ptr_deref_93_word_address_calculated_213_symbol;
          ptr_deref_93_trigger_x_x208_predecessors(1) <= ptr_deref_93_base_address_calculated_210_symbol;
          ptr_deref_93_trigger_x_x208_predecessors(2) <= ptr_deref_79_active_x_x62_symbol;
          ptr_deref_93_trigger_x_x208_join: join -- 
            port map( -- 
              preds => ptr_deref_93_trigger_x_x208_predecessors,
              symbol_out => ptr_deref_93_trigger_x_x208_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_trigger_
        ptr_deref_93_active_x_x209_symbol <= ptr_deref_93_request_256_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_active_
        ptr_deref_93_base_address_calculated_210_symbol <= simple_obj_ref_92_complete_211_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_address_calculated
        simple_obj_ref_92_complete_211_symbol <= assign_stmt_90_completed_x_x182_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_92_complete
        ptr_deref_93_root_address_calculated_212_symbol <= ptr_deref_93_base_plus_offset_220_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_root_address_calculated
        ptr_deref_93_word_address_calculated_213_symbol <= ptr_deref_93_word_addrgen_225_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_address_calculated
        ptr_deref_93_base_address_resized_214_symbol <= ptr_deref_93_base_addr_resize_215_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_address_resized
        ptr_deref_93_base_addr_resize_215: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize 
          signal ptr_deref_93_base_addr_resize_215_start: Boolean;
          signal Xentry_216_symbol: Boolean;
          signal Xexit_217_symbol: Boolean;
          signal base_resize_req_218_symbol : Boolean;
          signal base_resize_ack_219_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_base_addr_resize_215_start <= ptr_deref_93_base_address_calculated_210_symbol; -- control passed to block
          Xentry_216_symbol  <= ptr_deref_93_base_addr_resize_215_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/$entry
          base_resize_req_218_symbol <= Xentry_216_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/base_resize_req
          ptr_deref_93_base_resize_req_0 <= base_resize_req_218_symbol; -- link to DP
          base_resize_ack_219_symbol <= ptr_deref_93_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/base_resize_ack
          Xexit_217_symbol <= base_resize_ack_219_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/$exit
          ptr_deref_93_base_addr_resize_215_symbol <= Xexit_217_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize
        ptr_deref_93_base_plus_offset_220: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset 
          signal ptr_deref_93_base_plus_offset_220_start: Boolean;
          signal Xentry_221_symbol: Boolean;
          signal Xexit_222_symbol: Boolean;
          signal sum_rename_req_223_symbol : Boolean;
          signal sum_rename_ack_224_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_base_plus_offset_220_start <= ptr_deref_93_base_address_resized_214_symbol; -- control passed to block
          Xentry_221_symbol  <= ptr_deref_93_base_plus_offset_220_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/$entry
          sum_rename_req_223_symbol <= Xentry_221_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/sum_rename_req
          ptr_deref_93_root_address_inst_req_0 <= sum_rename_req_223_symbol; -- link to DP
          sum_rename_ack_224_symbol <= ptr_deref_93_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/sum_rename_ack
          Xexit_222_symbol <= sum_rename_ack_224_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/$exit
          ptr_deref_93_base_plus_offset_220_symbol <= Xexit_222_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset
        ptr_deref_93_word_addrgen_225: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen 
          signal ptr_deref_93_word_addrgen_225_start: Boolean;
          signal Xentry_226_symbol: Boolean;
          signal Xexit_227_symbol: Boolean;
          signal word_0_228_symbol : Boolean;
          signal word_1_235_symbol : Boolean;
          signal word_2_242_symbol : Boolean;
          signal word_3_249_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_word_addrgen_225_start <= ptr_deref_93_root_address_calculated_212_symbol; -- control passed to block
          Xentry_226_symbol  <= ptr_deref_93_word_addrgen_225_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/$entry
          word_0_228: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0 
            signal word_0_228_start: Boolean;
            signal Xentry_229_symbol: Boolean;
            signal Xexit_230_symbol: Boolean;
            signal rr_231_symbol : Boolean;
            signal ra_232_symbol : Boolean;
            signal cr_233_symbol : Boolean;
            signal ca_234_symbol : Boolean;
            -- 
          begin -- 
            word_0_228_start <= Xentry_226_symbol; -- control passed to block
            Xentry_229_symbol  <= word_0_228_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0/$entry
            rr_231_symbol <= Xentry_229_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0/rr
            ptr_deref_93_addr_0_req_0 <= rr_231_symbol; -- link to DP
            ra_232_symbol <= ptr_deref_93_addr_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0/ra
            cr_233_symbol <= ra_232_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0/cr
            ptr_deref_93_addr_0_req_1 <= cr_233_symbol; -- link to DP
            ca_234_symbol <= ptr_deref_93_addr_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0/ca
            Xexit_230_symbol <= ca_234_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0/$exit
            word_0_228_symbol <= Xexit_230_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_0
          word_1_235: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1 
            signal word_1_235_start: Boolean;
            signal Xentry_236_symbol: Boolean;
            signal Xexit_237_symbol: Boolean;
            signal rr_238_symbol : Boolean;
            signal ra_239_symbol : Boolean;
            signal cr_240_symbol : Boolean;
            signal ca_241_symbol : Boolean;
            -- 
          begin -- 
            word_1_235_start <= Xentry_226_symbol; -- control passed to block
            Xentry_236_symbol  <= word_1_235_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1/$entry
            rr_238_symbol <= Xentry_236_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1/rr
            ptr_deref_93_addr_1_req_0 <= rr_238_symbol; -- link to DP
            ra_239_symbol <= ptr_deref_93_addr_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1/ra
            cr_240_symbol <= ra_239_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1/cr
            ptr_deref_93_addr_1_req_1 <= cr_240_symbol; -- link to DP
            ca_241_symbol <= ptr_deref_93_addr_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1/ca
            Xexit_237_symbol <= ca_241_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1/$exit
            word_1_235_symbol <= Xexit_237_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_1
          word_2_242: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2 
            signal word_2_242_start: Boolean;
            signal Xentry_243_symbol: Boolean;
            signal Xexit_244_symbol: Boolean;
            signal rr_245_symbol : Boolean;
            signal ra_246_symbol : Boolean;
            signal cr_247_symbol : Boolean;
            signal ca_248_symbol : Boolean;
            -- 
          begin -- 
            word_2_242_start <= Xentry_226_symbol; -- control passed to block
            Xentry_243_symbol  <= word_2_242_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2/$entry
            rr_245_symbol <= Xentry_243_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2/rr
            ptr_deref_93_addr_2_req_0 <= rr_245_symbol; -- link to DP
            ra_246_symbol <= ptr_deref_93_addr_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2/ra
            cr_247_symbol <= ra_246_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2/cr
            ptr_deref_93_addr_2_req_1 <= cr_247_symbol; -- link to DP
            ca_248_symbol <= ptr_deref_93_addr_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2/ca
            Xexit_244_symbol <= ca_248_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2/$exit
            word_2_242_symbol <= Xexit_244_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_2
          word_3_249: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3 
            signal word_3_249_start: Boolean;
            signal Xentry_250_symbol: Boolean;
            signal Xexit_251_symbol: Boolean;
            signal rr_252_symbol : Boolean;
            signal ra_253_symbol : Boolean;
            signal cr_254_symbol : Boolean;
            signal ca_255_symbol : Boolean;
            -- 
          begin -- 
            word_3_249_start <= Xentry_226_symbol; -- control passed to block
            Xentry_250_symbol  <= word_3_249_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3/$entry
            rr_252_symbol <= Xentry_250_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3/rr
            ptr_deref_93_addr_3_req_0 <= rr_252_symbol; -- link to DP
            ra_253_symbol <= ptr_deref_93_addr_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3/ra
            cr_254_symbol <= ra_253_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3/cr
            ptr_deref_93_addr_3_req_1 <= cr_254_symbol; -- link to DP
            ca_255_symbol <= ptr_deref_93_addr_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3/ca
            Xexit_251_symbol <= ca_255_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3/$exit
            word_3_249_symbol <= Xexit_251_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/word_3
          Xexit_227_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/$exit 
            signal Xexit_227_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_227_predecessors(0) <= word_0_228_symbol;
            Xexit_227_predecessors(1) <= word_1_235_symbol;
            Xexit_227_predecessors(2) <= word_2_242_symbol;
            Xexit_227_predecessors(3) <= word_3_249_symbol;
            Xexit_227_join: join -- 
              port map( -- 
                preds => Xexit_227_predecessors,
                symbol_out => Xexit_227_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/$exit
          ptr_deref_93_word_addrgen_225_symbol <= Xexit_227_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen
        ptr_deref_93_request_256: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request 
          signal ptr_deref_93_request_256_start: Boolean;
          signal Xentry_257_symbol: Boolean;
          signal Xexit_258_symbol: Boolean;
          signal word_access_259_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_request_256_start <= ptr_deref_93_trigger_x_x208_symbol; -- control passed to block
          Xentry_257_symbol  <= ptr_deref_93_request_256_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/$entry
          word_access_259: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access 
            signal word_access_259_start: Boolean;
            signal Xentry_260_symbol: Boolean;
            signal Xexit_261_symbol: Boolean;
            signal word_access_0_262_symbol : Boolean;
            signal word_access_1_267_symbol : Boolean;
            signal word_access_2_272_symbol : Boolean;
            signal word_access_3_277_symbol : Boolean;
            -- 
          begin -- 
            word_access_259_start <= Xentry_257_symbol; -- control passed to block
            Xentry_260_symbol  <= word_access_259_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/$entry
            word_access_0_262: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0 
              signal word_access_0_262_start: Boolean;
              signal Xentry_263_symbol: Boolean;
              signal Xexit_264_symbol: Boolean;
              signal rr_265_symbol : Boolean;
              signal ra_266_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_262_start <= Xentry_260_symbol; -- control passed to block
              Xentry_263_symbol  <= word_access_0_262_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/$entry
              rr_265_symbol <= Xentry_263_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/rr
              ptr_deref_93_load_0_req_0 <= rr_265_symbol; -- link to DP
              ra_266_symbol <= ptr_deref_93_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/ra
              Xexit_264_symbol <= ra_266_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/$exit
              word_access_0_262_symbol <= Xexit_264_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0
            word_access_1_267: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_1 
              signal word_access_1_267_start: Boolean;
              signal Xentry_268_symbol: Boolean;
              signal Xexit_269_symbol: Boolean;
              signal rr_270_symbol : Boolean;
              signal ra_271_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_267_start <= Xentry_260_symbol; -- control passed to block
              Xentry_268_symbol  <= word_access_1_267_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_1/$entry
              rr_270_symbol <= Xentry_268_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_1/rr
              ptr_deref_93_load_1_req_0 <= rr_270_symbol; -- link to DP
              ra_271_symbol <= ptr_deref_93_load_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_1/ra
              Xexit_269_symbol <= ra_271_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_1/$exit
              word_access_1_267_symbol <= Xexit_269_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_1
            word_access_2_272: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_2 
              signal word_access_2_272_start: Boolean;
              signal Xentry_273_symbol: Boolean;
              signal Xexit_274_symbol: Boolean;
              signal rr_275_symbol : Boolean;
              signal ra_276_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_272_start <= Xentry_260_symbol; -- control passed to block
              Xentry_273_symbol  <= word_access_2_272_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_2/$entry
              rr_275_symbol <= Xentry_273_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_2/rr
              ptr_deref_93_load_2_req_0 <= rr_275_symbol; -- link to DP
              ra_276_symbol <= ptr_deref_93_load_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_2/ra
              Xexit_274_symbol <= ra_276_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_2/$exit
              word_access_2_272_symbol <= Xexit_274_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_2
            word_access_3_277: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_3 
              signal word_access_3_277_start: Boolean;
              signal Xentry_278_symbol: Boolean;
              signal Xexit_279_symbol: Boolean;
              signal rr_280_symbol : Boolean;
              signal ra_281_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_277_start <= Xentry_260_symbol; -- control passed to block
              Xentry_278_symbol  <= word_access_3_277_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_3/$entry
              rr_280_symbol <= Xentry_278_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_3/rr
              ptr_deref_93_load_3_req_0 <= rr_280_symbol; -- link to DP
              ra_281_symbol <= ptr_deref_93_load_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_3/ra
              Xexit_279_symbol <= ra_281_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_3/$exit
              word_access_3_277_symbol <= Xexit_279_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_3
            Xexit_261_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/$exit 
              signal Xexit_261_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_261_predecessors(0) <= word_access_0_262_symbol;
              Xexit_261_predecessors(1) <= word_access_1_267_symbol;
              Xexit_261_predecessors(2) <= word_access_2_272_symbol;
              Xexit_261_predecessors(3) <= word_access_3_277_symbol;
              Xexit_261_join: join -- 
                port map( -- 
                  preds => Xexit_261_predecessors,
                  symbol_out => Xexit_261_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/$exit
            word_access_259_symbol <= Xexit_261_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access
          Xexit_258_symbol <= word_access_259_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/$exit
          ptr_deref_93_request_256_symbol <= Xexit_258_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request
        ptr_deref_93_complete_282: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete 
          signal ptr_deref_93_complete_282_start: Boolean;
          signal Xentry_283_symbol: Boolean;
          signal Xexit_284_symbol: Boolean;
          signal word_access_285_symbol : Boolean;
          signal merge_req_308_symbol : Boolean;
          signal merge_ack_309_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_complete_282_start <= ptr_deref_93_active_x_x209_symbol; -- control passed to block
          Xentry_283_symbol  <= ptr_deref_93_complete_282_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/$entry
          word_access_285: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access 
            signal word_access_285_start: Boolean;
            signal Xentry_286_symbol: Boolean;
            signal Xexit_287_symbol: Boolean;
            signal word_access_0_288_symbol : Boolean;
            signal word_access_1_293_symbol : Boolean;
            signal word_access_2_298_symbol : Boolean;
            signal word_access_3_303_symbol : Boolean;
            -- 
          begin -- 
            word_access_285_start <= Xentry_283_symbol; -- control passed to block
            Xentry_286_symbol  <= word_access_285_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/$entry
            word_access_0_288: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0 
              signal word_access_0_288_start: Boolean;
              signal Xentry_289_symbol: Boolean;
              signal Xexit_290_symbol: Boolean;
              signal cr_291_symbol : Boolean;
              signal ca_292_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_288_start <= Xentry_286_symbol; -- control passed to block
              Xentry_289_symbol  <= word_access_0_288_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/$entry
              cr_291_symbol <= Xentry_289_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/cr
              ptr_deref_93_load_0_req_1 <= cr_291_symbol; -- link to DP
              ca_292_symbol <= ptr_deref_93_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/ca
              Xexit_290_symbol <= ca_292_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/$exit
              word_access_0_288_symbol <= Xexit_290_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0
            word_access_1_293: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_1 
              signal word_access_1_293_start: Boolean;
              signal Xentry_294_symbol: Boolean;
              signal Xexit_295_symbol: Boolean;
              signal cr_296_symbol : Boolean;
              signal ca_297_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_293_start <= Xentry_286_symbol; -- control passed to block
              Xentry_294_symbol  <= word_access_1_293_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_1/$entry
              cr_296_symbol <= Xentry_294_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_1/cr
              ptr_deref_93_load_1_req_1 <= cr_296_symbol; -- link to DP
              ca_297_symbol <= ptr_deref_93_load_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_1/ca
              Xexit_295_symbol <= ca_297_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_1/$exit
              word_access_1_293_symbol <= Xexit_295_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_1
            word_access_2_298: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_2 
              signal word_access_2_298_start: Boolean;
              signal Xentry_299_symbol: Boolean;
              signal Xexit_300_symbol: Boolean;
              signal cr_301_symbol : Boolean;
              signal ca_302_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_298_start <= Xentry_286_symbol; -- control passed to block
              Xentry_299_symbol  <= word_access_2_298_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_2/$entry
              cr_301_symbol <= Xentry_299_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_2/cr
              ptr_deref_93_load_2_req_1 <= cr_301_symbol; -- link to DP
              ca_302_symbol <= ptr_deref_93_load_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_2/ca
              Xexit_300_symbol <= ca_302_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_2/$exit
              word_access_2_298_symbol <= Xexit_300_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_2
            word_access_3_303: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_3 
              signal word_access_3_303_start: Boolean;
              signal Xentry_304_symbol: Boolean;
              signal Xexit_305_symbol: Boolean;
              signal cr_306_symbol : Boolean;
              signal ca_307_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_303_start <= Xentry_286_symbol; -- control passed to block
              Xentry_304_symbol  <= word_access_3_303_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_3/$entry
              cr_306_symbol <= Xentry_304_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_3/cr
              ptr_deref_93_load_3_req_1 <= cr_306_symbol; -- link to DP
              ca_307_symbol <= ptr_deref_93_load_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_3/ca
              Xexit_305_symbol <= ca_307_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_3/$exit
              word_access_3_303_symbol <= Xexit_305_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_3
            Xexit_287_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/$exit 
              signal Xexit_287_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_287_predecessors(0) <= word_access_0_288_symbol;
              Xexit_287_predecessors(1) <= word_access_1_293_symbol;
              Xexit_287_predecessors(2) <= word_access_2_298_symbol;
              Xexit_287_predecessors(3) <= word_access_3_303_symbol;
              Xexit_287_join: join -- 
                port map( -- 
                  preds => Xexit_287_predecessors,
                  symbol_out => Xexit_287_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/$exit
            word_access_285_symbol <= Xexit_287_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access
          merge_req_308_symbol <= word_access_285_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/merge_req
          ptr_deref_93_gather_scatter_req_0 <= merge_req_308_symbol; -- link to DP
          merge_ack_309_symbol <= ptr_deref_93_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/merge_ack
          Xexit_284_symbol <= merge_ack_309_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/$exit
          ptr_deref_93_complete_282_symbol <= Xexit_284_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete
        assign_stmt_99_active_x_x310_symbol <= binary_98_complete_315_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_99_active_
        assign_stmt_99_completed_x_x311_symbol <= assign_stmt_99_active_x_x310_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_99_completed_
        binary_98_active_x_x312_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_active_ 
          signal binary_98_active_x_x312_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_98_active_x_x312_predecessors(0) <= binary_98_trigger_x_x313_symbol;
          binary_98_active_x_x312_predecessors(1) <= simple_obj_ref_97_complete_314_symbol;
          binary_98_active_x_x312_join: join -- 
            port map( -- 
              preds => binary_98_active_x_x312_predecessors,
              symbol_out => binary_98_active_x_x312_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_active_
        binary_98_trigger_x_x313_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_trigger_
        simple_obj_ref_97_complete_314_symbol <= assign_stmt_94_completed_x_x207_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_97_complete
        binary_98_complete_315: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete 
          signal binary_98_complete_315_start: Boolean;
          signal Xentry_316_symbol: Boolean;
          signal Xexit_317_symbol: Boolean;
          signal rr_318_symbol : Boolean;
          signal ra_319_symbol : Boolean;
          signal cr_320_symbol : Boolean;
          signal ca_321_symbol : Boolean;
          -- 
        begin -- 
          binary_98_complete_315_start <= binary_98_active_x_x312_symbol; -- control passed to block
          Xentry_316_symbol  <= binary_98_complete_315_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/$entry
          rr_318_symbol <= Xentry_316_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/rr
          binary_98_inst_req_0 <= rr_318_symbol; -- link to DP
          ra_319_symbol <= binary_98_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/ra
          cr_320_symbol <= ra_319_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/cr
          binary_98_inst_req_1 <= cr_320_symbol; -- link to DP
          ca_321_symbol <= binary_98_inst_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/ca
          Xexit_317_symbol <= ca_321_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/$exit
          binary_98_complete_315_symbol <= Xexit_317_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete
        assign_stmt_103_active_x_x322_symbol <= ptr_deref_102_complete_355_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_103_active_
        assign_stmt_103_completed_x_x323_symbol <= assign_stmt_103_active_x_x322_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_103_completed_
        ptr_deref_102_trigger_x_x324_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_trigger_ 
          signal ptr_deref_102_trigger_x_x324_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_102_trigger_x_x324_predecessors(0) <= ptr_deref_102_word_address_calculated_328_symbol;
          ptr_deref_102_trigger_x_x324_predecessors(1) <= ptr_deref_79_active_x_x62_symbol;
          ptr_deref_102_trigger_x_x324_join: join -- 
            port map( -- 
              preds => ptr_deref_102_trigger_x_x324_predecessors,
              symbol_out => ptr_deref_102_trigger_x_x324_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_trigger_
        ptr_deref_102_active_x_x325_symbol <= ptr_deref_102_request_329_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_active_
        ptr_deref_102_base_address_calculated_326_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_base_address_calculated
        ptr_deref_102_root_address_calculated_327_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_root_address_calculated
        ptr_deref_102_word_address_calculated_328_symbol <= ptr_deref_102_root_address_calculated_327_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_word_address_calculated
        ptr_deref_102_request_329: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request 
          signal ptr_deref_102_request_329_start: Boolean;
          signal Xentry_330_symbol: Boolean;
          signal Xexit_331_symbol: Boolean;
          signal word_access_332_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_102_request_329_start <= ptr_deref_102_trigger_x_x324_symbol; -- control passed to block
          Xentry_330_symbol  <= ptr_deref_102_request_329_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/$entry
          word_access_332: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access 
            signal word_access_332_start: Boolean;
            signal Xentry_333_symbol: Boolean;
            signal Xexit_334_symbol: Boolean;
            signal word_access_0_335_symbol : Boolean;
            signal word_access_1_340_symbol : Boolean;
            signal word_access_2_345_symbol : Boolean;
            signal word_access_3_350_symbol : Boolean;
            -- 
          begin -- 
            word_access_332_start <= Xentry_330_symbol; -- control passed to block
            Xentry_333_symbol  <= word_access_332_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/$entry
            word_access_0_335: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0 
              signal word_access_0_335_start: Boolean;
              signal Xentry_336_symbol: Boolean;
              signal Xexit_337_symbol: Boolean;
              signal rr_338_symbol : Boolean;
              signal ra_339_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_335_start <= Xentry_333_symbol; -- control passed to block
              Xentry_336_symbol  <= word_access_0_335_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/$entry
              rr_338_symbol <= Xentry_336_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/rr
              ptr_deref_102_load_0_req_0 <= rr_338_symbol; -- link to DP
              ra_339_symbol <= ptr_deref_102_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/ra
              Xexit_337_symbol <= ra_339_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/$exit
              word_access_0_335_symbol <= Xexit_337_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0
            word_access_1_340: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_1 
              signal word_access_1_340_start: Boolean;
              signal Xentry_341_symbol: Boolean;
              signal Xexit_342_symbol: Boolean;
              signal rr_343_symbol : Boolean;
              signal ra_344_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_340_start <= Xentry_333_symbol; -- control passed to block
              Xentry_341_symbol  <= word_access_1_340_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_1/$entry
              rr_343_symbol <= Xentry_341_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_1/rr
              ptr_deref_102_load_1_req_0 <= rr_343_symbol; -- link to DP
              ra_344_symbol <= ptr_deref_102_load_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_1/ra
              Xexit_342_symbol <= ra_344_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_1/$exit
              word_access_1_340_symbol <= Xexit_342_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_1
            word_access_2_345: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_2 
              signal word_access_2_345_start: Boolean;
              signal Xentry_346_symbol: Boolean;
              signal Xexit_347_symbol: Boolean;
              signal rr_348_symbol : Boolean;
              signal ra_349_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_345_start <= Xentry_333_symbol; -- control passed to block
              Xentry_346_symbol  <= word_access_2_345_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_2/$entry
              rr_348_symbol <= Xentry_346_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_2/rr
              ptr_deref_102_load_2_req_0 <= rr_348_symbol; -- link to DP
              ra_349_symbol <= ptr_deref_102_load_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_2/ra
              Xexit_347_symbol <= ra_349_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_2/$exit
              word_access_2_345_symbol <= Xexit_347_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_2
            word_access_3_350: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_3 
              signal word_access_3_350_start: Boolean;
              signal Xentry_351_symbol: Boolean;
              signal Xexit_352_symbol: Boolean;
              signal rr_353_symbol : Boolean;
              signal ra_354_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_350_start <= Xentry_333_symbol; -- control passed to block
              Xentry_351_symbol  <= word_access_3_350_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_3/$entry
              rr_353_symbol <= Xentry_351_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_3/rr
              ptr_deref_102_load_3_req_0 <= rr_353_symbol; -- link to DP
              ra_354_symbol <= ptr_deref_102_load_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_3/ra
              Xexit_352_symbol <= ra_354_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_3/$exit
              word_access_3_350_symbol <= Xexit_352_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_3
            Xexit_334_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/$exit 
              signal Xexit_334_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_334_predecessors(0) <= word_access_0_335_symbol;
              Xexit_334_predecessors(1) <= word_access_1_340_symbol;
              Xexit_334_predecessors(2) <= word_access_2_345_symbol;
              Xexit_334_predecessors(3) <= word_access_3_350_symbol;
              Xexit_334_join: join -- 
                port map( -- 
                  preds => Xexit_334_predecessors,
                  symbol_out => Xexit_334_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/$exit
            word_access_332_symbol <= Xexit_334_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access
          Xexit_331_symbol <= word_access_332_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/$exit
          ptr_deref_102_request_329_symbol <= Xexit_331_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request
        ptr_deref_102_complete_355: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete 
          signal ptr_deref_102_complete_355_start: Boolean;
          signal Xentry_356_symbol: Boolean;
          signal Xexit_357_symbol: Boolean;
          signal word_access_358_symbol : Boolean;
          signal merge_req_381_symbol : Boolean;
          signal merge_ack_382_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_102_complete_355_start <= ptr_deref_102_active_x_x325_symbol; -- control passed to block
          Xentry_356_symbol  <= ptr_deref_102_complete_355_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/$entry
          word_access_358: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access 
            signal word_access_358_start: Boolean;
            signal Xentry_359_symbol: Boolean;
            signal Xexit_360_symbol: Boolean;
            signal word_access_0_361_symbol : Boolean;
            signal word_access_1_366_symbol : Boolean;
            signal word_access_2_371_symbol : Boolean;
            signal word_access_3_376_symbol : Boolean;
            -- 
          begin -- 
            word_access_358_start <= Xentry_356_symbol; -- control passed to block
            Xentry_359_symbol  <= word_access_358_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/$entry
            word_access_0_361: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0 
              signal word_access_0_361_start: Boolean;
              signal Xentry_362_symbol: Boolean;
              signal Xexit_363_symbol: Boolean;
              signal cr_364_symbol : Boolean;
              signal ca_365_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_361_start <= Xentry_359_symbol; -- control passed to block
              Xentry_362_symbol  <= word_access_0_361_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/$entry
              cr_364_symbol <= Xentry_362_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/cr
              ptr_deref_102_load_0_req_1 <= cr_364_symbol; -- link to DP
              ca_365_symbol <= ptr_deref_102_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/ca
              Xexit_363_symbol <= ca_365_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/$exit
              word_access_0_361_symbol <= Xexit_363_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0
            word_access_1_366: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_1 
              signal word_access_1_366_start: Boolean;
              signal Xentry_367_symbol: Boolean;
              signal Xexit_368_symbol: Boolean;
              signal cr_369_symbol : Boolean;
              signal ca_370_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_366_start <= Xentry_359_symbol; -- control passed to block
              Xentry_367_symbol  <= word_access_1_366_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_1/$entry
              cr_369_symbol <= Xentry_367_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_1/cr
              ptr_deref_102_load_1_req_1 <= cr_369_symbol; -- link to DP
              ca_370_symbol <= ptr_deref_102_load_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_1/ca
              Xexit_368_symbol <= ca_370_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_1/$exit
              word_access_1_366_symbol <= Xexit_368_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_1
            word_access_2_371: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_2 
              signal word_access_2_371_start: Boolean;
              signal Xentry_372_symbol: Boolean;
              signal Xexit_373_symbol: Boolean;
              signal cr_374_symbol : Boolean;
              signal ca_375_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_371_start <= Xentry_359_symbol; -- control passed to block
              Xentry_372_symbol  <= word_access_2_371_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_2/$entry
              cr_374_symbol <= Xentry_372_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_2/cr
              ptr_deref_102_load_2_req_1 <= cr_374_symbol; -- link to DP
              ca_375_symbol <= ptr_deref_102_load_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_2/ca
              Xexit_373_symbol <= ca_375_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_2/$exit
              word_access_2_371_symbol <= Xexit_373_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_2
            word_access_3_376: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_3 
              signal word_access_3_376_start: Boolean;
              signal Xentry_377_symbol: Boolean;
              signal Xexit_378_symbol: Boolean;
              signal cr_379_symbol : Boolean;
              signal ca_380_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_376_start <= Xentry_359_symbol; -- control passed to block
              Xentry_377_symbol  <= word_access_3_376_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_3/$entry
              cr_379_symbol <= Xentry_377_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_3/cr
              ptr_deref_102_load_3_req_1 <= cr_379_symbol; -- link to DP
              ca_380_symbol <= ptr_deref_102_load_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_3/ca
              Xexit_378_symbol <= ca_380_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_3/$exit
              word_access_3_376_symbol <= Xexit_378_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_3
            Xexit_360_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/$exit 
              signal Xexit_360_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_360_predecessors(0) <= word_access_0_361_symbol;
              Xexit_360_predecessors(1) <= word_access_1_366_symbol;
              Xexit_360_predecessors(2) <= word_access_2_371_symbol;
              Xexit_360_predecessors(3) <= word_access_3_376_symbol;
              Xexit_360_join: join -- 
                port map( -- 
                  preds => Xexit_360_predecessors,
                  symbol_out => Xexit_360_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/$exit
            word_access_358_symbol <= Xexit_360_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access
          merge_req_381_symbol <= word_access_358_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/merge_req
          ptr_deref_102_gather_scatter_req_0 <= merge_req_381_symbol; -- link to DP
          merge_ack_382_symbol <= ptr_deref_102_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/merge_ack
          Xexit_357_symbol <= merge_ack_382_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/$exit
          ptr_deref_102_complete_355_symbol <= Xexit_357_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete
        assign_stmt_108_active_x_x383_symbol <= array_obj_ref_107_complete_403_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_108_active_
        assign_stmt_108_completed_x_x384_symbol <= assign_stmt_108_active_x_x383_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_108_completed_
        array_obj_ref_107_trigger_x_x385_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_trigger_
        array_obj_ref_107_active_x_x386_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_active_ 
          signal array_obj_ref_107_active_x_x386_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_107_active_x_x386_predecessors(0) <= array_obj_ref_107_trigger_x_x385_symbol;
          array_obj_ref_107_active_x_x386_predecessors(1) <= array_obj_ref_107_root_address_calculated_388_symbol;
          array_obj_ref_107_active_x_x386_join: join -- 
            port map( -- 
              preds => array_obj_ref_107_active_x_x386_predecessors,
              symbol_out => array_obj_ref_107_active_x_x386_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_active_
        array_obj_ref_107_base_address_calculated_387_symbol <= assign_stmt_103_completed_x_x323_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_address_calculated
        array_obj_ref_107_root_address_calculated_388_symbol <= array_obj_ref_107_base_plus_offset_396_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_root_address_calculated
        array_obj_ref_107_base_address_resized_389_symbol <= array_obj_ref_107_base_addr_resize_390_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_address_resized
        array_obj_ref_107_base_addr_resize_390: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize 
          signal array_obj_ref_107_base_addr_resize_390_start: Boolean;
          signal Xentry_391_symbol: Boolean;
          signal Xexit_392_symbol: Boolean;
          signal base_resize_req_393_symbol : Boolean;
          signal base_resize_ack_394_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_107_base_addr_resize_390_start <= array_obj_ref_107_base_address_calculated_387_symbol; -- control passed to block
          Xentry_391_symbol  <= array_obj_ref_107_base_addr_resize_390_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/$entry
          base_resize_req_393_symbol <= Xentry_391_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/base_resize_req
          array_obj_ref_107_base_resize_req_0 <= base_resize_req_393_symbol; -- link to DP
          base_resize_ack_394_symbol <= array_obj_ref_107_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/base_resize_ack
          Xexit_392_symbol <= base_resize_ack_394_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/$exit
          array_obj_ref_107_base_addr_resize_390_symbol <= Xexit_392_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize
        array_obj_ref_107_base_plus_offset_trigger_395_symbol <= array_obj_ref_107_base_address_resized_389_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset_trigger
        array_obj_ref_107_base_plus_offset_396: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset 
          signal array_obj_ref_107_base_plus_offset_396_start: Boolean;
          signal Xentry_397_symbol: Boolean;
          signal Xexit_398_symbol: Boolean;
          signal plus_base_rr_399_symbol : Boolean;
          signal plus_base_ra_400_symbol : Boolean;
          signal plus_base_cr_401_symbol : Boolean;
          signal plus_base_ca_402_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_107_base_plus_offset_396_start <= array_obj_ref_107_base_plus_offset_trigger_395_symbol; -- control passed to block
          Xentry_397_symbol  <= array_obj_ref_107_base_plus_offset_396_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/$entry
          plus_base_rr_399_symbol <= Xentry_397_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_rr
          array_obj_ref_107_root_address_inst_req_0 <= plus_base_rr_399_symbol; -- link to DP
          plus_base_ra_400_symbol <= array_obj_ref_107_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_ra
          plus_base_cr_401_symbol <= plus_base_ra_400_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_cr
          array_obj_ref_107_root_address_inst_req_1 <= plus_base_cr_401_symbol; -- link to DP
          plus_base_ca_402_symbol <= array_obj_ref_107_root_address_inst_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_ca
          Xexit_398_symbol <= plus_base_ca_402_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/$exit
          array_obj_ref_107_base_plus_offset_396_symbol <= Xexit_398_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset
        array_obj_ref_107_complete_403: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete 
          signal array_obj_ref_107_complete_403_start: Boolean;
          signal Xentry_404_symbol: Boolean;
          signal Xexit_405_symbol: Boolean;
          signal final_reg_req_406_symbol : Boolean;
          signal final_reg_ack_407_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_107_complete_403_start <= array_obj_ref_107_active_x_x386_symbol; -- control passed to block
          Xentry_404_symbol  <= array_obj_ref_107_complete_403_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/$entry
          final_reg_req_406_symbol <= Xentry_404_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/final_reg_req
          array_obj_ref_107_final_reg_req_0 <= final_reg_req_406_symbol; -- link to DP
          final_reg_ack_407_symbol <= array_obj_ref_107_final_reg_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/final_reg_ack
          Xexit_405_symbol <= final_reg_ack_407_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/$exit
          array_obj_ref_107_complete_403_symbol <= Xexit_405_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete
        assign_stmt_112_active_x_x408_symbol <= simple_obj_ref_111_complete_410_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_112_active_
        assign_stmt_112_completed_x_x409_symbol <= ptr_deref_110_complete_487_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_112_completed_
        simple_obj_ref_111_complete_410_symbol <= assign_stmt_99_completed_x_x311_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_111_complete
        ptr_deref_110_trigger_x_x411_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_trigger_ 
          signal ptr_deref_110_trigger_x_x411_predecessors: BooleanArray(5 downto 0);
          -- 
        begin -- 
          ptr_deref_110_trigger_x_x411_predecessors(0) <= ptr_deref_110_word_address_calculated_416_symbol;
          ptr_deref_110_trigger_x_x411_predecessors(1) <= ptr_deref_110_base_address_calculated_413_symbol;
          ptr_deref_110_trigger_x_x411_predecessors(2) <= assign_stmt_112_active_x_x408_symbol;
          ptr_deref_110_trigger_x_x411_predecessors(3) <= ptr_deref_84_active_x_x123_symbol;
          ptr_deref_110_trigger_x_x411_predecessors(4) <= ptr_deref_93_active_x_x209_symbol;
          ptr_deref_110_trigger_x_x411_predecessors(5) <= ptr_deref_102_active_x_x325_symbol;
          ptr_deref_110_trigger_x_x411_join: join -- 
            port map( -- 
              preds => ptr_deref_110_trigger_x_x411_predecessors,
              symbol_out => ptr_deref_110_trigger_x_x411_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_trigger_
        ptr_deref_110_active_x_x412_symbol <= ptr_deref_110_request_459_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_active_
        ptr_deref_110_base_address_calculated_413_symbol <= simple_obj_ref_109_complete_414_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_address_calculated
        simple_obj_ref_109_complete_414_symbol <= assign_stmt_108_completed_x_x384_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_109_complete
        ptr_deref_110_root_address_calculated_415_symbol <= ptr_deref_110_base_plus_offset_423_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_root_address_calculated
        ptr_deref_110_word_address_calculated_416_symbol <= ptr_deref_110_word_addrgen_428_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_address_calculated
        ptr_deref_110_base_address_resized_417_symbol <= ptr_deref_110_base_addr_resize_418_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_address_resized
        ptr_deref_110_base_addr_resize_418: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize 
          signal ptr_deref_110_base_addr_resize_418_start: Boolean;
          signal Xentry_419_symbol: Boolean;
          signal Xexit_420_symbol: Boolean;
          signal base_resize_req_421_symbol : Boolean;
          signal base_resize_ack_422_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_base_addr_resize_418_start <= ptr_deref_110_base_address_calculated_413_symbol; -- control passed to block
          Xentry_419_symbol  <= ptr_deref_110_base_addr_resize_418_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/$entry
          base_resize_req_421_symbol <= Xentry_419_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/base_resize_req
          ptr_deref_110_base_resize_req_0 <= base_resize_req_421_symbol; -- link to DP
          base_resize_ack_422_symbol <= ptr_deref_110_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/base_resize_ack
          Xexit_420_symbol <= base_resize_ack_422_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/$exit
          ptr_deref_110_base_addr_resize_418_symbol <= Xexit_420_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize
        ptr_deref_110_base_plus_offset_423: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset 
          signal ptr_deref_110_base_plus_offset_423_start: Boolean;
          signal Xentry_424_symbol: Boolean;
          signal Xexit_425_symbol: Boolean;
          signal sum_rename_req_426_symbol : Boolean;
          signal sum_rename_ack_427_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_base_plus_offset_423_start <= ptr_deref_110_base_address_resized_417_symbol; -- control passed to block
          Xentry_424_symbol  <= ptr_deref_110_base_plus_offset_423_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/$entry
          sum_rename_req_426_symbol <= Xentry_424_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/sum_rename_req
          ptr_deref_110_root_address_inst_req_0 <= sum_rename_req_426_symbol; -- link to DP
          sum_rename_ack_427_symbol <= ptr_deref_110_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/sum_rename_ack
          Xexit_425_symbol <= sum_rename_ack_427_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/$exit
          ptr_deref_110_base_plus_offset_423_symbol <= Xexit_425_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset
        ptr_deref_110_word_addrgen_428: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen 
          signal ptr_deref_110_word_addrgen_428_start: Boolean;
          signal Xentry_429_symbol: Boolean;
          signal Xexit_430_symbol: Boolean;
          signal word_0_431_symbol : Boolean;
          signal word_1_438_symbol : Boolean;
          signal word_2_445_symbol : Boolean;
          signal word_3_452_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_word_addrgen_428_start <= ptr_deref_110_root_address_calculated_415_symbol; -- control passed to block
          Xentry_429_symbol  <= ptr_deref_110_word_addrgen_428_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/$entry
          word_0_431: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0 
            signal word_0_431_start: Boolean;
            signal Xentry_432_symbol: Boolean;
            signal Xexit_433_symbol: Boolean;
            signal rr_434_symbol : Boolean;
            signal ra_435_symbol : Boolean;
            signal cr_436_symbol : Boolean;
            signal ca_437_symbol : Boolean;
            -- 
          begin -- 
            word_0_431_start <= Xentry_429_symbol; -- control passed to block
            Xentry_432_symbol  <= word_0_431_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0/$entry
            rr_434_symbol <= Xentry_432_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0/rr
            ptr_deref_110_addr_0_req_0 <= rr_434_symbol; -- link to DP
            ra_435_symbol <= ptr_deref_110_addr_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0/ra
            cr_436_symbol <= ra_435_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0/cr
            ptr_deref_110_addr_0_req_1 <= cr_436_symbol; -- link to DP
            ca_437_symbol <= ptr_deref_110_addr_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0/ca
            Xexit_433_symbol <= ca_437_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0/$exit
            word_0_431_symbol <= Xexit_433_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_0
          word_1_438: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1 
            signal word_1_438_start: Boolean;
            signal Xentry_439_symbol: Boolean;
            signal Xexit_440_symbol: Boolean;
            signal rr_441_symbol : Boolean;
            signal ra_442_symbol : Boolean;
            signal cr_443_symbol : Boolean;
            signal ca_444_symbol : Boolean;
            -- 
          begin -- 
            word_1_438_start <= Xentry_429_symbol; -- control passed to block
            Xentry_439_symbol  <= word_1_438_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1/$entry
            rr_441_symbol <= Xentry_439_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1/rr
            ptr_deref_110_addr_1_req_0 <= rr_441_symbol; -- link to DP
            ra_442_symbol <= ptr_deref_110_addr_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1/ra
            cr_443_symbol <= ra_442_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1/cr
            ptr_deref_110_addr_1_req_1 <= cr_443_symbol; -- link to DP
            ca_444_symbol <= ptr_deref_110_addr_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1/ca
            Xexit_440_symbol <= ca_444_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1/$exit
            word_1_438_symbol <= Xexit_440_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_1
          word_2_445: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2 
            signal word_2_445_start: Boolean;
            signal Xentry_446_symbol: Boolean;
            signal Xexit_447_symbol: Boolean;
            signal rr_448_symbol : Boolean;
            signal ra_449_symbol : Boolean;
            signal cr_450_symbol : Boolean;
            signal ca_451_symbol : Boolean;
            -- 
          begin -- 
            word_2_445_start <= Xentry_429_symbol; -- control passed to block
            Xentry_446_symbol  <= word_2_445_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2/$entry
            rr_448_symbol <= Xentry_446_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2/rr
            ptr_deref_110_addr_2_req_0 <= rr_448_symbol; -- link to DP
            ra_449_symbol <= ptr_deref_110_addr_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2/ra
            cr_450_symbol <= ra_449_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2/cr
            ptr_deref_110_addr_2_req_1 <= cr_450_symbol; -- link to DP
            ca_451_symbol <= ptr_deref_110_addr_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2/ca
            Xexit_447_symbol <= ca_451_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2/$exit
            word_2_445_symbol <= Xexit_447_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_2
          word_3_452: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3 
            signal word_3_452_start: Boolean;
            signal Xentry_453_symbol: Boolean;
            signal Xexit_454_symbol: Boolean;
            signal rr_455_symbol : Boolean;
            signal ra_456_symbol : Boolean;
            signal cr_457_symbol : Boolean;
            signal ca_458_symbol : Boolean;
            -- 
          begin -- 
            word_3_452_start <= Xentry_429_symbol; -- control passed to block
            Xentry_453_symbol  <= word_3_452_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3/$entry
            rr_455_symbol <= Xentry_453_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3/rr
            ptr_deref_110_addr_3_req_0 <= rr_455_symbol; -- link to DP
            ra_456_symbol <= ptr_deref_110_addr_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3/ra
            cr_457_symbol <= ra_456_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3/cr
            ptr_deref_110_addr_3_req_1 <= cr_457_symbol; -- link to DP
            ca_458_symbol <= ptr_deref_110_addr_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3/ca
            Xexit_454_symbol <= ca_458_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3/$exit
            word_3_452_symbol <= Xexit_454_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/word_3
          Xexit_430_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/$exit 
            signal Xexit_430_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_430_predecessors(0) <= word_0_431_symbol;
            Xexit_430_predecessors(1) <= word_1_438_symbol;
            Xexit_430_predecessors(2) <= word_2_445_symbol;
            Xexit_430_predecessors(3) <= word_3_452_symbol;
            Xexit_430_join: join -- 
              port map( -- 
                preds => Xexit_430_predecessors,
                symbol_out => Xexit_430_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/$exit
          ptr_deref_110_word_addrgen_428_symbol <= Xexit_430_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen
        ptr_deref_110_request_459: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request 
          signal ptr_deref_110_request_459_start: Boolean;
          signal Xentry_460_symbol: Boolean;
          signal Xexit_461_symbol: Boolean;
          signal split_req_462_symbol : Boolean;
          signal split_ack_463_symbol : Boolean;
          signal word_access_464_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_request_459_start <= ptr_deref_110_trigger_x_x411_symbol; -- control passed to block
          Xentry_460_symbol  <= ptr_deref_110_request_459_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/$entry
          split_req_462_symbol <= Xentry_460_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/split_req
          ptr_deref_110_gather_scatter_req_0 <= split_req_462_symbol; -- link to DP
          split_ack_463_symbol <= ptr_deref_110_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/split_ack
          word_access_464: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access 
            signal word_access_464_start: Boolean;
            signal Xentry_465_symbol: Boolean;
            signal Xexit_466_symbol: Boolean;
            signal word_access_0_467_symbol : Boolean;
            signal word_access_1_472_symbol : Boolean;
            signal word_access_2_477_symbol : Boolean;
            signal word_access_3_482_symbol : Boolean;
            -- 
          begin -- 
            word_access_464_start <= split_ack_463_symbol; -- control passed to block
            Xentry_465_symbol  <= word_access_464_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/$entry
            word_access_0_467: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0 
              signal word_access_0_467_start: Boolean;
              signal Xentry_468_symbol: Boolean;
              signal Xexit_469_symbol: Boolean;
              signal rr_470_symbol : Boolean;
              signal ra_471_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_467_start <= Xentry_465_symbol; -- control passed to block
              Xentry_468_symbol  <= word_access_0_467_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/$entry
              rr_470_symbol <= Xentry_468_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/rr
              ptr_deref_110_store_0_req_0 <= rr_470_symbol; -- link to DP
              ra_471_symbol <= ptr_deref_110_store_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/ra
              Xexit_469_symbol <= ra_471_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/$exit
              word_access_0_467_symbol <= Xexit_469_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0
            word_access_1_472: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_1 
              signal word_access_1_472_start: Boolean;
              signal Xentry_473_symbol: Boolean;
              signal Xexit_474_symbol: Boolean;
              signal rr_475_symbol : Boolean;
              signal ra_476_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_472_start <= Xentry_465_symbol; -- control passed to block
              Xentry_473_symbol  <= word_access_1_472_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_1/$entry
              rr_475_symbol <= Xentry_473_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_1/rr
              ptr_deref_110_store_1_req_0 <= rr_475_symbol; -- link to DP
              ra_476_symbol <= ptr_deref_110_store_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_1/ra
              Xexit_474_symbol <= ra_476_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_1/$exit
              word_access_1_472_symbol <= Xexit_474_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_1
            word_access_2_477: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_2 
              signal word_access_2_477_start: Boolean;
              signal Xentry_478_symbol: Boolean;
              signal Xexit_479_symbol: Boolean;
              signal rr_480_symbol : Boolean;
              signal ra_481_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_477_start <= Xentry_465_symbol; -- control passed to block
              Xentry_478_symbol  <= word_access_2_477_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_2/$entry
              rr_480_symbol <= Xentry_478_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_2/rr
              ptr_deref_110_store_2_req_0 <= rr_480_symbol; -- link to DP
              ra_481_symbol <= ptr_deref_110_store_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_2/ra
              Xexit_479_symbol <= ra_481_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_2/$exit
              word_access_2_477_symbol <= Xexit_479_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_2
            word_access_3_482: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_3 
              signal word_access_3_482_start: Boolean;
              signal Xentry_483_symbol: Boolean;
              signal Xexit_484_symbol: Boolean;
              signal rr_485_symbol : Boolean;
              signal ra_486_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_482_start <= Xentry_465_symbol; -- control passed to block
              Xentry_483_symbol  <= word_access_3_482_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_3/$entry
              rr_485_symbol <= Xentry_483_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_3/rr
              ptr_deref_110_store_3_req_0 <= rr_485_symbol; -- link to DP
              ra_486_symbol <= ptr_deref_110_store_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_3/ra
              Xexit_484_symbol <= ra_486_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_3/$exit
              word_access_3_482_symbol <= Xexit_484_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_3
            Xexit_466_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/$exit 
              signal Xexit_466_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_466_predecessors(0) <= word_access_0_467_symbol;
              Xexit_466_predecessors(1) <= word_access_1_472_symbol;
              Xexit_466_predecessors(2) <= word_access_2_477_symbol;
              Xexit_466_predecessors(3) <= word_access_3_482_symbol;
              Xexit_466_join: join -- 
                port map( -- 
                  preds => Xexit_466_predecessors,
                  symbol_out => Xexit_466_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/$exit
            word_access_464_symbol <= Xexit_466_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access
          Xexit_461_symbol <= word_access_464_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/$exit
          ptr_deref_110_request_459_symbol <= Xexit_461_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request
        ptr_deref_110_complete_487: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete 
          signal ptr_deref_110_complete_487_start: Boolean;
          signal Xentry_488_symbol: Boolean;
          signal Xexit_489_symbol: Boolean;
          signal word_access_490_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_complete_487_start <= ptr_deref_110_active_x_x412_symbol; -- control passed to block
          Xentry_488_symbol  <= ptr_deref_110_complete_487_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/$entry
          word_access_490: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access 
            signal word_access_490_start: Boolean;
            signal Xentry_491_symbol: Boolean;
            signal Xexit_492_symbol: Boolean;
            signal word_access_0_493_symbol : Boolean;
            signal word_access_1_498_symbol : Boolean;
            signal word_access_2_503_symbol : Boolean;
            signal word_access_3_508_symbol : Boolean;
            -- 
          begin -- 
            word_access_490_start <= Xentry_488_symbol; -- control passed to block
            Xentry_491_symbol  <= word_access_490_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/$entry
            word_access_0_493: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0 
              signal word_access_0_493_start: Boolean;
              signal Xentry_494_symbol: Boolean;
              signal Xexit_495_symbol: Boolean;
              signal cr_496_symbol : Boolean;
              signal ca_497_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_493_start <= Xentry_491_symbol; -- control passed to block
              Xentry_494_symbol  <= word_access_0_493_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/$entry
              cr_496_symbol <= Xentry_494_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/cr
              ptr_deref_110_store_0_req_1 <= cr_496_symbol; -- link to DP
              ca_497_symbol <= ptr_deref_110_store_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/ca
              Xexit_495_symbol <= ca_497_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/$exit
              word_access_0_493_symbol <= Xexit_495_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0
            word_access_1_498: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_1 
              signal word_access_1_498_start: Boolean;
              signal Xentry_499_symbol: Boolean;
              signal Xexit_500_symbol: Boolean;
              signal cr_501_symbol : Boolean;
              signal ca_502_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_498_start <= Xentry_491_symbol; -- control passed to block
              Xentry_499_symbol  <= word_access_1_498_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_1/$entry
              cr_501_symbol <= Xentry_499_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_1/cr
              ptr_deref_110_store_1_req_1 <= cr_501_symbol; -- link to DP
              ca_502_symbol <= ptr_deref_110_store_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_1/ca
              Xexit_500_symbol <= ca_502_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_1/$exit
              word_access_1_498_symbol <= Xexit_500_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_1
            word_access_2_503: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_2 
              signal word_access_2_503_start: Boolean;
              signal Xentry_504_symbol: Boolean;
              signal Xexit_505_symbol: Boolean;
              signal cr_506_symbol : Boolean;
              signal ca_507_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_503_start <= Xentry_491_symbol; -- control passed to block
              Xentry_504_symbol  <= word_access_2_503_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_2/$entry
              cr_506_symbol <= Xentry_504_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_2/cr
              ptr_deref_110_store_2_req_1 <= cr_506_symbol; -- link to DP
              ca_507_symbol <= ptr_deref_110_store_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_2/ca
              Xexit_505_symbol <= ca_507_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_2/$exit
              word_access_2_503_symbol <= Xexit_505_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_2
            word_access_3_508: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_3 
              signal word_access_3_508_start: Boolean;
              signal Xentry_509_symbol: Boolean;
              signal Xexit_510_symbol: Boolean;
              signal cr_511_symbol : Boolean;
              signal ca_512_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_508_start <= Xentry_491_symbol; -- control passed to block
              Xentry_509_symbol  <= word_access_3_508_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_3/$entry
              cr_511_symbol <= Xentry_509_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_3/cr
              ptr_deref_110_store_3_req_1 <= cr_511_symbol; -- link to DP
              ca_512_symbol <= ptr_deref_110_store_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_3/ca
              Xexit_510_symbol <= ca_512_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_3/$exit
              word_access_3_508_symbol <= Xexit_510_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_3
            Xexit_492_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/$exit 
              signal Xexit_492_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_492_predecessors(0) <= word_access_0_493_symbol;
              Xexit_492_predecessors(1) <= word_access_1_498_symbol;
              Xexit_492_predecessors(2) <= word_access_2_503_symbol;
              Xexit_492_predecessors(3) <= word_access_3_508_symbol;
              Xexit_492_join: join -- 
                port map( -- 
                  preds => Xexit_492_predecessors,
                  symbol_out => Xexit_492_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/$exit
            word_access_490_symbol <= Xexit_492_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access
          Xexit_489_symbol <= word_access_490_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/$exit
          ptr_deref_110_complete_487_symbol <= Xexit_489_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete
        assign_stmt_116_active_x_x513_symbol <= ptr_deref_115_complete_546_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_116_active_
        assign_stmt_116_completed_x_x514_symbol <= assign_stmt_116_active_x_x513_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_116_completed_
        ptr_deref_115_trigger_x_x515_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_trigger_ 
          signal ptr_deref_115_trigger_x_x515_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_115_trigger_x_x515_predecessors(0) <= ptr_deref_115_word_address_calculated_519_symbol;
          ptr_deref_115_trigger_x_x515_predecessors(1) <= ptr_deref_110_active_x_x412_symbol;
          ptr_deref_115_trigger_x_x515_join: join -- 
            port map( -- 
              preds => ptr_deref_115_trigger_x_x515_predecessors,
              symbol_out => ptr_deref_115_trigger_x_x515_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_trigger_
        ptr_deref_115_active_x_x516_symbol <= ptr_deref_115_request_520_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_active_
        ptr_deref_115_base_address_calculated_517_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_base_address_calculated
        ptr_deref_115_root_address_calculated_518_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_root_address_calculated
        ptr_deref_115_word_address_calculated_519_symbol <= ptr_deref_115_root_address_calculated_518_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_word_address_calculated
        ptr_deref_115_request_520: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request 
          signal ptr_deref_115_request_520_start: Boolean;
          signal Xentry_521_symbol: Boolean;
          signal Xexit_522_symbol: Boolean;
          signal word_access_523_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_115_request_520_start <= ptr_deref_115_trigger_x_x515_symbol; -- control passed to block
          Xentry_521_symbol  <= ptr_deref_115_request_520_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/$entry
          word_access_523: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access 
            signal word_access_523_start: Boolean;
            signal Xentry_524_symbol: Boolean;
            signal Xexit_525_symbol: Boolean;
            signal word_access_0_526_symbol : Boolean;
            signal word_access_1_531_symbol : Boolean;
            signal word_access_2_536_symbol : Boolean;
            signal word_access_3_541_symbol : Boolean;
            -- 
          begin -- 
            word_access_523_start <= Xentry_521_symbol; -- control passed to block
            Xentry_524_symbol  <= word_access_523_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/$entry
            word_access_0_526: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0 
              signal word_access_0_526_start: Boolean;
              signal Xentry_527_symbol: Boolean;
              signal Xexit_528_symbol: Boolean;
              signal rr_529_symbol : Boolean;
              signal ra_530_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_526_start <= Xentry_524_symbol; -- control passed to block
              Xentry_527_symbol  <= word_access_0_526_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/$entry
              rr_529_symbol <= Xentry_527_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/rr
              ptr_deref_115_load_0_req_0 <= rr_529_symbol; -- link to DP
              ra_530_symbol <= ptr_deref_115_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/ra
              Xexit_528_symbol <= ra_530_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/$exit
              word_access_0_526_symbol <= Xexit_528_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0
            word_access_1_531: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_1 
              signal word_access_1_531_start: Boolean;
              signal Xentry_532_symbol: Boolean;
              signal Xexit_533_symbol: Boolean;
              signal rr_534_symbol : Boolean;
              signal ra_535_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_531_start <= Xentry_524_symbol; -- control passed to block
              Xentry_532_symbol  <= word_access_1_531_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_1/$entry
              rr_534_symbol <= Xentry_532_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_1/rr
              ptr_deref_115_load_1_req_0 <= rr_534_symbol; -- link to DP
              ra_535_symbol <= ptr_deref_115_load_1_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_1/ra
              Xexit_533_symbol <= ra_535_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_1/$exit
              word_access_1_531_symbol <= Xexit_533_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_1
            word_access_2_536: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_2 
              signal word_access_2_536_start: Boolean;
              signal Xentry_537_symbol: Boolean;
              signal Xexit_538_symbol: Boolean;
              signal rr_539_symbol : Boolean;
              signal ra_540_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_536_start <= Xentry_524_symbol; -- control passed to block
              Xentry_537_symbol  <= word_access_2_536_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_2/$entry
              rr_539_symbol <= Xentry_537_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_2/rr
              ptr_deref_115_load_2_req_0 <= rr_539_symbol; -- link to DP
              ra_540_symbol <= ptr_deref_115_load_2_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_2/ra
              Xexit_538_symbol <= ra_540_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_2/$exit
              word_access_2_536_symbol <= Xexit_538_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_2
            word_access_3_541: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_3 
              signal word_access_3_541_start: Boolean;
              signal Xentry_542_symbol: Boolean;
              signal Xexit_543_symbol: Boolean;
              signal rr_544_symbol : Boolean;
              signal ra_545_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_541_start <= Xentry_524_symbol; -- control passed to block
              Xentry_542_symbol  <= word_access_3_541_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_3/$entry
              rr_544_symbol <= Xentry_542_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_3/rr
              ptr_deref_115_load_3_req_0 <= rr_544_symbol; -- link to DP
              ra_545_symbol <= ptr_deref_115_load_3_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_3/ra
              Xexit_543_symbol <= ra_545_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_3/$exit
              word_access_3_541_symbol <= Xexit_543_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_3
            Xexit_525_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/$exit 
              signal Xexit_525_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_525_predecessors(0) <= word_access_0_526_symbol;
              Xexit_525_predecessors(1) <= word_access_1_531_symbol;
              Xexit_525_predecessors(2) <= word_access_2_536_symbol;
              Xexit_525_predecessors(3) <= word_access_3_541_symbol;
              Xexit_525_join: join -- 
                port map( -- 
                  preds => Xexit_525_predecessors,
                  symbol_out => Xexit_525_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/$exit
            word_access_523_symbol <= Xexit_525_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access
          Xexit_522_symbol <= word_access_523_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/$exit
          ptr_deref_115_request_520_symbol <= Xexit_522_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request
        ptr_deref_115_complete_546: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete 
          signal ptr_deref_115_complete_546_start: Boolean;
          signal Xentry_547_symbol: Boolean;
          signal Xexit_548_symbol: Boolean;
          signal word_access_549_symbol : Boolean;
          signal merge_req_572_symbol : Boolean;
          signal merge_ack_573_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_115_complete_546_start <= ptr_deref_115_active_x_x516_symbol; -- control passed to block
          Xentry_547_symbol  <= ptr_deref_115_complete_546_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/$entry
          word_access_549: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access 
            signal word_access_549_start: Boolean;
            signal Xentry_550_symbol: Boolean;
            signal Xexit_551_symbol: Boolean;
            signal word_access_0_552_symbol : Boolean;
            signal word_access_1_557_symbol : Boolean;
            signal word_access_2_562_symbol : Boolean;
            signal word_access_3_567_symbol : Boolean;
            -- 
          begin -- 
            word_access_549_start <= Xentry_547_symbol; -- control passed to block
            Xentry_550_symbol  <= word_access_549_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/$entry
            word_access_0_552: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0 
              signal word_access_0_552_start: Boolean;
              signal Xentry_553_symbol: Boolean;
              signal Xexit_554_symbol: Boolean;
              signal cr_555_symbol : Boolean;
              signal ca_556_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_552_start <= Xentry_550_symbol; -- control passed to block
              Xentry_553_symbol  <= word_access_0_552_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/$entry
              cr_555_symbol <= Xentry_553_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/cr
              ptr_deref_115_load_0_req_1 <= cr_555_symbol; -- link to DP
              ca_556_symbol <= ptr_deref_115_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/ca
              Xexit_554_symbol <= ca_556_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/$exit
              word_access_0_552_symbol <= Xexit_554_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0
            word_access_1_557: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_1 
              signal word_access_1_557_start: Boolean;
              signal Xentry_558_symbol: Boolean;
              signal Xexit_559_symbol: Boolean;
              signal cr_560_symbol : Boolean;
              signal ca_561_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_557_start <= Xentry_550_symbol; -- control passed to block
              Xentry_558_symbol  <= word_access_1_557_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_1/$entry
              cr_560_symbol <= Xentry_558_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_1/cr
              ptr_deref_115_load_1_req_1 <= cr_560_symbol; -- link to DP
              ca_561_symbol <= ptr_deref_115_load_1_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_1/ca
              Xexit_559_symbol <= ca_561_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_1/$exit
              word_access_1_557_symbol <= Xexit_559_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_1
            word_access_2_562: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_2 
              signal word_access_2_562_start: Boolean;
              signal Xentry_563_symbol: Boolean;
              signal Xexit_564_symbol: Boolean;
              signal cr_565_symbol : Boolean;
              signal ca_566_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_562_start <= Xentry_550_symbol; -- control passed to block
              Xentry_563_symbol  <= word_access_2_562_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_2/$entry
              cr_565_symbol <= Xentry_563_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_2/cr
              ptr_deref_115_load_2_req_1 <= cr_565_symbol; -- link to DP
              ca_566_symbol <= ptr_deref_115_load_2_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_2/ca
              Xexit_564_symbol <= ca_566_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_2/$exit
              word_access_2_562_symbol <= Xexit_564_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_2
            word_access_3_567: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_3 
              signal word_access_3_567_start: Boolean;
              signal Xentry_568_symbol: Boolean;
              signal Xexit_569_symbol: Boolean;
              signal cr_570_symbol : Boolean;
              signal ca_571_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_567_start <= Xentry_550_symbol; -- control passed to block
              Xentry_568_symbol  <= word_access_3_567_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_3/$entry
              cr_570_symbol <= Xentry_568_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_3/cr
              ptr_deref_115_load_3_req_1 <= cr_570_symbol; -- link to DP
              ca_571_symbol <= ptr_deref_115_load_3_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_3/ca
              Xexit_569_symbol <= ca_571_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_3/$exit
              word_access_3_567_symbol <= Xexit_569_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_3
            Xexit_551_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/$exit 
              signal Xexit_551_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_551_predecessors(0) <= word_access_0_552_symbol;
              Xexit_551_predecessors(1) <= word_access_1_557_symbol;
              Xexit_551_predecessors(2) <= word_access_2_562_symbol;
              Xexit_551_predecessors(3) <= word_access_3_567_symbol;
              Xexit_551_join: join -- 
                port map( -- 
                  preds => Xexit_551_predecessors,
                  symbol_out => Xexit_551_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/$exit
            word_access_549_symbol <= Xexit_551_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access
          merge_req_572_symbol <= word_access_549_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/merge_req
          ptr_deref_115_gather_scatter_req_0 <= merge_req_572_symbol; -- link to DP
          merge_ack_573_symbol <= ptr_deref_115_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/merge_ack
          Xexit_548_symbol <= merge_ack_573_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/$exit
          ptr_deref_115_complete_546_symbol <= Xexit_548_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete
        assign_stmt_120_active_x_x574_symbol <= type_cast_119_complete_579_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_120_active_
        assign_stmt_120_completed_x_x575_symbol <= assign_stmt_120_active_x_x574_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_120_completed_
        type_cast_119_active_x_x576_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_active_ 
          signal type_cast_119_active_x_x576_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_119_active_x_x576_predecessors(0) <= type_cast_119_trigger_x_x577_symbol;
          type_cast_119_active_x_x576_predecessors(1) <= simple_obj_ref_118_complete_578_symbol;
          type_cast_119_active_x_x576_join: join -- 
            port map( -- 
              preds => type_cast_119_active_x_x576_predecessors,
              symbol_out => type_cast_119_active_x_x576_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_active_
        type_cast_119_trigger_x_x577_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_trigger_
        simple_obj_ref_118_complete_578_symbol <= assign_stmt_116_completed_x_x514_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_118_complete
        type_cast_119_complete_579: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete 
          signal type_cast_119_complete_579_start: Boolean;
          signal Xentry_580_symbol: Boolean;
          signal Xexit_581_symbol: Boolean;
          signal req_582_symbol : Boolean;
          signal ack_583_symbol : Boolean;
          -- 
        begin -- 
          type_cast_119_complete_579_start <= type_cast_119_active_x_x576_symbol; -- control passed to block
          Xentry_580_symbol  <= type_cast_119_complete_579_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/$entry
          req_582_symbol <= Xentry_580_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/req
          type_cast_119_inst_req_0 <= req_582_symbol; -- link to DP
          ack_583_symbol <= type_cast_119_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/ack
          Xexit_581_symbol <= ack_583_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/$exit
          type_cast_119_complete_579_symbol <= Xexit_581_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete
        Xexit_47_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/$exit 
          signal Xexit_47_predecessors: BooleanArray(6 downto 0);
          -- 
        begin -- 
          Xexit_47_predecessors(0) <= assign_stmt_81_completed_x_x59_symbol;
          Xexit_47_predecessors(1) <= ptr_deref_79_base_address_calculated_63_symbol;
          Xexit_47_predecessors(2) <= ptr_deref_84_base_address_calculated_124_symbol;
          Xexit_47_predecessors(3) <= ptr_deref_102_base_address_calculated_326_symbol;
          Xexit_47_predecessors(4) <= assign_stmt_112_completed_x_x409_symbol;
          Xexit_47_predecessors(5) <= ptr_deref_115_base_address_calculated_517_symbol;
          Xexit_47_predecessors(6) <= assign_stmt_120_completed_x_x575_symbol;
          Xexit_47_join: join -- 
            port map( -- 
              preds => Xexit_47_predecessors,
              symbol_out => Xexit_47_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/$exit
        assign_stmt_77_to_assign_stmt_125_45_symbol <= Xexit_47_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125
      assign_stmt_129_584: Block -- branch_block_stmt_56/assign_stmt_129 
        signal assign_stmt_129_584_start: Boolean;
        signal Xentry_585_symbol: Boolean;
        signal Xexit_586_symbol: Boolean;
        signal assign_stmt_129_active_x_x587_symbol : Boolean;
        signal assign_stmt_129_completed_x_x588_symbol : Boolean;
        signal type_cast_128_active_x_x589_symbol : Boolean;
        signal type_cast_128_trigger_x_x590_symbol : Boolean;
        signal simple_obj_ref_127_complete_591_symbol : Boolean;
        signal type_cast_128_complete_592_symbol : Boolean;
        signal simple_obj_ref_126_trigger_x_x597_symbol : Boolean;
        signal simple_obj_ref_126_complete_598_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_129_584_start <= assign_stmt_129_x_xentry_x_xx_x18_symbol; -- control passed to block
        Xentry_585_symbol  <= assign_stmt_129_584_start; -- transition branch_block_stmt_56/assign_stmt_129/$entry
        assign_stmt_129_active_x_x587_symbol <= type_cast_128_complete_592_symbol; -- transition branch_block_stmt_56/assign_stmt_129/assign_stmt_129_active_
        assign_stmt_129_completed_x_x588_symbol <= simple_obj_ref_126_complete_598_symbol; -- transition branch_block_stmt_56/assign_stmt_129/assign_stmt_129_completed_
        type_cast_128_active_x_x589_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_129/type_cast_128_active_ 
          signal type_cast_128_active_x_x589_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_128_active_x_x589_predecessors(0) <= type_cast_128_trigger_x_x590_symbol;
          type_cast_128_active_x_x589_predecessors(1) <= simple_obj_ref_127_complete_591_symbol;
          type_cast_128_active_x_x589_join: join -- 
            port map( -- 
              preds => type_cast_128_active_x_x589_predecessors,
              symbol_out => type_cast_128_active_x_x589_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_129/type_cast_128_active_
        type_cast_128_trigger_x_x590_symbol <= Xentry_585_symbol; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_trigger_
        simple_obj_ref_127_complete_591_symbol <= Xentry_585_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_127_complete
        type_cast_128_complete_592: Block -- branch_block_stmt_56/assign_stmt_129/type_cast_128_complete 
          signal type_cast_128_complete_592_start: Boolean;
          signal Xentry_593_symbol: Boolean;
          signal Xexit_594_symbol: Boolean;
          signal req_595_symbol : Boolean;
          signal ack_596_symbol : Boolean;
          -- 
        begin -- 
          type_cast_128_complete_592_start <= type_cast_128_active_x_x589_symbol; -- control passed to block
          Xentry_593_symbol  <= type_cast_128_complete_592_start; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/$entry
          req_595_symbol <= Xentry_593_symbol; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/req
          type_cast_128_inst_req_0 <= req_595_symbol; -- link to DP
          ack_596_symbol <= type_cast_128_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/ack
          Xexit_594_symbol <= ack_596_symbol; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/$exit
          type_cast_128_complete_592_symbol <= Xexit_594_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_129/type_cast_128_complete
        simple_obj_ref_126_trigger_x_x597_symbol <= assign_stmt_129_active_x_x587_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_trigger_
        simple_obj_ref_126_complete_598: Block -- branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete 
          signal simple_obj_ref_126_complete_598_start: Boolean;
          signal Xentry_599_symbol: Boolean;
          signal Xexit_600_symbol: Boolean;
          signal pipe_wreq_601_symbol : Boolean;
          signal pipe_wack_602_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_126_complete_598_start <= simple_obj_ref_126_trigger_x_x597_symbol; -- control passed to block
          Xentry_599_symbol  <= simple_obj_ref_126_complete_598_start; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/$entry
          pipe_wreq_601_symbol <= Xentry_599_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/pipe_wreq
          simple_obj_ref_126_inst_req_0 <= pipe_wreq_601_symbol; -- link to DP
          pipe_wack_602_symbol <= simple_obj_ref_126_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/pipe_wack
          Xexit_600_symbol <= pipe_wack_602_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/$exit
          simple_obj_ref_126_complete_598_symbol <= Xexit_600_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete
        Xexit_586_symbol <= assign_stmt_129_completed_x_x588_symbol; -- transition branch_block_stmt_56/assign_stmt_129/$exit
        assign_stmt_129_584_symbol <= Xexit_586_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_129
      bb_0_bb_1_PhiReq_603: Block -- branch_block_stmt_56/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_603_start: Boolean;
        signal Xentry_604_symbol: Boolean;
        signal Xexit_605_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_603_start <= bb_0_bb_1_10_symbol; -- control passed to block
        Xentry_604_symbol  <= bb_0_bb_1_PhiReq_603_start; -- transition branch_block_stmt_56/bb_0_bb_1_PhiReq/$entry
        Xexit_605_symbol <= Xentry_604_symbol; -- transition branch_block_stmt_56/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_603_symbol <= Xexit_605_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/bb_0_bb_1_PhiReq
      bb_1_bb_1_PhiReq_606: Block -- branch_block_stmt_56/bb_1_bb_1_PhiReq 
        signal bb_1_bb_1_PhiReq_606_start: Boolean;
        signal Xentry_607_symbol: Boolean;
        signal Xexit_608_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_1_PhiReq_606_start <= bb_1_bb_1_20_symbol; -- control passed to block
        Xentry_607_symbol  <= bb_1_bb_1_PhiReq_606_start; -- transition branch_block_stmt_56/bb_1_bb_1_PhiReq/$entry
        Xexit_608_symbol <= Xentry_607_symbol; -- transition branch_block_stmt_56/bb_1_bb_1_PhiReq/$exit
        bb_1_bb_1_PhiReq_606_symbol <= Xexit_608_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/bb_1_bb_1_PhiReq
      merge_stmt_63_PhiReqMerge_609_symbol  <=  bb_0_bb_1_PhiReq_603_symbol or bb_1_bb_1_PhiReq_606_symbol; -- place branch_block_stmt_56/merge_stmt_63_PhiReqMerge (optimized away) 
      merge_stmt_63_PhiAck_610: Block -- branch_block_stmt_56/merge_stmt_63_PhiAck 
        signal merge_stmt_63_PhiAck_610_start: Boolean;
        signal Xentry_611_symbol: Boolean;
        signal Xexit_612_symbol: Boolean;
        signal dummy_613_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_63_PhiAck_610_start <= merge_stmt_63_PhiReqMerge_609_symbol; -- control passed to block
        Xentry_611_symbol  <= merge_stmt_63_PhiAck_610_start; -- transition branch_block_stmt_56/merge_stmt_63_PhiAck/$entry
        dummy_613_symbol <= Xentry_611_symbol; -- transition branch_block_stmt_56/merge_stmt_63_PhiAck/dummy
        Xexit_612_symbol <= dummy_613_symbol; -- transition branch_block_stmt_56/merge_stmt_63_PhiAck/$exit
        merge_stmt_63_PhiAck_610_symbol <= Xexit_612_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/merge_stmt_63_PhiAck
      Xexit_5_symbol <= branch_block_stmt_56_x_xexit_x_xx_x7_symbol; -- transition branch_block_stmt_56/$exit
      branch_block_stmt_56_3_symbol <= Xexit_5_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_56
    Xexit_2_symbol <= branch_block_stmt_56_3_symbol; -- transition $exit
    fin  <=  '1' when Xexit_2_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_107_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_107_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_107_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_89_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_89_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_89_root_address : std_logic_vector(5 downto 0);
    signal expr_96_wire_constant : std_logic_vector(31 downto 0);
    signal iNsTr_10_108 : std_logic_vector(31 downto 0);
    signal iNsTr_12_116 : std_logic_vector(31 downto 0);
    signal iNsTr_13_120 : std_logic_vector(31 downto 0);
    signal iNsTr_14_125 : std_logic_vector(31 downto 0);
    signal iNsTr_1_68 : std_logic_vector(31 downto 0);
    signal iNsTr_2_73 : std_logic_vector(31 downto 0);
    signal iNsTr_3_77 : std_logic_vector(31 downto 0);
    signal iNsTr_5_85 : std_logic_vector(31 downto 0);
    signal iNsTr_6_90 : std_logic_vector(31 downto 0);
    signal iNsTr_7_94 : std_logic_vector(31 downto 0);
    signal iNsTr_8_99 : std_logic_vector(31 downto 0);
    signal iNsTr_9_103 : std_logic_vector(31 downto 0);
    signal lptr_61 : std_logic_vector(31 downto 0);
    signal ptr_deref_102_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_102_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_102_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_102_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_102_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_102_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_102_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_102_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_110_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_110_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_110_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_110_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_110_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_110_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_110_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_110_word_offset_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_115_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_115_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_115_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_115_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_115_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_115_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_115_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_115_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_79_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_79_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_79_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_79_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_79_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_79_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_79_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_79_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_79_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_84_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_84_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_84_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_84_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_84_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_84_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_84_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_84_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_93_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_93_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_93_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_93_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_93_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_93_word_offset_3 : std_logic_vector(5 downto 0);
    signal simple_obj_ref_71_wire : std_logic_vector(31 downto 0);
    signal type_cast_128_wire : std_logic_vector(31 downto 0);
    signal xxfooxxbodyxxlptr_alloc_base_address : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    array_obj_ref_107_final_offset <= "000100";
    array_obj_ref_89_final_offset <= "000100";
    expr_96_wire_constant <= "00000000000000000000000000000010";
    iNsTr_14_125 <= "00000000000000000000000000000000";
    iNsTr_1_68 <= "00000000000000000000000000000000";
    lptr_61 <= "00000000000000000000000000011000";
    ptr_deref_102_word_address_0 <= "011000";
    ptr_deref_102_word_address_1 <= "011001";
    ptr_deref_102_word_address_2 <= "011010";
    ptr_deref_102_word_address_3 <= "011011";
    ptr_deref_110_word_offset_0 <= "000000";
    ptr_deref_110_word_offset_1 <= "000001";
    ptr_deref_110_word_offset_2 <= "000010";
    ptr_deref_110_word_offset_3 <= "000011";
    ptr_deref_115_word_address_0 <= "011000";
    ptr_deref_115_word_address_1 <= "011001";
    ptr_deref_115_word_address_2 <= "011010";
    ptr_deref_115_word_address_3 <= "011011";
    ptr_deref_79_word_address_0 <= "011000";
    ptr_deref_79_word_address_1 <= "011001";
    ptr_deref_79_word_address_2 <= "011010";
    ptr_deref_79_word_address_3 <= "011011";
    ptr_deref_84_word_address_0 <= "011000";
    ptr_deref_84_word_address_1 <= "011001";
    ptr_deref_84_word_address_2 <= "011010";
    ptr_deref_84_word_address_3 <= "011011";
    ptr_deref_93_word_offset_0 <= "000000";
    ptr_deref_93_word_offset_1 <= "000001";
    ptr_deref_93_word_offset_2 <= "000010";
    ptr_deref_93_word_offset_3 <= "000011";
    xxfooxxbodyxxlptr_alloc_base_address <= "011000";
    array_obj_ref_107_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_9_103, dout => array_obj_ref_107_resized_base_address, req => array_obj_ref_107_base_resize_req_0, ack => array_obj_ref_107_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_107_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_107_root_address, dout => iNsTr_10_108, req => array_obj_ref_107_final_reg_req_0, ack => array_obj_ref_107_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_89_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_5_85, dout => array_obj_ref_89_resized_base_address, req => array_obj_ref_89_base_resize_req_0, ack => array_obj_ref_89_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_89_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_89_root_address, dout => iNsTr_6_90, req => array_obj_ref_89_final_reg_req_0, ack => array_obj_ref_89_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_110_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_10_108, dout => ptr_deref_110_resized_base_address, req => ptr_deref_110_base_resize_req_0, ack => ptr_deref_110_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_93_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_6_90, dout => ptr_deref_93_resized_base_address, req => ptr_deref_93_base_resize_req_0, ack => ptr_deref_93_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_119_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_12_116, dout => iNsTr_13_120, req => type_cast_119_inst_req_0, ack => type_cast_119_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_128_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_13_120, dout => type_cast_128_wire, req => type_cast_128_inst_req_0, ack => type_cast_128_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_72_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_71_wire, dout => iNsTr_2_73, req => type_cast_72_inst_req_0, ack => type_cast_72_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_76_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_2_73, dout => iNsTr_3_77, req => type_cast_76_inst_req_0, ack => type_cast_76_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_102_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_102_gather_scatter_ack_0 <= ptr_deref_102_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_102_data_0 & ptr_deref_102_data_1 & ptr_deref_102_data_2 & ptr_deref_102_data_3;
      iNsTr_9_103 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_110_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_110_gather_scatter_ack_0 <= ptr_deref_110_gather_scatter_req_0;
      aggregated_sig <= iNsTr_8_99;
      ptr_deref_110_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_110_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_110_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_110_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_110_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_110_root_address_inst_ack_0 <= ptr_deref_110_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_110_resized_base_address;
      ptr_deref_110_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_115_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_115_gather_scatter_ack_0 <= ptr_deref_115_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_115_data_0 & ptr_deref_115_data_1 & ptr_deref_115_data_2 & ptr_deref_115_data_3;
      iNsTr_12_116 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_79_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_79_gather_scatter_ack_0 <= ptr_deref_79_gather_scatter_req_0;
      aggregated_sig <= iNsTr_3_77;
      ptr_deref_79_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_79_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_79_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_79_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_84_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_84_gather_scatter_ack_0 <= ptr_deref_84_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_84_data_0 & ptr_deref_84_data_1 & ptr_deref_84_data_2 & ptr_deref_84_data_3;
      iNsTr_5_85 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_93_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_93_gather_scatter_ack_0 <= ptr_deref_93_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_93_data_0 & ptr_deref_93_data_1 & ptr_deref_93_data_2 & ptr_deref_93_data_3;
      iNsTr_7_94 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_93_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_93_root_address_inst_ack_0 <= ptr_deref_93_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_93_resized_base_address;
      ptr_deref_93_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_107_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_107_resized_base_address;
      array_obj_ref_107_root_address <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000100",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_107_root_address_inst_req_0,
          ackL => array_obj_ref_107_root_address_inst_ack_0,
          reqR => array_obj_ref_107_root_address_inst_req_1,
          ackR => array_obj_ref_107_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_89_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_89_resized_base_address;
      array_obj_ref_89_root_address <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000100",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_89_root_address_inst_req_0,
          ackL => array_obj_ref_89_root_address_inst_ack_0,
          reqR => array_obj_ref_89_root_address_inst_req_1,
          ackR => array_obj_ref_89_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_98_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_7_94;
      iNsTr_8_99 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_98_inst_req_0,
          ackL => binary_98_inst_ack_0,
          reqR => binary_98_inst_req_1,
          ackR => binary_98_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ptr_deref_110_addr_0 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_110_root_address;
      ptr_deref_110_word_address_0 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_110_addr_0_req_0,
          ackL => ptr_deref_110_addr_0_ack_0,
          reqR => ptr_deref_110_addr_0_req_1,
          ackR => ptr_deref_110_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ptr_deref_110_addr_1 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_110_root_address;
      ptr_deref_110_word_address_1 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_110_addr_1_req_0,
          ackL => ptr_deref_110_addr_1_ack_0,
          reqR => ptr_deref_110_addr_1_req_1,
          ackR => ptr_deref_110_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : ptr_deref_110_addr_2 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_110_root_address;
      ptr_deref_110_word_address_2 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_110_addr_2_req_0,
          ackL => ptr_deref_110_addr_2_ack_0,
          reqR => ptr_deref_110_addr_2_req_1,
          ackR => ptr_deref_110_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : ptr_deref_110_addr_3 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_110_root_address;
      ptr_deref_110_word_address_3 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000011",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_110_addr_3_req_0,
          ackL => ptr_deref_110_addr_3_ack_0,
          reqR => ptr_deref_110_addr_3_req_1,
          ackR => ptr_deref_110_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : ptr_deref_93_addr_0 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_93_root_address;
      ptr_deref_93_word_address_0 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_93_addr_0_req_0,
          ackL => ptr_deref_93_addr_0_ack_0,
          reqR => ptr_deref_93_addr_0_req_1,
          ackR => ptr_deref_93_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : ptr_deref_93_addr_1 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_93_root_address;
      ptr_deref_93_word_address_1 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_93_addr_1_req_0,
          ackL => ptr_deref_93_addr_1_ack_0,
          reqR => ptr_deref_93_addr_1_req_1,
          ackR => ptr_deref_93_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : ptr_deref_93_addr_2 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_93_root_address;
      ptr_deref_93_word_address_2 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_93_addr_2_req_0,
          ackL => ptr_deref_93_addr_2_ack_0,
          reqR => ptr_deref_93_addr_2_req_1,
          ackR => ptr_deref_93_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : ptr_deref_93_addr_3 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_93_root_address;
      ptr_deref_93_word_address_3 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000011",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_93_addr_3_req_0,
          ackL => ptr_deref_93_addr_3_ack_0,
          reqR => ptr_deref_93_addr_3_req_1,
          ackR => ptr_deref_93_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared load operator group (0) : ptr_deref_102_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_102_load_0_req_0;
      ptr_deref_102_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_102_load_0_req_1;
      ptr_deref_102_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_102_word_address_0;
      ptr_deref_102_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(15),
          mack => memory_space_1_lr_ack(15),
          maddr => memory_space_1_lr_addr(95 downto 90),
          mtag => memory_space_1_lr_tag(47 downto 45),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(15),
          mack => memory_space_1_lc_ack(15),
          mdata => memory_space_1_lc_data(127 downto 120),
          mtag => memory_space_1_lc_tag(47 downto 45),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_102_load_1 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_102_load_1_req_0;
      ptr_deref_102_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_102_load_1_req_1;
      ptr_deref_102_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_102_word_address_1;
      ptr_deref_102_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(14),
          mack => memory_space_1_lr_ack(14),
          maddr => memory_space_1_lr_addr(89 downto 84),
          mtag => memory_space_1_lr_tag(44 downto 42),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(14),
          mack => memory_space_1_lc_ack(14),
          mdata => memory_space_1_lc_data(119 downto 112),
          mtag => memory_space_1_lc_tag(44 downto 42),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_102_load_2 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_102_load_2_req_0;
      ptr_deref_102_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_102_load_2_req_1;
      ptr_deref_102_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_102_word_address_2;
      ptr_deref_102_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(13),
          mack => memory_space_1_lr_ack(13),
          maddr => memory_space_1_lr_addr(83 downto 78),
          mtag => memory_space_1_lr_tag(41 downto 39),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(13),
          mack => memory_space_1_lc_ack(13),
          mdata => memory_space_1_lc_data(111 downto 104),
          mtag => memory_space_1_lc_tag(41 downto 39),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_102_load_3 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_102_load_3_req_0;
      ptr_deref_102_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_102_load_3_req_1;
      ptr_deref_102_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_102_word_address_3;
      ptr_deref_102_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(12),
          mack => memory_space_1_lr_ack(12),
          maddr => memory_space_1_lr_addr(77 downto 72),
          mtag => memory_space_1_lr_tag(38 downto 36),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(12),
          mack => memory_space_1_lc_ack(12),
          mdata => memory_space_1_lc_data(103 downto 96),
          mtag => memory_space_1_lc_tag(38 downto 36),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_115_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_115_load_0_req_0;
      ptr_deref_115_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_115_load_0_req_1;
      ptr_deref_115_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_115_word_address_0;
      ptr_deref_115_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(11),
          mack => memory_space_1_lr_ack(11),
          maddr => memory_space_1_lr_addr(71 downto 66),
          mtag => memory_space_1_lr_tag(35 downto 33),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(11),
          mack => memory_space_1_lc_ack(11),
          mdata => memory_space_1_lc_data(95 downto 88),
          mtag => memory_space_1_lc_tag(35 downto 33),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_115_load_1 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_115_load_1_req_0;
      ptr_deref_115_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_115_load_1_req_1;
      ptr_deref_115_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_115_word_address_1;
      ptr_deref_115_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(10),
          mack => memory_space_1_lr_ack(10),
          maddr => memory_space_1_lr_addr(65 downto 60),
          mtag => memory_space_1_lr_tag(32 downto 30),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(10),
          mack => memory_space_1_lc_ack(10),
          mdata => memory_space_1_lc_data(87 downto 80),
          mtag => memory_space_1_lc_tag(32 downto 30),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_115_load_2 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_115_load_2_req_0;
      ptr_deref_115_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_115_load_2_req_1;
      ptr_deref_115_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_115_word_address_2;
      ptr_deref_115_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(9),
          mack => memory_space_1_lr_ack(9),
          maddr => memory_space_1_lr_addr(59 downto 54),
          mtag => memory_space_1_lr_tag(29 downto 27),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(9),
          mack => memory_space_1_lc_ack(9),
          mdata => memory_space_1_lc_data(79 downto 72),
          mtag => memory_space_1_lc_tag(29 downto 27),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_115_load_3 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_115_load_3_req_0;
      ptr_deref_115_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_115_load_3_req_1;
      ptr_deref_115_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_115_word_address_3;
      ptr_deref_115_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(8),
          mack => memory_space_1_lr_ack(8),
          maddr => memory_space_1_lr_addr(53 downto 48),
          mtag => memory_space_1_lr_tag(26 downto 24),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(8),
          mack => memory_space_1_lc_ack(8),
          mdata => memory_space_1_lc_data(71 downto 64),
          mtag => memory_space_1_lc_tag(26 downto 24),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared load operator group (8) : ptr_deref_84_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_84_load_0_req_0;
      ptr_deref_84_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_84_load_0_req_1;
      ptr_deref_84_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_84_word_address_0;
      ptr_deref_84_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(7),
          mack => memory_space_1_lr_ack(7),
          maddr => memory_space_1_lr_addr(47 downto 42),
          mtag => memory_space_1_lr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(7),
          mack => memory_space_1_lc_ack(7),
          mdata => memory_space_1_lc_data(63 downto 56),
          mtag => memory_space_1_lc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- shared load operator group (9) : ptr_deref_84_load_1 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_84_load_1_req_0;
      ptr_deref_84_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_84_load_1_req_1;
      ptr_deref_84_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_84_word_address_1;
      ptr_deref_84_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(6),
          mack => memory_space_1_lr_ack(6),
          maddr => memory_space_1_lr_addr(41 downto 36),
          mtag => memory_space_1_lr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(6),
          mack => memory_space_1_lc_ack(6),
          mdata => memory_space_1_lc_data(55 downto 48),
          mtag => memory_space_1_lc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    -- shared load operator group (10) : ptr_deref_84_load_2 
    LoadGroup10: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_84_load_2_req_0;
      ptr_deref_84_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_84_load_2_req_1;
      ptr_deref_84_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_84_word_address_2;
      ptr_deref_84_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(5),
          mack => memory_space_1_lr_ack(5),
          maddr => memory_space_1_lr_addr(35 downto 30),
          mtag => memory_space_1_lr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(5),
          mack => memory_space_1_lc_ack(5),
          mdata => memory_space_1_lc_data(47 downto 40),
          mtag => memory_space_1_lc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 10
    -- shared load operator group (11) : ptr_deref_84_load_3 
    LoadGroup11: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_84_load_3_req_0;
      ptr_deref_84_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_84_load_3_req_1;
      ptr_deref_84_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_84_word_address_3;
      ptr_deref_84_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(4),
          mack => memory_space_1_lr_ack(4),
          maddr => memory_space_1_lr_addr(29 downto 24),
          mtag => memory_space_1_lr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(4),
          mack => memory_space_1_lc_ack(4),
          mdata => memory_space_1_lc_data(39 downto 32),
          mtag => memory_space_1_lc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 11
    -- shared load operator group (12) : ptr_deref_93_load_0 
    LoadGroup12: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_93_load_0_req_0;
      ptr_deref_93_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_93_load_0_req_1;
      ptr_deref_93_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_93_word_address_0;
      ptr_deref_93_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(3),
          mack => memory_space_1_lr_ack(3),
          maddr => memory_space_1_lr_addr(23 downto 18),
          mtag => memory_space_1_lr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(3),
          mack => memory_space_1_lc_ack(3),
          mdata => memory_space_1_lc_data(31 downto 24),
          mtag => memory_space_1_lc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 12
    -- shared load operator group (13) : ptr_deref_93_load_1 
    LoadGroup13: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_93_load_1_req_0;
      ptr_deref_93_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_93_load_1_req_1;
      ptr_deref_93_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_93_word_address_1;
      ptr_deref_93_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(2),
          mack => memory_space_1_lr_ack(2),
          maddr => memory_space_1_lr_addr(17 downto 12),
          mtag => memory_space_1_lr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(2),
          mack => memory_space_1_lc_ack(2),
          mdata => memory_space_1_lc_data(23 downto 16),
          mtag => memory_space_1_lc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 13
    -- shared load operator group (14) : ptr_deref_93_load_2 
    LoadGroup14: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_93_load_2_req_0;
      ptr_deref_93_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_93_load_2_req_1;
      ptr_deref_93_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_93_word_address_2;
      ptr_deref_93_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(1),
          mack => memory_space_1_lr_ack(1),
          maddr => memory_space_1_lr_addr(11 downto 6),
          mtag => memory_space_1_lr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(1),
          mack => memory_space_1_lc_ack(1),
          mdata => memory_space_1_lc_data(15 downto 8),
          mtag => memory_space_1_lc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 14
    -- shared load operator group (15) : ptr_deref_93_load_3 
    LoadGroup15: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_93_load_3_req_0;
      ptr_deref_93_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_93_load_3_req_1;
      ptr_deref_93_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_93_word_address_3;
      ptr_deref_93_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(5 downto 0),
          mtag => memory_space_1_lr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 15
    -- shared store operator group (0) : ptr_deref_110_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_110_store_0_req_0;
      ptr_deref_110_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_110_store_0_req_1;
      ptr_deref_110_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_110_word_address_0;
      data_in <= ptr_deref_110_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(7),
          mack => memory_space_1_sr_ack(7),
          maddr => memory_space_1_sr_addr(47 downto 42),
          mdata => memory_space_1_sr_data(63 downto 56),
          mtag => memory_space_1_sr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(7),
          mack => memory_space_1_sc_ack(7),
          mtag => memory_space_1_sc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_110_store_1 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_110_store_1_req_0;
      ptr_deref_110_store_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_110_store_1_req_1;
      ptr_deref_110_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_110_word_address_1;
      data_in <= ptr_deref_110_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(6),
          mack => memory_space_1_sr_ack(6),
          maddr => memory_space_1_sr_addr(41 downto 36),
          mdata => memory_space_1_sr_data(55 downto 48),
          mtag => memory_space_1_sr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(6),
          mack => memory_space_1_sc_ack(6),
          mtag => memory_space_1_sc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_110_store_2 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_110_store_2_req_0;
      ptr_deref_110_store_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_110_store_2_req_1;
      ptr_deref_110_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_110_word_address_2;
      data_in <= ptr_deref_110_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(5),
          mack => memory_space_1_sr_ack(5),
          maddr => memory_space_1_sr_addr(35 downto 30),
          mdata => memory_space_1_sr_data(47 downto 40),
          mtag => memory_space_1_sr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(5),
          mack => memory_space_1_sc_ack(5),
          mtag => memory_space_1_sc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_110_store_3 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_110_store_3_req_0;
      ptr_deref_110_store_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_110_store_3_req_1;
      ptr_deref_110_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_110_word_address_3;
      data_in <= ptr_deref_110_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(4),
          mack => memory_space_1_sr_ack(4),
          maddr => memory_space_1_sr_addr(29 downto 24),
          mdata => memory_space_1_sr_data(39 downto 32),
          mtag => memory_space_1_sr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(4),
          mack => memory_space_1_sc_ack(4),
          mtag => memory_space_1_sc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_79_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_79_store_0_req_0;
      ptr_deref_79_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_79_store_0_req_1;
      ptr_deref_79_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_79_word_address_0;
      data_in <= ptr_deref_79_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(3),
          mack => memory_space_1_sr_ack(3),
          maddr => memory_space_1_sr_addr(23 downto 18),
          mdata => memory_space_1_sr_data(31 downto 24),
          mtag => memory_space_1_sr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(3),
          mack => memory_space_1_sc_ack(3),
          mtag => memory_space_1_sc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_79_store_1 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_79_store_1_req_0;
      ptr_deref_79_store_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_79_store_1_req_1;
      ptr_deref_79_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_79_word_address_1;
      data_in <= ptr_deref_79_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(2),
          mack => memory_space_1_sr_ack(2),
          maddr => memory_space_1_sr_addr(17 downto 12),
          mdata => memory_space_1_sr_data(23 downto 16),
          mtag => memory_space_1_sr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(2),
          mack => memory_space_1_sc_ack(2),
          mtag => memory_space_1_sc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_79_store_2 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_79_store_2_req_0;
      ptr_deref_79_store_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_79_store_2_req_1;
      ptr_deref_79_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_79_word_address_2;
      data_in <= ptr_deref_79_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(1),
          mack => memory_space_1_sr_ack(1),
          maddr => memory_space_1_sr_addr(11 downto 6),
          mdata => memory_space_1_sr_data(15 downto 8),
          mtag => memory_space_1_sr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(1),
          mack => memory_space_1_sc_ack(1),
          mtag => memory_space_1_sc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_79_store_3 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_79_store_3_req_0;
      ptr_deref_79_store_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_79_store_3_req_1;
      ptr_deref_79_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_79_word_address_3;
      data_in <= ptr_deref_79_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(5 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : simple_obj_ref_71_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_71_inst_req_0;
      simple_obj_ref_71_inst_ack_0 <= ack(0);
      simple_obj_ref_71_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => foo_in_pipe_read_req(0),
          oack => foo_in_pipe_read_ack(0),
          odata => foo_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : simple_obj_ref_126_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_126_inst_req_0;
      simple_obj_ref_126_inst_ack_0 <= ack(0);
      data_in <= type_cast_128_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => foo_out_pipe_write_req(0),
          oack => foo_out_pipe_write_ack(0),
          odata => foo_out_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_manager is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(1 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(1 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(1 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(1 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(1 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(11 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(11 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(71 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(35 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(11 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(11 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(95 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(35 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(47 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(23 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(7 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(23 downto 0);
    free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity free_queue_manager;
architecture Default of free_queue_manager is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_197_load_0_req_0 : boolean;
  signal ptr_deref_210_addr_1_req_1 : boolean;
  signal ptr_deref_183_load_2_ack_1 : boolean;
  signal simple_obj_ref_317_store_0_req_0 : boolean;
  signal ptr_deref_210_base_resize_req_0 : boolean;
  signal ptr_deref_315_addr_1_req_1 : boolean;
  signal ptr_deref_210_store_1_req_0 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal ptr_deref_210_store_1_ack_0 : boolean;
  signal ptr_deref_210_addr_2_ack_0 : boolean;
  signal addr_of_202_final_reg_ack_0 : boolean;
  signal ptr_deref_210_addr_0_req_0 : boolean;
  signal ptr_deref_183_load_2_req_1 : boolean;
  signal ptr_deref_210_addr_0_ack_1 : boolean;
  signal ptr_deref_210_addr_2_ack_1 : boolean;
  signal ptr_deref_210_addr_2_req_0 : boolean;
  signal ptr_deref_210_addr_1_ack_0 : boolean;
  signal ptr_deref_210_addr_0_ack_0 : boolean;
  signal ptr_deref_210_addr_0_req_1 : boolean;
  signal ptr_deref_210_addr_1_ack_1 : boolean;
  signal array_obj_ref_201_offset_inst_ack_0 : boolean;
  signal simple_obj_ref_306_load_0_ack_0 : boolean;
  signal ptr_deref_315_addr_1_ack_1 : boolean;
  signal ptr_deref_210_store_0_req_0 : boolean;
  signal ptr_deref_210_store_0_ack_0 : boolean;
  signal ptr_deref_210_store_3_req_0 : boolean;
  signal ptr_deref_210_store_3_ack_0 : boolean;
  signal ptr_deref_210_addr_2_req_1 : boolean;
  signal ptr_deref_210_store_2_req_0 : boolean;
  signal ptr_deref_210_store_2_ack_0 : boolean;
  signal ptr_deref_210_addr_3_req_1 : boolean;
  signal ptr_deref_210_addr_3_ack_1 : boolean;
  signal simple_obj_ref_317_gather_scatter_ack_0 : boolean;
  signal ptr_deref_324_load_0_req_0 : boolean;
  signal ptr_deref_210_addr_3_req_0 : boolean;
  signal ptr_deref_210_addr_3_ack_0 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal ptr_deref_210_gather_scatter_req_0 : boolean;
  signal ptr_deref_210_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_317_gather_scatter_req_0 : boolean;
  signal ptr_deref_324_load_0_ack_0 : boolean;
  signal simple_obj_ref_317_store_0_ack_0 : boolean;
  signal simple_obj_ref_317_store_0_req_1 : boolean;
  signal array_obj_ref_207_final_reg_ack_0 : boolean;
  signal array_obj_ref_201_offset_inst_req_0 : boolean;
  signal simple_obj_ref_306_load_0_req_1 : boolean;
  signal ptr_deref_210_addr_1_req_0 : boolean;
  signal ptr_deref_183_load_1_ack_1 : boolean;
  signal simple_obj_ref_306_load_0_ack_1 : boolean;
  signal array_obj_ref_201_root_address_inst_ack_0 : boolean;
  signal ptr_deref_324_load_2_req_0 : boolean;
  signal if_stmt_354_branch_req_0 : boolean;
  signal ptr_deref_197_load_1_ack_1 : boolean;
  signal ptr_deref_183_load_1_req_1 : boolean;
  signal array_obj_ref_201_index_0_scale_ack_1 : boolean;
  signal ptr_deref_324_load_1_req_0 : boolean;
  signal array_obj_ref_201_root_address_inst_req_0 : boolean;
  signal ptr_deref_197_load_1_req_1 : boolean;
  signal ptr_deref_210_base_resize_ack_0 : boolean;
  signal ptr_deref_183_load_0_ack_1 : boolean;
  signal ptr_deref_183_load_0_req_1 : boolean;
  signal ptr_deref_315_addr_3_ack_0 : boolean;
  signal ptr_deref_315_load_3_req_1 : boolean;
  signal array_obj_ref_201_index_0_scale_req_1 : boolean;
  signal ptr_deref_315_addr_2_req_0 : boolean;
  signal simple_obj_ref_306_gather_scatter_req_0 : boolean;
  signal ptr_deref_315_addr_3_req_1 : boolean;
  signal ptr_deref_315_addr_3_ack_1 : boolean;
  signal simple_obj_ref_306_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_201_index_0_scale_ack_0 : boolean;
  signal ptr_deref_324_load_2_req_1 : boolean;
  signal ptr_deref_324_load_2_ack_0 : boolean;
  signal ptr_deref_197_load_0_ack_1 : boolean;
  signal ptr_deref_315_gather_scatter_req_0 : boolean;
  signal ptr_deref_197_load_1_ack_0 : boolean;
  signal ptr_deref_197_load_1_req_0 : boolean;
  signal ptr_deref_197_load_2_ack_1 : boolean;
  signal addr_of_202_final_reg_req_0 : boolean;
  signal array_obj_ref_201_index_0_scale_req_0 : boolean;
  signal array_obj_ref_207_final_reg_req_0 : boolean;
  signal ptr_deref_343_load_0_ack_0 : boolean;
  signal addr_of_193_final_reg_ack_0 : boolean;
  signal ptr_deref_315_addr_2_ack_0 : boolean;
  signal addr_of_193_final_reg_req_0 : boolean;
  signal ptr_deref_315_load_3_ack_1 : boolean;
  signal ptr_deref_315_addr_3_req_0 : boolean;
  signal ptr_deref_197_load_0_req_1 : boolean;
  signal ptr_deref_210_root_address_inst_ack_0 : boolean;
  signal ptr_deref_183_load_3_ack_0 : boolean;
  signal array_obj_ref_192_root_address_inst_ack_0 : boolean;
  signal ptr_deref_183_load_3_req_0 : boolean;
  signal array_obj_ref_192_root_address_inst_req_0 : boolean;
  signal ptr_deref_210_root_address_inst_req_0 : boolean;
  signal array_obj_ref_207_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_207_root_address_inst_req_0 : boolean;
  signal ptr_deref_315_addr_0_req_0 : boolean;
  signal ptr_deref_183_load_2_ack_0 : boolean;
  signal binary_188_inst_ack_1 : boolean;
  signal ptr_deref_315_addr_2_ack_1 : boolean;
  signal array_obj_ref_192_offset_inst_ack_0 : boolean;
  signal ptr_deref_315_addr_2_req_1 : boolean;
  signal array_obj_ref_192_offset_inst_req_0 : boolean;
  signal binary_188_inst_req_1 : boolean;
  signal ptr_deref_183_load_2_req_0 : boolean;
  signal ptr_deref_343_load_0_req_0 : boolean;
  signal array_obj_ref_207_base_resize_ack_0 : boolean;
  signal binary_188_inst_ack_0 : boolean;
  signal array_obj_ref_207_base_resize_req_0 : boolean;
  signal simple_obj_ref_306_load_0_req_0 : boolean;
  signal array_obj_ref_192_index_0_scale_ack_1 : boolean;
  signal binary_188_inst_req_0 : boolean;
  signal array_obj_ref_192_index_0_scale_req_1 : boolean;
  signal array_obj_ref_192_index_0_scale_ack_0 : boolean;
  signal ptr_deref_197_gather_scatter_ack_0 : boolean;
  signal ptr_deref_197_load_3_ack_0 : boolean;
  signal ptr_deref_197_gather_scatter_req_0 : boolean;
  signal ptr_deref_197_load_3_req_0 : boolean;
  signal ptr_deref_324_load_1_ack_0 : boolean;
  signal array_obj_ref_192_index_0_scale_req_0 : boolean;
  signal ptr_deref_343_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_201_index_0_resize_ack_0 : boolean;
  signal ptr_deref_183_load_1_ack_0 : boolean;
  signal array_obj_ref_201_index_0_resize_req_0 : boolean;
  signal ptr_deref_197_load_3_ack_1 : boolean;
  signal ptr_deref_197_load_2_ack_0 : boolean;
  signal ptr_deref_183_load_1_req_0 : boolean;
  signal simple_obj_ref_317_store_0_ack_1 : boolean;
  signal array_obj_ref_192_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_192_index_0_resize_req_0 : boolean;
  signal ptr_deref_197_load_3_req_1 : boolean;
  signal ptr_deref_197_load_2_req_0 : boolean;
  signal ptr_deref_343_load_0_ack_1 : boolean;
  signal ptr_deref_324_load_3_req_1 : boolean;
  signal ptr_deref_324_gather_scatter_ack_0 : boolean;
  signal ptr_deref_324_load_2_ack_1 : boolean;
  signal ptr_deref_324_load_3_req_0 : boolean;
  signal ptr_deref_183_load_0_ack_0 : boolean;
  signal ptr_deref_183_load_0_req_0 : boolean;
  signal ptr_deref_183_gather_scatter_ack_0 : boolean;
  signal ptr_deref_324_load_1_req_1 : boolean;
  signal ptr_deref_315_root_address_inst_ack_0 : boolean;
  signal ptr_deref_375_store_1_req_0 : boolean;
  signal ptr_deref_375_store_2_ack_1 : boolean;
  signal ptr_deref_375_store_1_ack_0 : boolean;
  signal ptr_deref_383_load_1_ack_0 : boolean;
  signal if_stmt_174_branch_ack_0 : boolean;
  signal ptr_deref_183_gather_scatter_req_0 : boolean;
  signal ptr_deref_197_load_2_req_1 : boolean;
  signal ptr_deref_315_load_0_req_0 : boolean;
  signal ptr_deref_183_load_3_ack_1 : boolean;
  signal type_cast_347_inst_req_0 : boolean;
  signal ptr_deref_315_gather_scatter_ack_0 : boolean;
  signal ptr_deref_197_load_0_ack_0 : boolean;
  signal ptr_deref_183_load_3_req_1 : boolean;
  signal ptr_deref_324_load_3_ack_0 : boolean;
  signal type_cast_337_inst_req_0 : boolean;
  signal type_cast_337_inst_ack_0 : boolean;
  signal array_obj_ref_311_base_resize_req_0 : boolean;
  signal ptr_deref_315_load_0_ack_0 : boolean;
  signal ptr_deref_315_addr_0_ack_0 : boolean;
  signal array_obj_ref_311_base_resize_ack_0 : boolean;
  signal ptr_deref_315_load_1_req_0 : boolean;
  signal ptr_deref_315_load_1_ack_0 : boolean;
  signal ptr_deref_315_addr_0_req_1 : boolean;
  signal ptr_deref_375_store_3_ack_0 : boolean;
  signal array_obj_ref_311_root_address_inst_req_0 : boolean;
  signal array_obj_ref_311_root_address_inst_ack_0 : boolean;
  signal if_stmt_354_branch_ack_0 : boolean;
  signal simple_obj_ref_367_inst_req_0 : boolean;
  signal array_obj_ref_311_final_reg_req_0 : boolean;
  signal type_cast_368_inst_req_0 : boolean;
  signal array_obj_ref_311_final_reg_ack_0 : boolean;
  signal ptr_deref_315_load_2_req_0 : boolean;
  signal ptr_deref_315_load_2_ack_0 : boolean;
  signal ptr_deref_324_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_367_inst_ack_0 : boolean;
  signal ptr_deref_324_load_0_req_1 : boolean;
  signal ptr_deref_315_addr_0_ack_1 : boolean;
  signal ptr_deref_315_load_3_req_0 : boolean;
  signal ptr_deref_324_load_0_ack_1 : boolean;
  signal simple_obj_ref_335_inst_req_0 : boolean;
  signal type_cast_368_inst_ack_0 : boolean;
  signal simple_obj_ref_335_inst_ack_0 : boolean;
  signal ptr_deref_315_load_3_ack_0 : boolean;
  signal ptr_deref_375_store_3_req_1 : boolean;
  signal type_cast_372_inst_req_0 : boolean;
  signal type_cast_347_inst_ack_0 : boolean;
  signal ptr_deref_375_store_1_req_1 : boolean;
  signal ptr_deref_315_load_0_req_1 : boolean;
  signal type_cast_372_inst_ack_0 : boolean;
  signal ptr_deref_315_load_0_ack_1 : boolean;
  signal ptr_deref_315_base_resize_req_0 : boolean;
  signal ptr_deref_315_base_resize_ack_0 : boolean;
  signal simple_obj_ref_379_load_0_req_1 : boolean;
  signal simple_obj_ref_379_load_0_ack_1 : boolean;
  signal ptr_deref_343_load_0_req_1 : boolean;
  signal ptr_deref_375_store_0_ack_1 : boolean;
  signal ptr_deref_315_load_1_req_1 : boolean;
  signal ptr_deref_375_store_1_ack_1 : boolean;
  signal simple_obj_ref_379_load_0_ack_0 : boolean;
  signal ptr_deref_375_store_0_req_1 : boolean;
  signal ptr_deref_375_store_3_req_0 : boolean;
  signal ptr_deref_375_store_2_req_1 : boolean;
  signal ptr_deref_315_load_1_ack_1 : boolean;
  signal ptr_deref_375_gather_scatter_req_0 : boolean;
  signal ptr_deref_375_store_0_req_0 : boolean;
  signal ptr_deref_315_root_address_inst_req_0 : boolean;
  signal binary_352_inst_req_0 : boolean;
  signal binary_352_inst_ack_0 : boolean;
  signal ptr_deref_375_gather_scatter_ack_0 : boolean;
  signal binary_352_inst_req_1 : boolean;
  signal ptr_deref_383_load_2_ack_0 : boolean;
  signal binary_352_inst_ack_1 : boolean;
  signal if_stmt_354_branch_ack_1 : boolean;
  signal ptr_deref_375_store_3_ack_1 : boolean;
  signal ptr_deref_324_load_1_ack_1 : boolean;
  signal ptr_deref_343_gather_scatter_req_0 : boolean;
  signal ptr_deref_375_store_2_req_0 : boolean;
  signal ptr_deref_375_store_2_ack_0 : boolean;
  signal simple_obj_ref_379_load_0_req_0 : boolean;
  signal ptr_deref_383_load_1_req_0 : boolean;
  signal ptr_deref_375_store_0_ack_0 : boolean;
  signal ptr_deref_383_load_3_req_1 : boolean;
  signal ptr_deref_383_load_3_ack_1 : boolean;
  signal ptr_deref_383_gather_scatter_req_0 : boolean;
  signal ptr_deref_383_gather_scatter_ack_0 : boolean;
  signal ptr_deref_315_load_2_req_1 : boolean;
  signal ptr_deref_383_load_2_req_0 : boolean;
  signal ptr_deref_383_load_0_ack_1 : boolean;
  signal ptr_deref_383_load_3_ack_0 : boolean;
  signal ptr_deref_324_load_3_ack_1 : boolean;
  signal ptr_deref_383_load_0_req_1 : boolean;
  signal ptr_deref_383_load_3_req_0 : boolean;
  signal ptr_deref_383_load_0_req_0 : boolean;
  signal ptr_deref_383_load_0_ack_0 : boolean;
  signal simple_obj_ref_379_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_379_gather_scatter_ack_0 : boolean;
  signal ptr_deref_315_addr_1_ack_0 : boolean;
  signal ptr_deref_383_load_1_req_1 : boolean;
  signal ptr_deref_383_load_1_ack_1 : boolean;
  signal ptr_deref_315_load_2_ack_1 : boolean;
  signal ptr_deref_315_addr_1_req_0 : boolean;
  signal ptr_deref_383_load_2_req_1 : boolean;
  signal ptr_deref_383_load_2_ack_1 : boolean;
  signal array_obj_ref_388_base_resize_req_0 : boolean;
  signal ptr_deref_156_gather_scatter_req_0 : boolean;
  signal ptr_deref_156_gather_scatter_ack_0 : boolean;
  signal ptr_deref_156_store_0_req_0 : boolean;
  signal ptr_deref_156_store_0_ack_0 : boolean;
  signal ptr_deref_156_store_1_req_0 : boolean;
  signal ptr_deref_156_store_1_ack_0 : boolean;
  signal ptr_deref_156_store_2_req_0 : boolean;
  signal ptr_deref_156_store_2_ack_0 : boolean;
  signal ptr_deref_156_store_3_req_0 : boolean;
  signal ptr_deref_156_store_3_ack_0 : boolean;
  signal ptr_deref_156_store_0_req_1 : boolean;
  signal ptr_deref_156_store_0_ack_1 : boolean;
  signal ptr_deref_156_store_1_req_1 : boolean;
  signal ptr_deref_156_store_1_ack_1 : boolean;
  signal ptr_deref_156_store_2_req_1 : boolean;
  signal ptr_deref_156_store_2_ack_1 : boolean;
  signal ptr_deref_156_store_3_req_1 : boolean;
  signal ptr_deref_156_store_3_ack_1 : boolean;
  signal ptr_deref_163_load_0_req_0 : boolean;
  signal ptr_deref_163_load_0_ack_0 : boolean;
  signal ptr_deref_163_load_1_req_0 : boolean;
  signal ptr_deref_163_load_1_ack_0 : boolean;
  signal ptr_deref_163_load_2_req_0 : boolean;
  signal ptr_deref_163_load_2_ack_0 : boolean;
  signal ptr_deref_163_load_3_req_0 : boolean;
  signal ptr_deref_163_load_3_ack_0 : boolean;
  signal ptr_deref_163_load_0_req_1 : boolean;
  signal ptr_deref_163_load_0_ack_1 : boolean;
  signal ptr_deref_163_load_1_req_1 : boolean;
  signal ptr_deref_163_load_1_ack_1 : boolean;
  signal ptr_deref_163_load_2_req_1 : boolean;
  signal ptr_deref_163_load_2_ack_1 : boolean;
  signal ptr_deref_163_load_3_req_1 : boolean;
  signal ptr_deref_163_load_3_ack_1 : boolean;
  signal ptr_deref_163_gather_scatter_req_0 : boolean;
  signal ptr_deref_163_gather_scatter_ack_0 : boolean;
  signal type_cast_168_inst_req_0 : boolean;
  signal type_cast_168_inst_ack_0 : boolean;
  signal type_cast_168_inst_req_1 : boolean;
  signal type_cast_168_inst_ack_1 : boolean;
  signal binary_171_inst_req_0 : boolean;
  signal binary_171_inst_ack_0 : boolean;
  signal binary_171_inst_req_1 : boolean;
  signal binary_171_inst_ack_1 : boolean;
  signal if_stmt_174_branch_req_0 : boolean;
  signal if_stmt_174_branch_ack_1 : boolean;
  signal ptr_deref_210_store_0_req_1 : boolean;
  signal ptr_deref_210_store_0_ack_1 : boolean;
  signal ptr_deref_210_store_1_req_1 : boolean;
  signal ptr_deref_210_store_1_ack_1 : boolean;
  signal ptr_deref_210_store_2_req_1 : boolean;
  signal ptr_deref_210_store_2_ack_1 : boolean;
  signal ptr_deref_210_store_3_req_1 : boolean;
  signal ptr_deref_210_store_3_ack_1 : boolean;
  signal ptr_deref_215_load_0_req_0 : boolean;
  signal ptr_deref_215_load_0_ack_0 : boolean;
  signal ptr_deref_215_load_1_req_0 : boolean;
  signal ptr_deref_215_load_1_ack_0 : boolean;
  signal ptr_deref_215_load_2_req_0 : boolean;
  signal ptr_deref_215_load_2_ack_0 : boolean;
  signal ptr_deref_215_load_3_req_0 : boolean;
  signal ptr_deref_215_load_3_ack_0 : boolean;
  signal ptr_deref_215_load_0_req_1 : boolean;
  signal ptr_deref_215_load_0_ack_1 : boolean;
  signal ptr_deref_215_load_1_req_1 : boolean;
  signal ptr_deref_215_load_1_ack_1 : boolean;
  signal ptr_deref_215_load_2_req_1 : boolean;
  signal ptr_deref_215_load_2_ack_1 : boolean;
  signal ptr_deref_215_load_3_req_1 : boolean;
  signal ptr_deref_215_load_3_ack_1 : boolean;
  signal ptr_deref_215_gather_scatter_req_0 : boolean;
  signal ptr_deref_215_gather_scatter_ack_0 : boolean;
  signal binary_220_inst_req_0 : boolean;
  signal binary_220_inst_ack_0 : boolean;
  signal binary_220_inst_req_1 : boolean;
  signal binary_220_inst_ack_1 : boolean;
  signal ptr_deref_223_gather_scatter_req_0 : boolean;
  signal ptr_deref_223_gather_scatter_ack_0 : boolean;
  signal ptr_deref_223_store_0_req_0 : boolean;
  signal ptr_deref_223_store_0_ack_0 : boolean;
  signal ptr_deref_223_store_1_req_0 : boolean;
  signal ptr_deref_223_store_1_ack_0 : boolean;
  signal ptr_deref_223_store_2_req_0 : boolean;
  signal ptr_deref_223_store_2_ack_0 : boolean;
  signal ptr_deref_223_store_3_req_0 : boolean;
  signal ptr_deref_223_store_3_ack_0 : boolean;
  signal ptr_deref_223_store_0_req_1 : boolean;
  signal ptr_deref_223_store_0_ack_1 : boolean;
  signal ptr_deref_223_store_1_req_1 : boolean;
  signal ptr_deref_223_store_1_ack_1 : boolean;
  signal ptr_deref_223_store_2_req_1 : boolean;
  signal ptr_deref_223_store_2_ack_1 : boolean;
  signal ptr_deref_223_store_3_req_1 : boolean;
  signal ptr_deref_223_store_3_ack_1 : boolean;
  signal ptr_deref_235_gather_scatter_req_0 : boolean;
  signal ptr_deref_235_gather_scatter_ack_0 : boolean;
  signal ptr_deref_235_store_0_req_0 : boolean;
  signal ptr_deref_235_store_0_ack_0 : boolean;
  signal ptr_deref_235_store_1_req_0 : boolean;
  signal ptr_deref_235_store_1_ack_0 : boolean;
  signal ptr_deref_235_store_2_req_0 : boolean;
  signal ptr_deref_235_store_2_ack_0 : boolean;
  signal ptr_deref_235_store_3_req_0 : boolean;
  signal ptr_deref_235_store_3_ack_0 : boolean;
  signal ptr_deref_235_store_0_req_1 : boolean;
  signal ptr_deref_235_store_0_ack_1 : boolean;
  signal ptr_deref_235_store_1_req_1 : boolean;
  signal ptr_deref_235_store_1_ack_1 : boolean;
  signal ptr_deref_235_store_2_req_1 : boolean;
  signal ptr_deref_235_store_2_ack_1 : boolean;
  signal ptr_deref_235_store_3_req_1 : boolean;
  signal ptr_deref_235_store_3_ack_1 : boolean;
  signal simple_obj_ref_243_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_243_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_243_store_0_req_0 : boolean;
  signal simple_obj_ref_243_store_0_ack_0 : boolean;
  signal simple_obj_ref_243_store_0_req_1 : boolean;
  signal simple_obj_ref_243_store_0_ack_1 : boolean;
  signal simple_obj_ref_254_inst_req_0 : boolean;
  signal simple_obj_ref_254_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal ptr_deref_258_gather_scatter_req_0 : boolean;
  signal ptr_deref_258_gather_scatter_ack_0 : boolean;
  signal ptr_deref_258_store_0_req_0 : boolean;
  signal ptr_deref_258_store_0_ack_0 : boolean;
  signal ptr_deref_258_store_0_req_1 : boolean;
  signal ptr_deref_258_store_0_ack_1 : boolean;
  signal ptr_deref_263_load_0_req_0 : boolean;
  signal ptr_deref_263_load_0_ack_0 : boolean;
  signal ptr_deref_263_load_0_req_1 : boolean;
  signal ptr_deref_263_load_0_ack_1 : boolean;
  signal ptr_deref_263_gather_scatter_req_0 : boolean;
  signal ptr_deref_263_gather_scatter_ack_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal binary_272_inst_req_0 : boolean;
  signal binary_272_inst_ack_0 : boolean;
  signal binary_272_inst_req_1 : boolean;
  signal binary_272_inst_ack_1 : boolean;
  signal if_stmt_274_branch_req_0 : boolean;
  signal if_stmt_274_branch_ack_1 : boolean;
  signal if_stmt_274_branch_ack_0 : boolean;
  signal simple_obj_ref_282_load_0_req_0 : boolean;
  signal simple_obj_ref_282_load_0_ack_0 : boolean;
  signal simple_obj_ref_282_load_0_req_1 : boolean;
  signal simple_obj_ref_282_load_0_ack_1 : boolean;
  signal simple_obj_ref_282_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_282_gather_scatter_ack_0 : boolean;
  signal ptr_deref_285_gather_scatter_req_0 : boolean;
  signal ptr_deref_285_gather_scatter_ack_0 : boolean;
  signal ptr_deref_285_store_0_req_0 : boolean;
  signal ptr_deref_285_store_0_ack_0 : boolean;
  signal ptr_deref_285_store_1_req_0 : boolean;
  signal ptr_deref_285_store_1_ack_0 : boolean;
  signal ptr_deref_285_store_2_req_0 : boolean;
  signal ptr_deref_285_store_2_ack_0 : boolean;
  signal ptr_deref_285_store_3_req_0 : boolean;
  signal ptr_deref_285_store_3_ack_0 : boolean;
  signal ptr_deref_285_store_0_req_1 : boolean;
  signal ptr_deref_285_store_0_ack_1 : boolean;
  signal ptr_deref_285_store_1_req_1 : boolean;
  signal ptr_deref_285_store_1_ack_1 : boolean;
  signal ptr_deref_285_store_2_req_1 : boolean;
  signal ptr_deref_285_store_2_ack_1 : boolean;
  signal ptr_deref_285_store_3_req_1 : boolean;
  signal ptr_deref_285_store_3_ack_1 : boolean;
  signal simple_obj_ref_289_load_0_req_0 : boolean;
  signal simple_obj_ref_289_load_0_ack_0 : boolean;
  signal simple_obj_ref_289_load_0_req_1 : boolean;
  signal simple_obj_ref_289_load_0_ack_1 : boolean;
  signal simple_obj_ref_289_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_289_gather_scatter_ack_0 : boolean;
  signal type_cast_293_inst_req_0 : boolean;
  signal type_cast_293_inst_ack_0 : boolean;
  signal type_cast_293_inst_req_1 : boolean;
  signal type_cast_293_inst_ack_1 : boolean;
  signal binary_296_inst_req_0 : boolean;
  signal binary_296_inst_ack_0 : boolean;
  signal binary_296_inst_req_1 : boolean;
  signal binary_296_inst_ack_1 : boolean;
  signal if_stmt_298_branch_req_0 : boolean;
  signal if_stmt_298_branch_ack_1 : boolean;
  signal if_stmt_298_branch_ack_0 : boolean;
  signal array_obj_ref_388_base_resize_ack_0 : boolean;
  signal array_obj_ref_388_root_address_inst_req_0 : boolean;
  signal array_obj_ref_388_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_388_final_reg_req_0 : boolean;
  signal array_obj_ref_388_final_reg_ack_0 : boolean;
  signal ptr_deref_391_base_resize_req_0 : boolean;
  signal ptr_deref_391_base_resize_ack_0 : boolean;
  signal ptr_deref_391_root_address_inst_req_0 : boolean;
  signal ptr_deref_391_root_address_inst_ack_0 : boolean;
  signal ptr_deref_391_addr_0_req_0 : boolean;
  signal ptr_deref_391_addr_0_ack_0 : boolean;
  signal ptr_deref_391_addr_0_req_1 : boolean;
  signal ptr_deref_391_addr_0_ack_1 : boolean;
  signal ptr_deref_391_addr_1_req_0 : boolean;
  signal ptr_deref_391_addr_1_ack_0 : boolean;
  signal ptr_deref_391_addr_1_req_1 : boolean;
  signal ptr_deref_391_addr_1_ack_1 : boolean;
  signal ptr_deref_391_addr_2_req_0 : boolean;
  signal ptr_deref_391_addr_2_ack_0 : boolean;
  signal ptr_deref_391_addr_2_req_1 : boolean;
  signal ptr_deref_391_addr_2_ack_1 : boolean;
  signal ptr_deref_391_addr_3_req_0 : boolean;
  signal ptr_deref_391_addr_3_ack_0 : boolean;
  signal ptr_deref_391_addr_3_req_1 : boolean;
  signal ptr_deref_391_addr_3_ack_1 : boolean;
  signal ptr_deref_391_gather_scatter_req_0 : boolean;
  signal ptr_deref_391_gather_scatter_ack_0 : boolean;
  signal ptr_deref_391_store_0_req_0 : boolean;
  signal ptr_deref_391_store_0_ack_0 : boolean;
  signal ptr_deref_391_store_1_req_0 : boolean;
  signal ptr_deref_391_store_1_ack_0 : boolean;
  signal ptr_deref_391_store_2_req_0 : boolean;
  signal ptr_deref_391_store_2_ack_0 : boolean;
  signal ptr_deref_391_store_3_req_0 : boolean;
  signal ptr_deref_391_store_3_ack_0 : boolean;
  signal ptr_deref_391_store_0_req_1 : boolean;
  signal ptr_deref_391_store_0_ack_1 : boolean;
  signal ptr_deref_391_store_1_req_1 : boolean;
  signal ptr_deref_391_store_1_ack_1 : boolean;
  signal ptr_deref_391_store_2_req_1 : boolean;
  signal ptr_deref_391_store_2_ack_1 : boolean;
  signal ptr_deref_391_store_3_req_1 : boolean;
  signal ptr_deref_391_store_3_ack_1 : boolean;
  signal ptr_deref_396_load_0_req_0 : boolean;
  signal ptr_deref_396_load_0_ack_0 : boolean;
  signal ptr_deref_396_load_1_req_0 : boolean;
  signal ptr_deref_396_load_1_ack_0 : boolean;
  signal ptr_deref_396_load_2_req_0 : boolean;
  signal ptr_deref_396_load_2_ack_0 : boolean;
  signal ptr_deref_396_load_3_req_0 : boolean;
  signal ptr_deref_396_load_3_ack_0 : boolean;
  signal ptr_deref_396_load_0_req_1 : boolean;
  signal ptr_deref_396_load_0_ack_1 : boolean;
  signal ptr_deref_396_load_1_req_1 : boolean;
  signal ptr_deref_396_load_1_ack_1 : boolean;
  signal ptr_deref_396_load_2_req_1 : boolean;
  signal ptr_deref_396_load_2_ack_1 : boolean;
  signal ptr_deref_396_load_3_req_1 : boolean;
  signal ptr_deref_396_load_3_ack_1 : boolean;
  signal ptr_deref_396_gather_scatter_req_0 : boolean;
  signal ptr_deref_396_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_398_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_398_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_398_store_0_req_0 : boolean;
  signal simple_obj_ref_398_store_0_ack_0 : boolean;
  signal simple_obj_ref_398_store_0_req_1 : boolean;
  signal simple_obj_ref_398_store_0_ack_1 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  free_queue_manager_CP_614: Block -- control-path 
    signal free_queue_manager_CP_614_start: Boolean;
    signal Xentry_615_symbol: Boolean;
    signal Xexit_616_symbol: Boolean;
    signal branch_block_stmt_134_617_symbol : Boolean;
    -- 
  begin -- 
    free_queue_manager_CP_614_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_615_symbol  <= free_queue_manager_CP_614_start; -- transition $entry
    branch_block_stmt_134_617: Block -- branch_block_stmt_134 
      signal branch_block_stmt_134_617_start: Boolean;
      signal Xentry_618_symbol: Boolean;
      signal Xexit_619_symbol: Boolean;
      signal branch_block_stmt_134_x_xentry_x_xx_x620_symbol : Boolean;
      signal branch_block_stmt_134_x_xexit_x_xx_x621_symbol : Boolean;
      signal assign_stmt_142_to_assign_stmt_158_x_xentry_x_xx_x622_symbol : Boolean;
      signal assign_stmt_142_to_assign_stmt_158_x_xexit_x_xx_x623_symbol : Boolean;
      signal bb_0_bb_1_624_symbol : Boolean;
      signal merge_stmt_160_x_xexit_x_xx_x625_symbol : Boolean;
      signal assign_stmt_164_to_assign_stmt_173_x_xentry_x_xx_x626_symbol : Boolean;
      signal assign_stmt_164_to_assign_stmt_173_x_xexit_x_xx_x627_symbol : Boolean;
      signal if_stmt_174_x_xentry_x_xx_x628_symbol : Boolean;
      signal if_stmt_174_x_xexit_x_xx_x629_symbol : Boolean;
      signal merge_stmt_180_x_xentry_x_xx_x630_symbol : Boolean;
      signal merge_stmt_180_x_xexit_x_xx_x631_symbol : Boolean;
      signal assign_stmt_184_to_assign_stmt_225_x_xentry_x_xx_x632_symbol : Boolean;
      signal assign_stmt_184_to_assign_stmt_225_x_xexit_x_xx_x633_symbol : Boolean;
      signal bb_2_bb_1_634_symbol : Boolean;
      signal merge_stmt_227_x_xexit_x_xx_x635_symbol : Boolean;
      signal assign_stmt_233_to_assign_stmt_245_x_xentry_x_xx_x636_symbol : Boolean;
      signal assign_stmt_233_to_assign_stmt_245_x_xexit_x_xx_x637_symbol : Boolean;
      signal bb_3_bb_4_638_symbol : Boolean;
      signal merge_stmt_247_x_xexit_x_xx_x639_symbol : Boolean;
      signal assign_stmt_252_x_xentry_x_xx_x640_symbol : Boolean;
      signal assign_stmt_252_x_xexit_x_xx_x641_symbol : Boolean;
      signal assign_stmt_256_x_xentry_x_xx_x642_symbol : Boolean;
      signal assign_stmt_256_x_xexit_x_xx_x643_symbol : Boolean;
      signal assign_stmt_260_to_assign_stmt_273_x_xentry_x_xx_x644_symbol : Boolean;
      signal assign_stmt_260_to_assign_stmt_273_x_xexit_x_xx_x645_symbol : Boolean;
      signal if_stmt_274_x_xentry_x_xx_x646_symbol : Boolean;
      signal if_stmt_274_x_xexit_x_xx_x647_symbol : Boolean;
      signal merge_stmt_280_x_xentry_x_xx_x648_symbol : Boolean;
      signal merge_stmt_280_x_xexit_x_xx_x649_symbol : Boolean;
      signal assign_stmt_283_to_assign_stmt_297_x_xentry_x_xx_x650_symbol : Boolean;
      signal assign_stmt_283_to_assign_stmt_297_x_xexit_x_xx_x651_symbol : Boolean;
      signal if_stmt_298_x_xentry_x_xx_x652_symbol : Boolean;
      signal if_stmt_298_x_xexit_x_xx_x653_symbol : Boolean;
      signal merge_stmt_304_x_xentry_x_xx_x654_symbol : Boolean;
      signal merge_stmt_304_x_xexit_x_xx_x655_symbol : Boolean;
      signal assign_stmt_307_to_assign_stmt_319_x_xentry_x_xx_x656_symbol : Boolean;
      signal assign_stmt_307_to_assign_stmt_319_x_xexit_x_xx_x657_symbol : Boolean;
      signal bb_6_bb_7_658_symbol : Boolean;
      signal merge_stmt_321_x_xexit_x_xx_x659_symbol : Boolean;
      signal assign_stmt_325_to_assign_stmt_334_x_xentry_x_xx_x660_symbol : Boolean;
      signal assign_stmt_325_to_assign_stmt_334_x_xexit_x_xx_x661_symbol : Boolean;
      signal assign_stmt_338_x_xentry_x_xx_x662_symbol : Boolean;
      signal assign_stmt_338_x_xexit_x_xx_x663_symbol : Boolean;
      signal bb_7_bb_4_664_symbol : Boolean;
      signal merge_stmt_340_x_xexit_x_xx_x665_symbol : Boolean;
      signal assign_stmt_344_to_assign_stmt_353_x_xentry_x_xx_x666_symbol : Boolean;
      signal assign_stmt_344_to_assign_stmt_353_x_xexit_x_xx_x667_symbol : Boolean;
      signal if_stmt_354_x_xentry_x_xx_x668_symbol : Boolean;
      signal if_stmt_354_x_xexit_x_xx_x669_symbol : Boolean;
      signal merge_stmt_360_x_xentry_x_xx_x670_symbol : Boolean;
      signal merge_stmt_360_x_xexit_x_xx_x671_symbol : Boolean;
      signal assign_stmt_365_x_xentry_x_xx_x672_symbol : Boolean;
      signal assign_stmt_365_x_xexit_x_xx_x673_symbol : Boolean;
      signal assign_stmt_369_x_xentry_x_xx_x674_symbol : Boolean;
      signal assign_stmt_369_x_xexit_x_xx_x675_symbol : Boolean;
      signal assign_stmt_373_to_assign_stmt_400_x_xentry_x_xx_x676_symbol : Boolean;
      signal assign_stmt_373_to_assign_stmt_400_x_xexit_x_xx_x677_symbol : Boolean;
      signal bb_9_bb_4_678_symbol : Boolean;
      signal assign_stmt_142_to_assign_stmt_158_679_symbol : Boolean;
      signal assign_stmt_164_to_assign_stmt_173_743_symbol : Boolean;
      signal if_stmt_174_dead_link_828_symbol : Boolean;
      signal if_stmt_174_eval_test_832_symbol : Boolean;
      signal simple_obj_ref_175_place_836_symbol : Boolean;
      signal if_stmt_174_if_link_837_symbol : Boolean;
      signal if_stmt_174_else_link_841_symbol : Boolean;
      signal bb_1_bb_2_845_symbol : Boolean;
      signal bb_1_bb_3_846_symbol : Boolean;
      signal assign_stmt_184_to_assign_stmt_225_847_symbol : Boolean;
      signal assign_stmt_233_to_assign_stmt_245_1320_symbol : Boolean;
      signal assign_stmt_252_1414_symbol : Boolean;
      signal assign_stmt_256_1417_symbol : Boolean;
      signal assign_stmt_260_to_assign_stmt_273_1435_symbol : Boolean;
      signal if_stmt_274_dead_link_1523_symbol : Boolean;
      signal if_stmt_274_eval_test_1527_symbol : Boolean;
      signal simple_obj_ref_275_place_1531_symbol : Boolean;
      signal if_stmt_274_if_link_1532_symbol : Boolean;
      signal if_stmt_274_else_link_1536_symbol : Boolean;
      signal bb_4_bb_5_1540_symbol : Boolean;
      signal bb_4_bb_8_1541_symbol : Boolean;
      signal assign_stmt_283_to_assign_stmt_297_1542_symbol : Boolean;
      signal if_stmt_298_dead_link_1688_symbol : Boolean;
      signal if_stmt_298_eval_test_1692_symbol : Boolean;
      signal simple_obj_ref_299_place_1696_symbol : Boolean;
      signal if_stmt_298_if_link_1697_symbol : Boolean;
      signal if_stmt_298_else_link_1701_symbol : Boolean;
      signal bb_5_bb_6_1705_symbol : Boolean;
      signal bb_5_bb_7_1706_symbol : Boolean;
      signal assign_stmt_307_to_assign_stmt_319_1707_symbol : Boolean;
      signal assign_stmt_325_to_assign_stmt_334_1897_symbol : Boolean;
      signal assign_stmt_338_1971_symbol : Boolean;
      signal assign_stmt_344_to_assign_stmt_353_1990_symbol : Boolean;
      signal if_stmt_354_dead_link_2046_symbol : Boolean;
      signal if_stmt_354_eval_test_2050_symbol : Boolean;
      signal simple_obj_ref_355_place_2054_symbol : Boolean;
      signal if_stmt_354_if_link_2055_symbol : Boolean;
      signal if_stmt_354_else_link_2059_symbol : Boolean;
      signal bb_8_bb_9_2063_symbol : Boolean;
      signal bb_8_bb_4_2064_symbol : Boolean;
      signal assign_stmt_365_2065_symbol : Boolean;
      signal assign_stmt_369_2068_symbol : Boolean;
      signal assign_stmt_373_to_assign_stmt_400_2086_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_2471_symbol : Boolean;
      signal bb_2_bb_1_PhiReq_2474_symbol : Boolean;
      signal merge_stmt_160_PhiReqMerge_2477_symbol : Boolean;
      signal merge_stmt_160_PhiAck_2478_symbol : Boolean;
      signal merge_stmt_180_dead_link_2482_symbol : Boolean;
      signal bb_1_bb_2_PhiReq_2486_symbol : Boolean;
      signal merge_stmt_180_PhiReqMerge_2489_symbol : Boolean;
      signal merge_stmt_180_PhiAck_2490_symbol : Boolean;
      signal bb_1_bb_3_PhiReq_2494_symbol : Boolean;
      signal merge_stmt_227_PhiReqMerge_2497_symbol : Boolean;
      signal merge_stmt_227_PhiAck_2498_symbol : Boolean;
      signal bb_3_bb_4_PhiReq_2502_symbol : Boolean;
      signal bb_7_bb_4_PhiReq_2505_symbol : Boolean;
      signal bb_8_bb_4_PhiReq_2508_symbol : Boolean;
      signal bb_9_bb_4_PhiReq_2511_symbol : Boolean;
      signal merge_stmt_247_PhiReqMerge_2514_symbol : Boolean;
      signal merge_stmt_247_PhiAck_2515_symbol : Boolean;
      signal merge_stmt_280_dead_link_2519_symbol : Boolean;
      signal bb_4_bb_5_PhiReq_2523_symbol : Boolean;
      signal merge_stmt_280_PhiReqMerge_2526_symbol : Boolean;
      signal merge_stmt_280_PhiAck_2527_symbol : Boolean;
      signal merge_stmt_304_dead_link_2531_symbol : Boolean;
      signal bb_5_bb_6_PhiReq_2535_symbol : Boolean;
      signal merge_stmt_304_PhiReqMerge_2538_symbol : Boolean;
      signal merge_stmt_304_PhiAck_2539_symbol : Boolean;
      signal bb_5_bb_7_PhiReq_2543_symbol : Boolean;
      signal bb_6_bb_7_PhiReq_2546_symbol : Boolean;
      signal merge_stmt_321_PhiReqMerge_2549_symbol : Boolean;
      signal merge_stmt_321_PhiAck_2550_symbol : Boolean;
      signal bb_4_bb_8_PhiReq_2554_symbol : Boolean;
      signal merge_stmt_340_PhiReqMerge_2557_symbol : Boolean;
      signal merge_stmt_340_PhiAck_2558_symbol : Boolean;
      signal merge_stmt_360_dead_link_2562_symbol : Boolean;
      signal bb_8_bb_9_PhiReq_2566_symbol : Boolean;
      signal merge_stmt_360_PhiReqMerge_2569_symbol : Boolean;
      signal merge_stmt_360_PhiAck_2570_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_134_617_start <= Xentry_615_symbol; -- control passed to block
      Xentry_618_symbol  <= branch_block_stmt_134_617_start; -- transition branch_block_stmt_134/$entry
      branch_block_stmt_134_x_xentry_x_xx_x620_symbol  <=  Xentry_618_symbol; -- place branch_block_stmt_134/branch_block_stmt_134__entry__ (optimized away) 
      branch_block_stmt_134_x_xexit_x_xx_x621_symbol  <=   false ; -- place branch_block_stmt_134/branch_block_stmt_134__exit__ (optimized away) 
      assign_stmt_142_to_assign_stmt_158_x_xentry_x_xx_x622_symbol  <=  branch_block_stmt_134_x_xentry_x_xx_x620_symbol; -- place branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158__entry__ (optimized away) 
      assign_stmt_142_to_assign_stmt_158_x_xexit_x_xx_x623_symbol  <=  assign_stmt_142_to_assign_stmt_158_679_symbol; -- place branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158__exit__ (optimized away) 
      bb_0_bb_1_624_symbol  <=  assign_stmt_142_to_assign_stmt_158_x_xexit_x_xx_x623_symbol; -- place branch_block_stmt_134/bb_0_bb_1 (optimized away) 
      merge_stmt_160_x_xexit_x_xx_x625_symbol  <=  merge_stmt_160_PhiAck_2478_symbol; -- place branch_block_stmt_134/merge_stmt_160__exit__ (optimized away) 
      assign_stmt_164_to_assign_stmt_173_x_xentry_x_xx_x626_symbol  <=  merge_stmt_160_x_xexit_x_xx_x625_symbol; -- place branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173__entry__ (optimized away) 
      assign_stmt_164_to_assign_stmt_173_x_xexit_x_xx_x627_symbol  <=  assign_stmt_164_to_assign_stmt_173_743_symbol; -- place branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173__exit__ (optimized away) 
      if_stmt_174_x_xentry_x_xx_x628_symbol  <=  assign_stmt_164_to_assign_stmt_173_x_xexit_x_xx_x627_symbol; -- place branch_block_stmt_134/if_stmt_174__entry__ (optimized away) 
      if_stmt_174_x_xexit_x_xx_x629_symbol  <=  if_stmt_174_dead_link_828_symbol; -- place branch_block_stmt_134/if_stmt_174__exit__ (optimized away) 
      merge_stmt_180_x_xentry_x_xx_x630_symbol  <=  if_stmt_174_x_xexit_x_xx_x629_symbol; -- place branch_block_stmt_134/merge_stmt_180__entry__ (optimized away) 
      merge_stmt_180_x_xexit_x_xx_x631_symbol  <=  merge_stmt_180_dead_link_2482_symbol or merge_stmt_180_PhiAck_2490_symbol; -- place branch_block_stmt_134/merge_stmt_180__exit__ (optimized away) 
      assign_stmt_184_to_assign_stmt_225_x_xentry_x_xx_x632_symbol  <=  merge_stmt_180_x_xexit_x_xx_x631_symbol; -- place branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225__entry__ (optimized away) 
      assign_stmt_184_to_assign_stmt_225_x_xexit_x_xx_x633_symbol  <=  assign_stmt_184_to_assign_stmt_225_847_symbol; -- place branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225__exit__ (optimized away) 
      bb_2_bb_1_634_symbol  <=  assign_stmt_184_to_assign_stmt_225_x_xexit_x_xx_x633_symbol; -- place branch_block_stmt_134/bb_2_bb_1 (optimized away) 
      merge_stmt_227_x_xexit_x_xx_x635_symbol  <=  merge_stmt_227_PhiAck_2498_symbol; -- place branch_block_stmt_134/merge_stmt_227__exit__ (optimized away) 
      assign_stmt_233_to_assign_stmt_245_x_xentry_x_xx_x636_symbol  <=  merge_stmt_227_x_xexit_x_xx_x635_symbol; -- place branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245__entry__ (optimized away) 
      assign_stmt_233_to_assign_stmt_245_x_xexit_x_xx_x637_symbol  <=  assign_stmt_233_to_assign_stmt_245_1320_symbol; -- place branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245__exit__ (optimized away) 
      bb_3_bb_4_638_symbol  <=  assign_stmt_233_to_assign_stmt_245_x_xexit_x_xx_x637_symbol; -- place branch_block_stmt_134/bb_3_bb_4 (optimized away) 
      merge_stmt_247_x_xexit_x_xx_x639_symbol  <=  merge_stmt_247_PhiAck_2515_symbol; -- place branch_block_stmt_134/merge_stmt_247__exit__ (optimized away) 
      assign_stmt_252_x_xentry_x_xx_x640_symbol  <=  merge_stmt_247_x_xexit_x_xx_x639_symbol; -- place branch_block_stmt_134/assign_stmt_252__entry__ (optimized away) 
      assign_stmt_252_x_xexit_x_xx_x641_symbol  <=  assign_stmt_252_1414_symbol; -- place branch_block_stmt_134/assign_stmt_252__exit__ (optimized away) 
      assign_stmt_256_x_xentry_x_xx_x642_symbol  <=  assign_stmt_252_x_xexit_x_xx_x641_symbol; -- place branch_block_stmt_134/assign_stmt_256__entry__ (optimized away) 
      assign_stmt_256_x_xexit_x_xx_x643_symbol  <=  assign_stmt_256_1417_symbol; -- place branch_block_stmt_134/assign_stmt_256__exit__ (optimized away) 
      assign_stmt_260_to_assign_stmt_273_x_xentry_x_xx_x644_symbol  <=  assign_stmt_256_x_xexit_x_xx_x643_symbol; -- place branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273__entry__ (optimized away) 
      assign_stmt_260_to_assign_stmt_273_x_xexit_x_xx_x645_symbol  <=  assign_stmt_260_to_assign_stmt_273_1435_symbol; -- place branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273__exit__ (optimized away) 
      if_stmt_274_x_xentry_x_xx_x646_symbol  <=  assign_stmt_260_to_assign_stmt_273_x_xexit_x_xx_x645_symbol; -- place branch_block_stmt_134/if_stmt_274__entry__ (optimized away) 
      if_stmt_274_x_xexit_x_xx_x647_symbol  <=  if_stmt_274_dead_link_1523_symbol; -- place branch_block_stmt_134/if_stmt_274__exit__ (optimized away) 
      merge_stmt_280_x_xentry_x_xx_x648_symbol  <=  if_stmt_274_x_xexit_x_xx_x647_symbol; -- place branch_block_stmt_134/merge_stmt_280__entry__ (optimized away) 
      merge_stmt_280_x_xexit_x_xx_x649_symbol  <=  merge_stmt_280_dead_link_2519_symbol or merge_stmt_280_PhiAck_2527_symbol; -- place branch_block_stmt_134/merge_stmt_280__exit__ (optimized away) 
      assign_stmt_283_to_assign_stmt_297_x_xentry_x_xx_x650_symbol  <=  merge_stmt_280_x_xexit_x_xx_x649_symbol; -- place branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297__entry__ (optimized away) 
      assign_stmt_283_to_assign_stmt_297_x_xexit_x_xx_x651_symbol  <=  assign_stmt_283_to_assign_stmt_297_1542_symbol; -- place branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297__exit__ (optimized away) 
      if_stmt_298_x_xentry_x_xx_x652_symbol  <=  assign_stmt_283_to_assign_stmt_297_x_xexit_x_xx_x651_symbol; -- place branch_block_stmt_134/if_stmt_298__entry__ (optimized away) 
      if_stmt_298_x_xexit_x_xx_x653_symbol  <=  if_stmt_298_dead_link_1688_symbol; -- place branch_block_stmt_134/if_stmt_298__exit__ (optimized away) 
      merge_stmt_304_x_xentry_x_xx_x654_symbol  <=  if_stmt_298_x_xexit_x_xx_x653_symbol; -- place branch_block_stmt_134/merge_stmt_304__entry__ (optimized away) 
      merge_stmt_304_x_xexit_x_xx_x655_symbol  <=  merge_stmt_304_dead_link_2531_symbol or merge_stmt_304_PhiAck_2539_symbol; -- place branch_block_stmt_134/merge_stmt_304__exit__ (optimized away) 
      assign_stmt_307_to_assign_stmt_319_x_xentry_x_xx_x656_symbol  <=  merge_stmt_304_x_xexit_x_xx_x655_symbol; -- place branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319__entry__ (optimized away) 
      assign_stmt_307_to_assign_stmt_319_x_xexit_x_xx_x657_symbol  <=  assign_stmt_307_to_assign_stmt_319_1707_symbol; -- place branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319__exit__ (optimized away) 
      bb_6_bb_7_658_symbol  <=  assign_stmt_307_to_assign_stmt_319_x_xexit_x_xx_x657_symbol; -- place branch_block_stmt_134/bb_6_bb_7 (optimized away) 
      merge_stmt_321_x_xexit_x_xx_x659_symbol  <=  merge_stmt_321_PhiAck_2550_symbol; -- place branch_block_stmt_134/merge_stmt_321__exit__ (optimized away) 
      assign_stmt_325_to_assign_stmt_334_x_xentry_x_xx_x660_symbol  <=  merge_stmt_321_x_xexit_x_xx_x659_symbol; -- place branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334__entry__ (optimized away) 
      assign_stmt_325_to_assign_stmt_334_x_xexit_x_xx_x661_symbol  <=  assign_stmt_325_to_assign_stmt_334_1897_symbol; -- place branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334__exit__ (optimized away) 
      assign_stmt_338_x_xentry_x_xx_x662_symbol  <=  assign_stmt_325_to_assign_stmt_334_x_xexit_x_xx_x661_symbol; -- place branch_block_stmt_134/assign_stmt_338__entry__ (optimized away) 
      assign_stmt_338_x_xexit_x_xx_x663_symbol  <=  assign_stmt_338_1971_symbol; -- place branch_block_stmt_134/assign_stmt_338__exit__ (optimized away) 
      bb_7_bb_4_664_symbol  <=  assign_stmt_338_x_xexit_x_xx_x663_symbol; -- place branch_block_stmt_134/bb_7_bb_4 (optimized away) 
      merge_stmt_340_x_xexit_x_xx_x665_symbol  <=  merge_stmt_340_PhiAck_2558_symbol; -- place branch_block_stmt_134/merge_stmt_340__exit__ (optimized away) 
      assign_stmt_344_to_assign_stmt_353_x_xentry_x_xx_x666_symbol  <=  merge_stmt_340_x_xexit_x_xx_x665_symbol; -- place branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353__entry__ (optimized away) 
      assign_stmt_344_to_assign_stmt_353_x_xexit_x_xx_x667_symbol  <=  assign_stmt_344_to_assign_stmt_353_1990_symbol; -- place branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353__exit__ (optimized away) 
      if_stmt_354_x_xentry_x_xx_x668_symbol  <=  assign_stmt_344_to_assign_stmt_353_x_xexit_x_xx_x667_symbol; -- place branch_block_stmt_134/if_stmt_354__entry__ (optimized away) 
      if_stmt_354_x_xexit_x_xx_x669_symbol  <=  if_stmt_354_dead_link_2046_symbol; -- place branch_block_stmt_134/if_stmt_354__exit__ (optimized away) 
      merge_stmt_360_x_xentry_x_xx_x670_symbol  <=  if_stmt_354_x_xexit_x_xx_x669_symbol; -- place branch_block_stmt_134/merge_stmt_360__entry__ (optimized away) 
      merge_stmt_360_x_xexit_x_xx_x671_symbol  <=  merge_stmt_360_dead_link_2562_symbol or merge_stmt_360_PhiAck_2570_symbol; -- place branch_block_stmt_134/merge_stmt_360__exit__ (optimized away) 
      assign_stmt_365_x_xentry_x_xx_x672_symbol  <=  merge_stmt_360_x_xexit_x_xx_x671_symbol; -- place branch_block_stmt_134/assign_stmt_365__entry__ (optimized away) 
      assign_stmt_365_x_xexit_x_xx_x673_symbol  <=  assign_stmt_365_2065_symbol; -- place branch_block_stmt_134/assign_stmt_365__exit__ (optimized away) 
      assign_stmt_369_x_xentry_x_xx_x674_symbol  <=  assign_stmt_365_x_xexit_x_xx_x673_symbol; -- place branch_block_stmt_134/assign_stmt_369__entry__ (optimized away) 
      assign_stmt_369_x_xexit_x_xx_x675_symbol  <=  assign_stmt_369_2068_symbol; -- place branch_block_stmt_134/assign_stmt_369__exit__ (optimized away) 
      assign_stmt_373_to_assign_stmt_400_x_xentry_x_xx_x676_symbol  <=  assign_stmt_369_x_xexit_x_xx_x675_symbol; -- place branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400__entry__ (optimized away) 
      assign_stmt_373_to_assign_stmt_400_x_xexit_x_xx_x677_symbol  <=  assign_stmt_373_to_assign_stmt_400_2086_symbol; -- place branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400__exit__ (optimized away) 
      bb_9_bb_4_678_symbol  <=  assign_stmt_373_to_assign_stmt_400_x_xexit_x_xx_x677_symbol; -- place branch_block_stmt_134/bb_9_bb_4 (optimized away) 
      assign_stmt_142_to_assign_stmt_158_679: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158 
        signal assign_stmt_142_to_assign_stmt_158_679_start: Boolean;
        signal Xentry_680_symbol: Boolean;
        signal Xexit_681_symbol: Boolean;
        signal assign_stmt_158_active_x_x682_symbol : Boolean;
        signal assign_stmt_158_completed_x_x683_symbol : Boolean;
        signal ptr_deref_156_trigger_x_x684_symbol : Boolean;
        signal ptr_deref_156_active_x_x685_symbol : Boolean;
        signal ptr_deref_156_base_address_calculated_686_symbol : Boolean;
        signal ptr_deref_156_root_address_calculated_687_symbol : Boolean;
        signal ptr_deref_156_word_address_calculated_688_symbol : Boolean;
        signal ptr_deref_156_request_689_symbol : Boolean;
        signal ptr_deref_156_complete_717_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_142_to_assign_stmt_158_679_start <= assign_stmt_142_to_assign_stmt_158_x_xentry_x_xx_x622_symbol; -- control passed to block
        Xentry_680_symbol  <= assign_stmt_142_to_assign_stmt_158_679_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/$entry
        assign_stmt_158_active_x_x682_symbol <= Xentry_680_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/assign_stmt_158_active_
        assign_stmt_158_completed_x_x683_symbol <= ptr_deref_156_complete_717_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/assign_stmt_158_completed_
        ptr_deref_156_trigger_x_x684_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_trigger_ 
          signal ptr_deref_156_trigger_x_x684_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_156_trigger_x_x684_predecessors(0) <= ptr_deref_156_word_address_calculated_688_symbol;
          ptr_deref_156_trigger_x_x684_predecessors(1) <= assign_stmt_158_active_x_x682_symbol;
          ptr_deref_156_trigger_x_x684_join: join -- 
            port map( -- 
              preds => ptr_deref_156_trigger_x_x684_predecessors,
              symbol_out => ptr_deref_156_trigger_x_x684_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_trigger_
        ptr_deref_156_active_x_x685_symbol <= ptr_deref_156_request_689_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_active_
        ptr_deref_156_base_address_calculated_686_symbol <= Xentry_680_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_base_address_calculated
        ptr_deref_156_root_address_calculated_687_symbol <= Xentry_680_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_root_address_calculated
        ptr_deref_156_word_address_calculated_688_symbol <= ptr_deref_156_root_address_calculated_687_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_word_address_calculated
        ptr_deref_156_request_689: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request 
          signal ptr_deref_156_request_689_start: Boolean;
          signal Xentry_690_symbol: Boolean;
          signal Xexit_691_symbol: Boolean;
          signal split_req_692_symbol : Boolean;
          signal split_ack_693_symbol : Boolean;
          signal word_access_694_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_156_request_689_start <= ptr_deref_156_trigger_x_x684_symbol; -- control passed to block
          Xentry_690_symbol  <= ptr_deref_156_request_689_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/$entry
          split_req_692_symbol <= Xentry_690_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/split_req
          ptr_deref_156_gather_scatter_req_0 <= split_req_692_symbol; -- link to DP
          split_ack_693_symbol <= ptr_deref_156_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/split_ack
          word_access_694: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access 
            signal word_access_694_start: Boolean;
            signal Xentry_695_symbol: Boolean;
            signal Xexit_696_symbol: Boolean;
            signal word_access_0_697_symbol : Boolean;
            signal word_access_1_702_symbol : Boolean;
            signal word_access_2_707_symbol : Boolean;
            signal word_access_3_712_symbol : Boolean;
            -- 
          begin -- 
            word_access_694_start <= split_ack_693_symbol; -- control passed to block
            Xentry_695_symbol  <= word_access_694_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/$entry
            word_access_0_697: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0 
              signal word_access_0_697_start: Boolean;
              signal Xentry_698_symbol: Boolean;
              signal Xexit_699_symbol: Boolean;
              signal rr_700_symbol : Boolean;
              signal ra_701_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_697_start <= Xentry_695_symbol; -- control passed to block
              Xentry_698_symbol  <= word_access_0_697_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/$entry
              rr_700_symbol <= Xentry_698_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/rr
              ptr_deref_156_store_0_req_0 <= rr_700_symbol; -- link to DP
              ra_701_symbol <= ptr_deref_156_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/ra
              Xexit_699_symbol <= ra_701_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/$exit
              word_access_0_697_symbol <= Xexit_699_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0
            word_access_1_702: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_1 
              signal word_access_1_702_start: Boolean;
              signal Xentry_703_symbol: Boolean;
              signal Xexit_704_symbol: Boolean;
              signal rr_705_symbol : Boolean;
              signal ra_706_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_702_start <= Xentry_695_symbol; -- control passed to block
              Xentry_703_symbol  <= word_access_1_702_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_1/$entry
              rr_705_symbol <= Xentry_703_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_1/rr
              ptr_deref_156_store_1_req_0 <= rr_705_symbol; -- link to DP
              ra_706_symbol <= ptr_deref_156_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_1/ra
              Xexit_704_symbol <= ra_706_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_1/$exit
              word_access_1_702_symbol <= Xexit_704_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_1
            word_access_2_707: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_2 
              signal word_access_2_707_start: Boolean;
              signal Xentry_708_symbol: Boolean;
              signal Xexit_709_symbol: Boolean;
              signal rr_710_symbol : Boolean;
              signal ra_711_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_707_start <= Xentry_695_symbol; -- control passed to block
              Xentry_708_symbol  <= word_access_2_707_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_2/$entry
              rr_710_symbol <= Xentry_708_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_2/rr
              ptr_deref_156_store_2_req_0 <= rr_710_symbol; -- link to DP
              ra_711_symbol <= ptr_deref_156_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_2/ra
              Xexit_709_symbol <= ra_711_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_2/$exit
              word_access_2_707_symbol <= Xexit_709_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_2
            word_access_3_712: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_3 
              signal word_access_3_712_start: Boolean;
              signal Xentry_713_symbol: Boolean;
              signal Xexit_714_symbol: Boolean;
              signal rr_715_symbol : Boolean;
              signal ra_716_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_712_start <= Xentry_695_symbol; -- control passed to block
              Xentry_713_symbol  <= word_access_3_712_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_3/$entry
              rr_715_symbol <= Xentry_713_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_3/rr
              ptr_deref_156_store_3_req_0 <= rr_715_symbol; -- link to DP
              ra_716_symbol <= ptr_deref_156_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_3/ra
              Xexit_714_symbol <= ra_716_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_3/$exit
              word_access_3_712_symbol <= Xexit_714_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_3
            Xexit_696_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/$exit 
              signal Xexit_696_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_696_predecessors(0) <= word_access_0_697_symbol;
              Xexit_696_predecessors(1) <= word_access_1_702_symbol;
              Xexit_696_predecessors(2) <= word_access_2_707_symbol;
              Xexit_696_predecessors(3) <= word_access_3_712_symbol;
              Xexit_696_join: join -- 
                port map( -- 
                  preds => Xexit_696_predecessors,
                  symbol_out => Xexit_696_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/$exit
            word_access_694_symbol <= Xexit_696_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access
          Xexit_691_symbol <= word_access_694_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/$exit
          ptr_deref_156_request_689_symbol <= Xexit_691_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request
        ptr_deref_156_complete_717: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete 
          signal ptr_deref_156_complete_717_start: Boolean;
          signal Xentry_718_symbol: Boolean;
          signal Xexit_719_symbol: Boolean;
          signal word_access_720_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_156_complete_717_start <= ptr_deref_156_active_x_x685_symbol; -- control passed to block
          Xentry_718_symbol  <= ptr_deref_156_complete_717_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/$entry
          word_access_720: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access 
            signal word_access_720_start: Boolean;
            signal Xentry_721_symbol: Boolean;
            signal Xexit_722_symbol: Boolean;
            signal word_access_0_723_symbol : Boolean;
            signal word_access_1_728_symbol : Boolean;
            signal word_access_2_733_symbol : Boolean;
            signal word_access_3_738_symbol : Boolean;
            -- 
          begin -- 
            word_access_720_start <= Xentry_718_symbol; -- control passed to block
            Xentry_721_symbol  <= word_access_720_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/$entry
            word_access_0_723: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0 
              signal word_access_0_723_start: Boolean;
              signal Xentry_724_symbol: Boolean;
              signal Xexit_725_symbol: Boolean;
              signal cr_726_symbol : Boolean;
              signal ca_727_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_723_start <= Xentry_721_symbol; -- control passed to block
              Xentry_724_symbol  <= word_access_0_723_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/$entry
              cr_726_symbol <= Xentry_724_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/cr
              ptr_deref_156_store_0_req_1 <= cr_726_symbol; -- link to DP
              ca_727_symbol <= ptr_deref_156_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/ca
              Xexit_725_symbol <= ca_727_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/$exit
              word_access_0_723_symbol <= Xexit_725_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0
            word_access_1_728: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_1 
              signal word_access_1_728_start: Boolean;
              signal Xentry_729_symbol: Boolean;
              signal Xexit_730_symbol: Boolean;
              signal cr_731_symbol : Boolean;
              signal ca_732_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_728_start <= Xentry_721_symbol; -- control passed to block
              Xentry_729_symbol  <= word_access_1_728_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_1/$entry
              cr_731_symbol <= Xentry_729_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_1/cr
              ptr_deref_156_store_1_req_1 <= cr_731_symbol; -- link to DP
              ca_732_symbol <= ptr_deref_156_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_1/ca
              Xexit_730_symbol <= ca_732_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_1/$exit
              word_access_1_728_symbol <= Xexit_730_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_1
            word_access_2_733: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_2 
              signal word_access_2_733_start: Boolean;
              signal Xentry_734_symbol: Boolean;
              signal Xexit_735_symbol: Boolean;
              signal cr_736_symbol : Boolean;
              signal ca_737_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_733_start <= Xentry_721_symbol; -- control passed to block
              Xentry_734_symbol  <= word_access_2_733_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_2/$entry
              cr_736_symbol <= Xentry_734_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_2/cr
              ptr_deref_156_store_2_req_1 <= cr_736_symbol; -- link to DP
              ca_737_symbol <= ptr_deref_156_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_2/ca
              Xexit_735_symbol <= ca_737_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_2/$exit
              word_access_2_733_symbol <= Xexit_735_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_2
            word_access_3_738: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_3 
              signal word_access_3_738_start: Boolean;
              signal Xentry_739_symbol: Boolean;
              signal Xexit_740_symbol: Boolean;
              signal cr_741_symbol : Boolean;
              signal ca_742_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_738_start <= Xentry_721_symbol; -- control passed to block
              Xentry_739_symbol  <= word_access_3_738_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_3/$entry
              cr_741_symbol <= Xentry_739_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_3/cr
              ptr_deref_156_store_3_req_1 <= cr_741_symbol; -- link to DP
              ca_742_symbol <= ptr_deref_156_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_3/ca
              Xexit_740_symbol <= ca_742_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_3/$exit
              word_access_3_738_symbol <= Xexit_740_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_3
            Xexit_722_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/$exit 
              signal Xexit_722_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_722_predecessors(0) <= word_access_0_723_symbol;
              Xexit_722_predecessors(1) <= word_access_1_728_symbol;
              Xexit_722_predecessors(2) <= word_access_2_733_symbol;
              Xexit_722_predecessors(3) <= word_access_3_738_symbol;
              Xexit_722_join: join -- 
                port map( -- 
                  preds => Xexit_722_predecessors,
                  symbol_out => Xexit_722_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/$exit
            word_access_720_symbol <= Xexit_722_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access
          Xexit_719_symbol <= word_access_720_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/$exit
          ptr_deref_156_complete_717_symbol <= Xexit_719_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete
        Xexit_681_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/$exit 
          signal Xexit_681_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_681_predecessors(0) <= assign_stmt_158_completed_x_x683_symbol;
          Xexit_681_predecessors(1) <= ptr_deref_156_base_address_calculated_686_symbol;
          Xexit_681_join: join -- 
            port map( -- 
              preds => Xexit_681_predecessors,
              symbol_out => Xexit_681_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/$exit
        assign_stmt_142_to_assign_stmt_158_679_symbol <= Xexit_681_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158
      assign_stmt_164_to_assign_stmt_173_743: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173 
        signal assign_stmt_164_to_assign_stmt_173_743_start: Boolean;
        signal Xentry_744_symbol: Boolean;
        signal Xexit_745_symbol: Boolean;
        signal assign_stmt_164_active_x_x746_symbol : Boolean;
        signal assign_stmt_164_completed_x_x747_symbol : Boolean;
        signal ptr_deref_163_trigger_x_x748_symbol : Boolean;
        signal ptr_deref_163_active_x_x749_symbol : Boolean;
        signal ptr_deref_163_base_address_calculated_750_symbol : Boolean;
        signal ptr_deref_163_root_address_calculated_751_symbol : Boolean;
        signal ptr_deref_163_word_address_calculated_752_symbol : Boolean;
        signal ptr_deref_163_request_753_symbol : Boolean;
        signal ptr_deref_163_complete_779_symbol : Boolean;
        signal assign_stmt_173_active_x_x807_symbol : Boolean;
        signal assign_stmt_173_completed_x_x808_symbol : Boolean;
        signal binary_171_active_x_x809_symbol : Boolean;
        signal binary_171_trigger_x_x810_symbol : Boolean;
        signal type_cast_168_active_x_x811_symbol : Boolean;
        signal type_cast_168_trigger_x_x812_symbol : Boolean;
        signal simple_obj_ref_167_complete_813_symbol : Boolean;
        signal type_cast_168_complete_814_symbol : Boolean;
        signal binary_171_complete_821_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_164_to_assign_stmt_173_743_start <= assign_stmt_164_to_assign_stmt_173_x_xentry_x_xx_x626_symbol; -- control passed to block
        Xentry_744_symbol  <= assign_stmt_164_to_assign_stmt_173_743_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/$entry
        assign_stmt_164_active_x_x746_symbol <= ptr_deref_163_complete_779_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_164_active_
        assign_stmt_164_completed_x_x747_symbol <= assign_stmt_164_active_x_x746_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_164_completed_
        ptr_deref_163_trigger_x_x748_symbol <= ptr_deref_163_word_address_calculated_752_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_trigger_
        ptr_deref_163_active_x_x749_symbol <= ptr_deref_163_request_753_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_active_
        ptr_deref_163_base_address_calculated_750_symbol <= Xentry_744_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_base_address_calculated
        ptr_deref_163_root_address_calculated_751_symbol <= Xentry_744_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_root_address_calculated
        ptr_deref_163_word_address_calculated_752_symbol <= ptr_deref_163_root_address_calculated_751_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_word_address_calculated
        ptr_deref_163_request_753: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request 
          signal ptr_deref_163_request_753_start: Boolean;
          signal Xentry_754_symbol: Boolean;
          signal Xexit_755_symbol: Boolean;
          signal word_access_756_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_163_request_753_start <= ptr_deref_163_trigger_x_x748_symbol; -- control passed to block
          Xentry_754_symbol  <= ptr_deref_163_request_753_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/$entry
          word_access_756: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access 
            signal word_access_756_start: Boolean;
            signal Xentry_757_symbol: Boolean;
            signal Xexit_758_symbol: Boolean;
            signal word_access_0_759_symbol : Boolean;
            signal word_access_1_764_symbol : Boolean;
            signal word_access_2_769_symbol : Boolean;
            signal word_access_3_774_symbol : Boolean;
            -- 
          begin -- 
            word_access_756_start <= Xentry_754_symbol; -- control passed to block
            Xentry_757_symbol  <= word_access_756_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/$entry
            word_access_0_759: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0 
              signal word_access_0_759_start: Boolean;
              signal Xentry_760_symbol: Boolean;
              signal Xexit_761_symbol: Boolean;
              signal rr_762_symbol : Boolean;
              signal ra_763_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_759_start <= Xentry_757_symbol; -- control passed to block
              Xentry_760_symbol  <= word_access_0_759_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/$entry
              rr_762_symbol <= Xentry_760_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/rr
              ptr_deref_163_load_0_req_0 <= rr_762_symbol; -- link to DP
              ra_763_symbol <= ptr_deref_163_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/ra
              Xexit_761_symbol <= ra_763_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/$exit
              word_access_0_759_symbol <= Xexit_761_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0
            word_access_1_764: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_1 
              signal word_access_1_764_start: Boolean;
              signal Xentry_765_symbol: Boolean;
              signal Xexit_766_symbol: Boolean;
              signal rr_767_symbol : Boolean;
              signal ra_768_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_764_start <= Xentry_757_symbol; -- control passed to block
              Xentry_765_symbol  <= word_access_1_764_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_1/$entry
              rr_767_symbol <= Xentry_765_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_1/rr
              ptr_deref_163_load_1_req_0 <= rr_767_symbol; -- link to DP
              ra_768_symbol <= ptr_deref_163_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_1/ra
              Xexit_766_symbol <= ra_768_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_1/$exit
              word_access_1_764_symbol <= Xexit_766_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_1
            word_access_2_769: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_2 
              signal word_access_2_769_start: Boolean;
              signal Xentry_770_symbol: Boolean;
              signal Xexit_771_symbol: Boolean;
              signal rr_772_symbol : Boolean;
              signal ra_773_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_769_start <= Xentry_757_symbol; -- control passed to block
              Xentry_770_symbol  <= word_access_2_769_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_2/$entry
              rr_772_symbol <= Xentry_770_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_2/rr
              ptr_deref_163_load_2_req_0 <= rr_772_symbol; -- link to DP
              ra_773_symbol <= ptr_deref_163_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_2/ra
              Xexit_771_symbol <= ra_773_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_2/$exit
              word_access_2_769_symbol <= Xexit_771_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_2
            word_access_3_774: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_3 
              signal word_access_3_774_start: Boolean;
              signal Xentry_775_symbol: Boolean;
              signal Xexit_776_symbol: Boolean;
              signal rr_777_symbol : Boolean;
              signal ra_778_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_774_start <= Xentry_757_symbol; -- control passed to block
              Xentry_775_symbol  <= word_access_3_774_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_3/$entry
              rr_777_symbol <= Xentry_775_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_3/rr
              ptr_deref_163_load_3_req_0 <= rr_777_symbol; -- link to DP
              ra_778_symbol <= ptr_deref_163_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_3/ra
              Xexit_776_symbol <= ra_778_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_3/$exit
              word_access_3_774_symbol <= Xexit_776_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_3
            Xexit_758_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/$exit 
              signal Xexit_758_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_758_predecessors(0) <= word_access_0_759_symbol;
              Xexit_758_predecessors(1) <= word_access_1_764_symbol;
              Xexit_758_predecessors(2) <= word_access_2_769_symbol;
              Xexit_758_predecessors(3) <= word_access_3_774_symbol;
              Xexit_758_join: join -- 
                port map( -- 
                  preds => Xexit_758_predecessors,
                  symbol_out => Xexit_758_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/$exit
            word_access_756_symbol <= Xexit_758_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access
          Xexit_755_symbol <= word_access_756_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/$exit
          ptr_deref_163_request_753_symbol <= Xexit_755_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request
        ptr_deref_163_complete_779: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete 
          signal ptr_deref_163_complete_779_start: Boolean;
          signal Xentry_780_symbol: Boolean;
          signal Xexit_781_symbol: Boolean;
          signal word_access_782_symbol : Boolean;
          signal merge_req_805_symbol : Boolean;
          signal merge_ack_806_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_163_complete_779_start <= ptr_deref_163_active_x_x749_symbol; -- control passed to block
          Xentry_780_symbol  <= ptr_deref_163_complete_779_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/$entry
          word_access_782: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access 
            signal word_access_782_start: Boolean;
            signal Xentry_783_symbol: Boolean;
            signal Xexit_784_symbol: Boolean;
            signal word_access_0_785_symbol : Boolean;
            signal word_access_1_790_symbol : Boolean;
            signal word_access_2_795_symbol : Boolean;
            signal word_access_3_800_symbol : Boolean;
            -- 
          begin -- 
            word_access_782_start <= Xentry_780_symbol; -- control passed to block
            Xentry_783_symbol  <= word_access_782_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/$entry
            word_access_0_785: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0 
              signal word_access_0_785_start: Boolean;
              signal Xentry_786_symbol: Boolean;
              signal Xexit_787_symbol: Boolean;
              signal cr_788_symbol : Boolean;
              signal ca_789_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_785_start <= Xentry_783_symbol; -- control passed to block
              Xentry_786_symbol  <= word_access_0_785_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/$entry
              cr_788_symbol <= Xentry_786_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/cr
              ptr_deref_163_load_0_req_1 <= cr_788_symbol; -- link to DP
              ca_789_symbol <= ptr_deref_163_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/ca
              Xexit_787_symbol <= ca_789_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/$exit
              word_access_0_785_symbol <= Xexit_787_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0
            word_access_1_790: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_1 
              signal word_access_1_790_start: Boolean;
              signal Xentry_791_symbol: Boolean;
              signal Xexit_792_symbol: Boolean;
              signal cr_793_symbol : Boolean;
              signal ca_794_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_790_start <= Xentry_783_symbol; -- control passed to block
              Xentry_791_symbol  <= word_access_1_790_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_1/$entry
              cr_793_symbol <= Xentry_791_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_1/cr
              ptr_deref_163_load_1_req_1 <= cr_793_symbol; -- link to DP
              ca_794_symbol <= ptr_deref_163_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_1/ca
              Xexit_792_symbol <= ca_794_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_1/$exit
              word_access_1_790_symbol <= Xexit_792_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_1
            word_access_2_795: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_2 
              signal word_access_2_795_start: Boolean;
              signal Xentry_796_symbol: Boolean;
              signal Xexit_797_symbol: Boolean;
              signal cr_798_symbol : Boolean;
              signal ca_799_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_795_start <= Xentry_783_symbol; -- control passed to block
              Xentry_796_symbol  <= word_access_2_795_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_2/$entry
              cr_798_symbol <= Xentry_796_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_2/cr
              ptr_deref_163_load_2_req_1 <= cr_798_symbol; -- link to DP
              ca_799_symbol <= ptr_deref_163_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_2/ca
              Xexit_797_symbol <= ca_799_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_2/$exit
              word_access_2_795_symbol <= Xexit_797_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_2
            word_access_3_800: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_3 
              signal word_access_3_800_start: Boolean;
              signal Xentry_801_symbol: Boolean;
              signal Xexit_802_symbol: Boolean;
              signal cr_803_symbol : Boolean;
              signal ca_804_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_800_start <= Xentry_783_symbol; -- control passed to block
              Xentry_801_symbol  <= word_access_3_800_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_3/$entry
              cr_803_symbol <= Xentry_801_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_3/cr
              ptr_deref_163_load_3_req_1 <= cr_803_symbol; -- link to DP
              ca_804_symbol <= ptr_deref_163_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_3/ca
              Xexit_802_symbol <= ca_804_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_3/$exit
              word_access_3_800_symbol <= Xexit_802_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_3
            Xexit_784_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/$exit 
              signal Xexit_784_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_784_predecessors(0) <= word_access_0_785_symbol;
              Xexit_784_predecessors(1) <= word_access_1_790_symbol;
              Xexit_784_predecessors(2) <= word_access_2_795_symbol;
              Xexit_784_predecessors(3) <= word_access_3_800_symbol;
              Xexit_784_join: join -- 
                port map( -- 
                  preds => Xexit_784_predecessors,
                  symbol_out => Xexit_784_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/$exit
            word_access_782_symbol <= Xexit_784_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access
          merge_req_805_symbol <= word_access_782_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/merge_req
          ptr_deref_163_gather_scatter_req_0 <= merge_req_805_symbol; -- link to DP
          merge_ack_806_symbol <= ptr_deref_163_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/merge_ack
          Xexit_781_symbol <= merge_ack_806_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/$exit
          ptr_deref_163_complete_779_symbol <= Xexit_781_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete
        assign_stmt_173_active_x_x807_symbol <= binary_171_complete_821_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_173_active_
        assign_stmt_173_completed_x_x808_symbol <= assign_stmt_173_active_x_x807_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_173_completed_
        binary_171_active_x_x809_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_active_ 
          signal binary_171_active_x_x809_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_171_active_x_x809_predecessors(0) <= binary_171_trigger_x_x810_symbol;
          binary_171_active_x_x809_predecessors(1) <= type_cast_168_complete_814_symbol;
          binary_171_active_x_x809_join: join -- 
            port map( -- 
              preds => binary_171_active_x_x809_predecessors,
              symbol_out => binary_171_active_x_x809_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_active_
        binary_171_trigger_x_x810_symbol <= Xentry_744_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_trigger_
        type_cast_168_active_x_x811_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_active_ 
          signal type_cast_168_active_x_x811_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_168_active_x_x811_predecessors(0) <= type_cast_168_trigger_x_x812_symbol;
          type_cast_168_active_x_x811_predecessors(1) <= simple_obj_ref_167_complete_813_symbol;
          type_cast_168_active_x_x811_join: join -- 
            port map( -- 
              preds => type_cast_168_active_x_x811_predecessors,
              symbol_out => type_cast_168_active_x_x811_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_active_
        type_cast_168_trigger_x_x812_symbol <= Xentry_744_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_trigger_
        simple_obj_ref_167_complete_813_symbol <= assign_stmt_164_completed_x_x747_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/simple_obj_ref_167_complete
        type_cast_168_complete_814: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete 
          signal type_cast_168_complete_814_start: Boolean;
          signal Xentry_815_symbol: Boolean;
          signal Xexit_816_symbol: Boolean;
          signal rr_817_symbol : Boolean;
          signal ra_818_symbol : Boolean;
          signal cr_819_symbol : Boolean;
          signal ca_820_symbol : Boolean;
          -- 
        begin -- 
          type_cast_168_complete_814_start <= type_cast_168_active_x_x811_symbol; -- control passed to block
          Xentry_815_symbol  <= type_cast_168_complete_814_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/$entry
          rr_817_symbol <= Xentry_815_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/rr
          type_cast_168_inst_req_0 <= rr_817_symbol; -- link to DP
          ra_818_symbol <= type_cast_168_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/ra
          cr_819_symbol <= ra_818_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/cr
          type_cast_168_inst_req_1 <= cr_819_symbol; -- link to DP
          ca_820_symbol <= type_cast_168_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/ca
          Xexit_816_symbol <= ca_820_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/$exit
          type_cast_168_complete_814_symbol <= Xexit_816_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete
        binary_171_complete_821: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete 
          signal binary_171_complete_821_start: Boolean;
          signal Xentry_822_symbol: Boolean;
          signal Xexit_823_symbol: Boolean;
          signal rr_824_symbol : Boolean;
          signal ra_825_symbol : Boolean;
          signal cr_826_symbol : Boolean;
          signal ca_827_symbol : Boolean;
          -- 
        begin -- 
          binary_171_complete_821_start <= binary_171_active_x_x809_symbol; -- control passed to block
          Xentry_822_symbol  <= binary_171_complete_821_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/$entry
          rr_824_symbol <= Xentry_822_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/rr
          binary_171_inst_req_0 <= rr_824_symbol; -- link to DP
          ra_825_symbol <= binary_171_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/ra
          cr_826_symbol <= ra_825_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/cr
          binary_171_inst_req_1 <= cr_826_symbol; -- link to DP
          ca_827_symbol <= binary_171_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/ca
          Xexit_823_symbol <= ca_827_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/$exit
          binary_171_complete_821_symbol <= Xexit_823_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete
        Xexit_745_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/$exit 
          signal Xexit_745_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_745_predecessors(0) <= ptr_deref_163_base_address_calculated_750_symbol;
          Xexit_745_predecessors(1) <= assign_stmt_173_completed_x_x808_symbol;
          Xexit_745_join: join -- 
            port map( -- 
              preds => Xexit_745_predecessors,
              symbol_out => Xexit_745_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/$exit
        assign_stmt_164_to_assign_stmt_173_743_symbol <= Xexit_745_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173
      if_stmt_174_dead_link_828: Block -- branch_block_stmt_134/if_stmt_174_dead_link 
        signal if_stmt_174_dead_link_828_start: Boolean;
        signal Xentry_829_symbol: Boolean;
        signal Xexit_830_symbol: Boolean;
        signal dead_transition_831_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_dead_link_828_start <= if_stmt_174_x_xentry_x_xx_x628_symbol; -- control passed to block
        Xentry_829_symbol  <= if_stmt_174_dead_link_828_start; -- transition branch_block_stmt_134/if_stmt_174_dead_link/$entry
        dead_transition_831_symbol <= false;
        Xexit_830_symbol <= dead_transition_831_symbol; -- transition branch_block_stmt_134/if_stmt_174_dead_link/$exit
        if_stmt_174_dead_link_828_symbol <= Xexit_830_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_dead_link
      if_stmt_174_eval_test_832: Block -- branch_block_stmt_134/if_stmt_174_eval_test 
        signal if_stmt_174_eval_test_832_start: Boolean;
        signal Xentry_833_symbol: Boolean;
        signal Xexit_834_symbol: Boolean;
        signal branch_req_835_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_eval_test_832_start <= if_stmt_174_x_xentry_x_xx_x628_symbol; -- control passed to block
        Xentry_833_symbol  <= if_stmt_174_eval_test_832_start; -- transition branch_block_stmt_134/if_stmt_174_eval_test/$entry
        branch_req_835_symbol <= Xentry_833_symbol; -- transition branch_block_stmt_134/if_stmt_174_eval_test/branch_req
        if_stmt_174_branch_req_0 <= branch_req_835_symbol; -- link to DP
        Xexit_834_symbol <= branch_req_835_symbol; -- transition branch_block_stmt_134/if_stmt_174_eval_test/$exit
        if_stmt_174_eval_test_832_symbol <= Xexit_834_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_eval_test
      simple_obj_ref_175_place_836_symbol  <=  if_stmt_174_eval_test_832_symbol; -- place branch_block_stmt_134/simple_obj_ref_175_place (optimized away) 
      if_stmt_174_if_link_837: Block -- branch_block_stmt_134/if_stmt_174_if_link 
        signal if_stmt_174_if_link_837_start: Boolean;
        signal Xentry_838_symbol: Boolean;
        signal Xexit_839_symbol: Boolean;
        signal if_choice_transition_840_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_if_link_837_start <= simple_obj_ref_175_place_836_symbol; -- control passed to block
        Xentry_838_symbol  <= if_stmt_174_if_link_837_start; -- transition branch_block_stmt_134/if_stmt_174_if_link/$entry
        if_choice_transition_840_symbol <= if_stmt_174_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_174_if_link/if_choice_transition
        Xexit_839_symbol <= if_choice_transition_840_symbol; -- transition branch_block_stmt_134/if_stmt_174_if_link/$exit
        if_stmt_174_if_link_837_symbol <= Xexit_839_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_if_link
      if_stmt_174_else_link_841: Block -- branch_block_stmt_134/if_stmt_174_else_link 
        signal if_stmt_174_else_link_841_start: Boolean;
        signal Xentry_842_symbol: Boolean;
        signal Xexit_843_symbol: Boolean;
        signal else_choice_transition_844_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_else_link_841_start <= simple_obj_ref_175_place_836_symbol; -- control passed to block
        Xentry_842_symbol  <= if_stmt_174_else_link_841_start; -- transition branch_block_stmt_134/if_stmt_174_else_link/$entry
        else_choice_transition_844_symbol <= if_stmt_174_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_174_else_link/else_choice_transition
        Xexit_843_symbol <= else_choice_transition_844_symbol; -- transition branch_block_stmt_134/if_stmt_174_else_link/$exit
        if_stmt_174_else_link_841_symbol <= Xexit_843_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_else_link
      bb_1_bb_2_845_symbol  <=  if_stmt_174_if_link_837_symbol; -- place branch_block_stmt_134/bb_1_bb_2 (optimized away) 
      bb_1_bb_3_846_symbol  <=  if_stmt_174_else_link_841_symbol; -- place branch_block_stmt_134/bb_1_bb_3 (optimized away) 
      assign_stmt_184_to_assign_stmt_225_847: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225 
        signal assign_stmt_184_to_assign_stmt_225_847_start: Boolean;
        signal Xentry_848_symbol: Boolean;
        signal Xexit_849_symbol: Boolean;
        signal assign_stmt_184_active_x_x850_symbol : Boolean;
        signal assign_stmt_184_completed_x_x851_symbol : Boolean;
        signal ptr_deref_183_trigger_x_x852_symbol : Boolean;
        signal ptr_deref_183_active_x_x853_symbol : Boolean;
        signal ptr_deref_183_base_address_calculated_854_symbol : Boolean;
        signal ptr_deref_183_root_address_calculated_855_symbol : Boolean;
        signal ptr_deref_183_word_address_calculated_856_symbol : Boolean;
        signal ptr_deref_183_request_857_symbol : Boolean;
        signal ptr_deref_183_complete_883_symbol : Boolean;
        signal assign_stmt_189_active_x_x911_symbol : Boolean;
        signal assign_stmt_189_completed_x_x912_symbol : Boolean;
        signal binary_188_active_x_x913_symbol : Boolean;
        signal binary_188_trigger_x_x914_symbol : Boolean;
        signal simple_obj_ref_186_complete_915_symbol : Boolean;
        signal binary_188_complete_916_symbol : Boolean;
        signal assign_stmt_194_active_x_x923_symbol : Boolean;
        signal assign_stmt_194_completed_x_x924_symbol : Boolean;
        signal addr_of_193_active_x_x925_symbol : Boolean;
        signal addr_of_193_trigger_x_x926_symbol : Boolean;
        signal array_obj_ref_192_root_address_calculated_927_symbol : Boolean;
        signal array_obj_ref_192_indices_scaled_928_symbol : Boolean;
        signal array_obj_ref_192_offset_calculated_929_symbol : Boolean;
        signal array_obj_ref_192_index_computed_0_930_symbol : Boolean;
        signal array_obj_ref_192_index_resized_0_931_symbol : Boolean;
        signal simple_obj_ref_191_complete_932_symbol : Boolean;
        signal array_obj_ref_192_index_resize_0_933_symbol : Boolean;
        signal array_obj_ref_192_index_scale_0_938_symbol : Boolean;
        signal array_obj_ref_192_add_indices_945_symbol : Boolean;
        signal array_obj_ref_192_base_plus_offset_950_symbol : Boolean;
        signal addr_of_193_complete_955_symbol : Boolean;
        signal assign_stmt_198_active_x_x960_symbol : Boolean;
        signal assign_stmt_198_completed_x_x961_symbol : Boolean;
        signal ptr_deref_197_trigger_x_x962_symbol : Boolean;
        signal ptr_deref_197_active_x_x963_symbol : Boolean;
        signal ptr_deref_197_base_address_calculated_964_symbol : Boolean;
        signal ptr_deref_197_root_address_calculated_965_symbol : Boolean;
        signal ptr_deref_197_word_address_calculated_966_symbol : Boolean;
        signal ptr_deref_197_request_967_symbol : Boolean;
        signal ptr_deref_197_complete_993_symbol : Boolean;
        signal assign_stmt_203_active_x_x1021_symbol : Boolean;
        signal assign_stmt_203_completed_x_x1022_symbol : Boolean;
        signal addr_of_202_active_x_x1023_symbol : Boolean;
        signal addr_of_202_trigger_x_x1024_symbol : Boolean;
        signal array_obj_ref_201_root_address_calculated_1025_symbol : Boolean;
        signal array_obj_ref_201_indices_scaled_1026_symbol : Boolean;
        signal array_obj_ref_201_offset_calculated_1027_symbol : Boolean;
        signal array_obj_ref_201_index_computed_0_1028_symbol : Boolean;
        signal array_obj_ref_201_index_resized_0_1029_symbol : Boolean;
        signal simple_obj_ref_200_complete_1030_symbol : Boolean;
        signal array_obj_ref_201_index_resize_0_1031_symbol : Boolean;
        signal array_obj_ref_201_index_scale_0_1036_symbol : Boolean;
        signal array_obj_ref_201_add_indices_1043_symbol : Boolean;
        signal array_obj_ref_201_base_plus_offset_1048_symbol : Boolean;
        signal addr_of_202_complete_1053_symbol : Boolean;
        signal assign_stmt_208_active_x_x1058_symbol : Boolean;
        signal assign_stmt_208_completed_x_x1059_symbol : Boolean;
        signal array_obj_ref_207_trigger_x_x1060_symbol : Boolean;
        signal array_obj_ref_207_active_x_x1061_symbol : Boolean;
        signal array_obj_ref_207_base_address_calculated_1062_symbol : Boolean;
        signal array_obj_ref_207_root_address_calculated_1063_symbol : Boolean;
        signal array_obj_ref_207_base_address_resized_1064_symbol : Boolean;
        signal array_obj_ref_207_base_addr_resize_1065_symbol : Boolean;
        signal array_obj_ref_207_base_plus_offset_1070_symbol : Boolean;
        signal array_obj_ref_207_complete_1075_symbol : Boolean;
        signal assign_stmt_212_active_x_x1080_symbol : Boolean;
        signal assign_stmt_212_completed_x_x1081_symbol : Boolean;
        signal simple_obj_ref_211_complete_1082_symbol : Boolean;
        signal ptr_deref_210_trigger_x_x1083_symbol : Boolean;
        signal ptr_deref_210_active_x_x1084_symbol : Boolean;
        signal ptr_deref_210_base_address_calculated_1085_symbol : Boolean;
        signal simple_obj_ref_209_complete_1086_symbol : Boolean;
        signal ptr_deref_210_root_address_calculated_1087_symbol : Boolean;
        signal ptr_deref_210_word_address_calculated_1088_symbol : Boolean;
        signal ptr_deref_210_base_address_resized_1089_symbol : Boolean;
        signal ptr_deref_210_base_addr_resize_1090_symbol : Boolean;
        signal ptr_deref_210_base_plus_offset_1095_symbol : Boolean;
        signal ptr_deref_210_word_addrgen_1100_symbol : Boolean;
        signal ptr_deref_210_request_1131_symbol : Boolean;
        signal ptr_deref_210_complete_1159_symbol : Boolean;
        signal assign_stmt_216_active_x_x1185_symbol : Boolean;
        signal assign_stmt_216_completed_x_x1186_symbol : Boolean;
        signal ptr_deref_215_trigger_x_x1187_symbol : Boolean;
        signal ptr_deref_215_active_x_x1188_symbol : Boolean;
        signal ptr_deref_215_base_address_calculated_1189_symbol : Boolean;
        signal ptr_deref_215_root_address_calculated_1190_symbol : Boolean;
        signal ptr_deref_215_word_address_calculated_1191_symbol : Boolean;
        signal ptr_deref_215_request_1192_symbol : Boolean;
        signal ptr_deref_215_complete_1218_symbol : Boolean;
        signal assign_stmt_221_active_x_x1246_symbol : Boolean;
        signal assign_stmt_221_completed_x_x1247_symbol : Boolean;
        signal binary_220_active_x_x1248_symbol : Boolean;
        signal binary_220_trigger_x_x1249_symbol : Boolean;
        signal simple_obj_ref_218_complete_1250_symbol : Boolean;
        signal binary_220_complete_1251_symbol : Boolean;
        signal assign_stmt_225_active_x_x1258_symbol : Boolean;
        signal assign_stmt_225_completed_x_x1259_symbol : Boolean;
        signal simple_obj_ref_224_complete_1260_symbol : Boolean;
        signal ptr_deref_223_trigger_x_x1261_symbol : Boolean;
        signal ptr_deref_223_active_x_x1262_symbol : Boolean;
        signal ptr_deref_223_base_address_calculated_1263_symbol : Boolean;
        signal ptr_deref_223_root_address_calculated_1264_symbol : Boolean;
        signal ptr_deref_223_word_address_calculated_1265_symbol : Boolean;
        signal ptr_deref_223_request_1266_symbol : Boolean;
        signal ptr_deref_223_complete_1294_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_184_to_assign_stmt_225_847_start <= assign_stmt_184_to_assign_stmt_225_x_xentry_x_xx_x632_symbol; -- control passed to block
        Xentry_848_symbol  <= assign_stmt_184_to_assign_stmt_225_847_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/$entry
        assign_stmt_184_active_x_x850_symbol <= ptr_deref_183_complete_883_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_184_active_
        assign_stmt_184_completed_x_x851_symbol <= assign_stmt_184_active_x_x850_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_184_completed_
        ptr_deref_183_trigger_x_x852_symbol <= ptr_deref_183_word_address_calculated_856_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_trigger_
        ptr_deref_183_active_x_x853_symbol <= ptr_deref_183_request_857_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_active_
        ptr_deref_183_base_address_calculated_854_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_base_address_calculated
        ptr_deref_183_root_address_calculated_855_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_root_address_calculated
        ptr_deref_183_word_address_calculated_856_symbol <= ptr_deref_183_root_address_calculated_855_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_word_address_calculated
        ptr_deref_183_request_857: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request 
          signal ptr_deref_183_request_857_start: Boolean;
          signal Xentry_858_symbol: Boolean;
          signal Xexit_859_symbol: Boolean;
          signal word_access_860_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_183_request_857_start <= ptr_deref_183_trigger_x_x852_symbol; -- control passed to block
          Xentry_858_symbol  <= ptr_deref_183_request_857_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/$entry
          word_access_860: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access 
            signal word_access_860_start: Boolean;
            signal Xentry_861_symbol: Boolean;
            signal Xexit_862_symbol: Boolean;
            signal word_access_0_863_symbol : Boolean;
            signal word_access_1_868_symbol : Boolean;
            signal word_access_2_873_symbol : Boolean;
            signal word_access_3_878_symbol : Boolean;
            -- 
          begin -- 
            word_access_860_start <= Xentry_858_symbol; -- control passed to block
            Xentry_861_symbol  <= word_access_860_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/$entry
            word_access_0_863: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0 
              signal word_access_0_863_start: Boolean;
              signal Xentry_864_symbol: Boolean;
              signal Xexit_865_symbol: Boolean;
              signal rr_866_symbol : Boolean;
              signal ra_867_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_863_start <= Xentry_861_symbol; -- control passed to block
              Xentry_864_symbol  <= word_access_0_863_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/$entry
              rr_866_symbol <= Xentry_864_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/rr
              ptr_deref_183_load_0_req_0 <= rr_866_symbol; -- link to DP
              ra_867_symbol <= ptr_deref_183_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/ra
              Xexit_865_symbol <= ra_867_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/$exit
              word_access_0_863_symbol <= Xexit_865_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0
            word_access_1_868: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_1 
              signal word_access_1_868_start: Boolean;
              signal Xentry_869_symbol: Boolean;
              signal Xexit_870_symbol: Boolean;
              signal rr_871_symbol : Boolean;
              signal ra_872_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_868_start <= Xentry_861_symbol; -- control passed to block
              Xentry_869_symbol  <= word_access_1_868_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_1/$entry
              rr_871_symbol <= Xentry_869_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_1/rr
              ptr_deref_183_load_1_req_0 <= rr_871_symbol; -- link to DP
              ra_872_symbol <= ptr_deref_183_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_1/ra
              Xexit_870_symbol <= ra_872_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_1/$exit
              word_access_1_868_symbol <= Xexit_870_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_1
            word_access_2_873: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_2 
              signal word_access_2_873_start: Boolean;
              signal Xentry_874_symbol: Boolean;
              signal Xexit_875_symbol: Boolean;
              signal rr_876_symbol : Boolean;
              signal ra_877_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_873_start <= Xentry_861_symbol; -- control passed to block
              Xentry_874_symbol  <= word_access_2_873_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_2/$entry
              rr_876_symbol <= Xentry_874_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_2/rr
              ptr_deref_183_load_2_req_0 <= rr_876_symbol; -- link to DP
              ra_877_symbol <= ptr_deref_183_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_2/ra
              Xexit_875_symbol <= ra_877_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_2/$exit
              word_access_2_873_symbol <= Xexit_875_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_2
            word_access_3_878: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_3 
              signal word_access_3_878_start: Boolean;
              signal Xentry_879_symbol: Boolean;
              signal Xexit_880_symbol: Boolean;
              signal rr_881_symbol : Boolean;
              signal ra_882_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_878_start <= Xentry_861_symbol; -- control passed to block
              Xentry_879_symbol  <= word_access_3_878_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_3/$entry
              rr_881_symbol <= Xentry_879_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_3/rr
              ptr_deref_183_load_3_req_0 <= rr_881_symbol; -- link to DP
              ra_882_symbol <= ptr_deref_183_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_3/ra
              Xexit_880_symbol <= ra_882_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_3/$exit
              word_access_3_878_symbol <= Xexit_880_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_3
            Xexit_862_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/$exit 
              signal Xexit_862_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_862_predecessors(0) <= word_access_0_863_symbol;
              Xexit_862_predecessors(1) <= word_access_1_868_symbol;
              Xexit_862_predecessors(2) <= word_access_2_873_symbol;
              Xexit_862_predecessors(3) <= word_access_3_878_symbol;
              Xexit_862_join: join -- 
                port map( -- 
                  preds => Xexit_862_predecessors,
                  symbol_out => Xexit_862_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/$exit
            word_access_860_symbol <= Xexit_862_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access
          Xexit_859_symbol <= word_access_860_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/$exit
          ptr_deref_183_request_857_symbol <= Xexit_859_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request
        ptr_deref_183_complete_883: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete 
          signal ptr_deref_183_complete_883_start: Boolean;
          signal Xentry_884_symbol: Boolean;
          signal Xexit_885_symbol: Boolean;
          signal word_access_886_symbol : Boolean;
          signal merge_req_909_symbol : Boolean;
          signal merge_ack_910_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_183_complete_883_start <= ptr_deref_183_active_x_x853_symbol; -- control passed to block
          Xentry_884_symbol  <= ptr_deref_183_complete_883_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/$entry
          word_access_886: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access 
            signal word_access_886_start: Boolean;
            signal Xentry_887_symbol: Boolean;
            signal Xexit_888_symbol: Boolean;
            signal word_access_0_889_symbol : Boolean;
            signal word_access_1_894_symbol : Boolean;
            signal word_access_2_899_symbol : Boolean;
            signal word_access_3_904_symbol : Boolean;
            -- 
          begin -- 
            word_access_886_start <= Xentry_884_symbol; -- control passed to block
            Xentry_887_symbol  <= word_access_886_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/$entry
            word_access_0_889: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0 
              signal word_access_0_889_start: Boolean;
              signal Xentry_890_symbol: Boolean;
              signal Xexit_891_symbol: Boolean;
              signal cr_892_symbol : Boolean;
              signal ca_893_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_889_start <= Xentry_887_symbol; -- control passed to block
              Xentry_890_symbol  <= word_access_0_889_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/$entry
              cr_892_symbol <= Xentry_890_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/cr
              ptr_deref_183_load_0_req_1 <= cr_892_symbol; -- link to DP
              ca_893_symbol <= ptr_deref_183_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/ca
              Xexit_891_symbol <= ca_893_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/$exit
              word_access_0_889_symbol <= Xexit_891_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0
            word_access_1_894: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_1 
              signal word_access_1_894_start: Boolean;
              signal Xentry_895_symbol: Boolean;
              signal Xexit_896_symbol: Boolean;
              signal cr_897_symbol : Boolean;
              signal ca_898_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_894_start <= Xentry_887_symbol; -- control passed to block
              Xentry_895_symbol  <= word_access_1_894_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_1/$entry
              cr_897_symbol <= Xentry_895_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_1/cr
              ptr_deref_183_load_1_req_1 <= cr_897_symbol; -- link to DP
              ca_898_symbol <= ptr_deref_183_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_1/ca
              Xexit_896_symbol <= ca_898_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_1/$exit
              word_access_1_894_symbol <= Xexit_896_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_1
            word_access_2_899: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_2 
              signal word_access_2_899_start: Boolean;
              signal Xentry_900_symbol: Boolean;
              signal Xexit_901_symbol: Boolean;
              signal cr_902_symbol : Boolean;
              signal ca_903_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_899_start <= Xentry_887_symbol; -- control passed to block
              Xentry_900_symbol  <= word_access_2_899_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_2/$entry
              cr_902_symbol <= Xentry_900_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_2/cr
              ptr_deref_183_load_2_req_1 <= cr_902_symbol; -- link to DP
              ca_903_symbol <= ptr_deref_183_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_2/ca
              Xexit_901_symbol <= ca_903_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_2/$exit
              word_access_2_899_symbol <= Xexit_901_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_2
            word_access_3_904: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_3 
              signal word_access_3_904_start: Boolean;
              signal Xentry_905_symbol: Boolean;
              signal Xexit_906_symbol: Boolean;
              signal cr_907_symbol : Boolean;
              signal ca_908_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_904_start <= Xentry_887_symbol; -- control passed to block
              Xentry_905_symbol  <= word_access_3_904_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_3/$entry
              cr_907_symbol <= Xentry_905_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_3/cr
              ptr_deref_183_load_3_req_1 <= cr_907_symbol; -- link to DP
              ca_908_symbol <= ptr_deref_183_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_3/ca
              Xexit_906_symbol <= ca_908_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_3/$exit
              word_access_3_904_symbol <= Xexit_906_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_3
            Xexit_888_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/$exit 
              signal Xexit_888_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_888_predecessors(0) <= word_access_0_889_symbol;
              Xexit_888_predecessors(1) <= word_access_1_894_symbol;
              Xexit_888_predecessors(2) <= word_access_2_899_symbol;
              Xexit_888_predecessors(3) <= word_access_3_904_symbol;
              Xexit_888_join: join -- 
                port map( -- 
                  preds => Xexit_888_predecessors,
                  symbol_out => Xexit_888_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/$exit
            word_access_886_symbol <= Xexit_888_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access
          merge_req_909_symbol <= word_access_886_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/merge_req
          ptr_deref_183_gather_scatter_req_0 <= merge_req_909_symbol; -- link to DP
          merge_ack_910_symbol <= ptr_deref_183_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/merge_ack
          Xexit_885_symbol <= merge_ack_910_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/$exit
          ptr_deref_183_complete_883_symbol <= Xexit_885_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete
        assign_stmt_189_active_x_x911_symbol <= binary_188_complete_916_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_189_active_
        assign_stmt_189_completed_x_x912_symbol <= assign_stmt_189_active_x_x911_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_189_completed_
        binary_188_active_x_x913_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_active_ 
          signal binary_188_active_x_x913_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_188_active_x_x913_predecessors(0) <= binary_188_trigger_x_x914_symbol;
          binary_188_active_x_x913_predecessors(1) <= simple_obj_ref_186_complete_915_symbol;
          binary_188_active_x_x913_join: join -- 
            port map( -- 
              preds => binary_188_active_x_x913_predecessors,
              symbol_out => binary_188_active_x_x913_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_active_
        binary_188_trigger_x_x914_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_trigger_
        simple_obj_ref_186_complete_915_symbol <= assign_stmt_184_completed_x_x851_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_186_complete
        binary_188_complete_916: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete 
          signal binary_188_complete_916_start: Boolean;
          signal Xentry_917_symbol: Boolean;
          signal Xexit_918_symbol: Boolean;
          signal rr_919_symbol : Boolean;
          signal ra_920_symbol : Boolean;
          signal cr_921_symbol : Boolean;
          signal ca_922_symbol : Boolean;
          -- 
        begin -- 
          binary_188_complete_916_start <= binary_188_active_x_x913_symbol; -- control passed to block
          Xentry_917_symbol  <= binary_188_complete_916_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/$entry
          rr_919_symbol <= Xentry_917_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/rr
          binary_188_inst_req_0 <= rr_919_symbol; -- link to DP
          ra_920_symbol <= binary_188_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/ra
          cr_921_symbol <= ra_920_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/cr
          binary_188_inst_req_1 <= cr_921_symbol; -- link to DP
          ca_922_symbol <= binary_188_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/ca
          Xexit_918_symbol <= ca_922_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/$exit
          binary_188_complete_916_symbol <= Xexit_918_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete
        assign_stmt_194_active_x_x923_symbol <= addr_of_193_complete_955_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_194_active_
        assign_stmt_194_completed_x_x924_symbol <= assign_stmt_194_active_x_x923_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_194_completed_
        addr_of_193_active_x_x925_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_active_ 
          signal addr_of_193_active_x_x925_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          addr_of_193_active_x_x925_predecessors(0) <= addr_of_193_trigger_x_x926_symbol;
          addr_of_193_active_x_x925_predecessors(1) <= array_obj_ref_192_root_address_calculated_927_symbol;
          addr_of_193_active_x_x925_join: join -- 
            port map( -- 
              preds => addr_of_193_active_x_x925_predecessors,
              symbol_out => addr_of_193_active_x_x925_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_active_
        addr_of_193_trigger_x_x926_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_trigger_
        array_obj_ref_192_root_address_calculated_927_symbol <= array_obj_ref_192_base_plus_offset_950_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_root_address_calculated
        array_obj_ref_192_indices_scaled_928_symbol <= array_obj_ref_192_index_scale_0_938_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_indices_scaled
        array_obj_ref_192_offset_calculated_929_symbol <= array_obj_ref_192_add_indices_945_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_offset_calculated
        array_obj_ref_192_index_computed_0_930_symbol <= simple_obj_ref_191_complete_932_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_computed_0
        array_obj_ref_192_index_resized_0_931_symbol <= array_obj_ref_192_index_resize_0_933_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resized_0
        simple_obj_ref_191_complete_932_symbol <= assign_stmt_189_completed_x_x912_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_191_complete
        array_obj_ref_192_index_resize_0_933: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0 
          signal array_obj_ref_192_index_resize_0_933_start: Boolean;
          signal Xentry_934_symbol: Boolean;
          signal Xexit_935_symbol: Boolean;
          signal index_resize_req_936_symbol : Boolean;
          signal index_resize_ack_937_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_index_resize_0_933_start <= array_obj_ref_192_index_computed_0_930_symbol; -- control passed to block
          Xentry_934_symbol  <= array_obj_ref_192_index_resize_0_933_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/$entry
          index_resize_req_936_symbol <= Xentry_934_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/index_resize_req
          array_obj_ref_192_index_0_resize_req_0 <= index_resize_req_936_symbol; -- link to DP
          index_resize_ack_937_symbol <= array_obj_ref_192_index_0_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/index_resize_ack
          Xexit_935_symbol <= index_resize_ack_937_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/$exit
          array_obj_ref_192_index_resize_0_933_symbol <= Xexit_935_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0
        array_obj_ref_192_index_scale_0_938: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0 
          signal array_obj_ref_192_index_scale_0_938_start: Boolean;
          signal Xentry_939_symbol: Boolean;
          signal Xexit_940_symbol: Boolean;
          signal scale_rr_941_symbol : Boolean;
          signal scale_ra_942_symbol : Boolean;
          signal scale_cr_943_symbol : Boolean;
          signal scale_ca_944_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_index_scale_0_938_start <= array_obj_ref_192_index_resized_0_931_symbol; -- control passed to block
          Xentry_939_symbol  <= array_obj_ref_192_index_scale_0_938_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/$entry
          scale_rr_941_symbol <= Xentry_939_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_rr
          array_obj_ref_192_index_0_scale_req_0 <= scale_rr_941_symbol; -- link to DP
          scale_ra_942_symbol <= array_obj_ref_192_index_0_scale_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_ra
          scale_cr_943_symbol <= scale_ra_942_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_cr
          array_obj_ref_192_index_0_scale_req_1 <= scale_cr_943_symbol; -- link to DP
          scale_ca_944_symbol <= array_obj_ref_192_index_0_scale_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_ca
          Xexit_940_symbol <= scale_ca_944_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/$exit
          array_obj_ref_192_index_scale_0_938_symbol <= Xexit_940_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0
        array_obj_ref_192_add_indices_945: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices 
          signal array_obj_ref_192_add_indices_945_start: Boolean;
          signal Xentry_946_symbol: Boolean;
          signal Xexit_947_symbol: Boolean;
          signal final_index_req_948_symbol : Boolean;
          signal final_index_ack_949_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_add_indices_945_start <= array_obj_ref_192_indices_scaled_928_symbol; -- control passed to block
          Xentry_946_symbol  <= array_obj_ref_192_add_indices_945_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/$entry
          final_index_req_948_symbol <= Xentry_946_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/final_index_req
          array_obj_ref_192_offset_inst_req_0 <= final_index_req_948_symbol; -- link to DP
          final_index_ack_949_symbol <= array_obj_ref_192_offset_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/final_index_ack
          Xexit_947_symbol <= final_index_ack_949_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/$exit
          array_obj_ref_192_add_indices_945_symbol <= Xexit_947_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices
        array_obj_ref_192_base_plus_offset_950: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset 
          signal array_obj_ref_192_base_plus_offset_950_start: Boolean;
          signal Xentry_951_symbol: Boolean;
          signal Xexit_952_symbol: Boolean;
          signal sum_rename_req_953_symbol : Boolean;
          signal sum_rename_ack_954_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_base_plus_offset_950_start <= array_obj_ref_192_offset_calculated_929_symbol; -- control passed to block
          Xentry_951_symbol  <= array_obj_ref_192_base_plus_offset_950_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/$entry
          sum_rename_req_953_symbol <= Xentry_951_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/sum_rename_req
          array_obj_ref_192_root_address_inst_req_0 <= sum_rename_req_953_symbol; -- link to DP
          sum_rename_ack_954_symbol <= array_obj_ref_192_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/sum_rename_ack
          Xexit_952_symbol <= sum_rename_ack_954_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/$exit
          array_obj_ref_192_base_plus_offset_950_symbol <= Xexit_952_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset
        addr_of_193_complete_955: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete 
          signal addr_of_193_complete_955_start: Boolean;
          signal Xentry_956_symbol: Boolean;
          signal Xexit_957_symbol: Boolean;
          signal final_reg_req_958_symbol : Boolean;
          signal final_reg_ack_959_symbol : Boolean;
          -- 
        begin -- 
          addr_of_193_complete_955_start <= addr_of_193_active_x_x925_symbol; -- control passed to block
          Xentry_956_symbol  <= addr_of_193_complete_955_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/$entry
          final_reg_req_958_symbol <= Xentry_956_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/final_reg_req
          addr_of_193_final_reg_req_0 <= final_reg_req_958_symbol; -- link to DP
          final_reg_ack_959_symbol <= addr_of_193_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/final_reg_ack
          Xexit_957_symbol <= final_reg_ack_959_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/$exit
          addr_of_193_complete_955_symbol <= Xexit_957_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete
        assign_stmt_198_active_x_x960_symbol <= ptr_deref_197_complete_993_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_198_active_
        assign_stmt_198_completed_x_x961_symbol <= assign_stmt_198_active_x_x960_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_198_completed_
        ptr_deref_197_trigger_x_x962_symbol <= ptr_deref_197_word_address_calculated_966_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_trigger_
        ptr_deref_197_active_x_x963_symbol <= ptr_deref_197_request_967_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_active_
        ptr_deref_197_base_address_calculated_964_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_base_address_calculated
        ptr_deref_197_root_address_calculated_965_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_root_address_calculated
        ptr_deref_197_word_address_calculated_966_symbol <= ptr_deref_197_root_address_calculated_965_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_word_address_calculated
        ptr_deref_197_request_967: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request 
          signal ptr_deref_197_request_967_start: Boolean;
          signal Xentry_968_symbol: Boolean;
          signal Xexit_969_symbol: Boolean;
          signal word_access_970_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_197_request_967_start <= ptr_deref_197_trigger_x_x962_symbol; -- control passed to block
          Xentry_968_symbol  <= ptr_deref_197_request_967_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/$entry
          word_access_970: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access 
            signal word_access_970_start: Boolean;
            signal Xentry_971_symbol: Boolean;
            signal Xexit_972_symbol: Boolean;
            signal word_access_0_973_symbol : Boolean;
            signal word_access_1_978_symbol : Boolean;
            signal word_access_2_983_symbol : Boolean;
            signal word_access_3_988_symbol : Boolean;
            -- 
          begin -- 
            word_access_970_start <= Xentry_968_symbol; -- control passed to block
            Xentry_971_symbol  <= word_access_970_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/$entry
            word_access_0_973: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0 
              signal word_access_0_973_start: Boolean;
              signal Xentry_974_symbol: Boolean;
              signal Xexit_975_symbol: Boolean;
              signal rr_976_symbol : Boolean;
              signal ra_977_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_973_start <= Xentry_971_symbol; -- control passed to block
              Xentry_974_symbol  <= word_access_0_973_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/$entry
              rr_976_symbol <= Xentry_974_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/rr
              ptr_deref_197_load_0_req_0 <= rr_976_symbol; -- link to DP
              ra_977_symbol <= ptr_deref_197_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/ra
              Xexit_975_symbol <= ra_977_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/$exit
              word_access_0_973_symbol <= Xexit_975_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0
            word_access_1_978: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_1 
              signal word_access_1_978_start: Boolean;
              signal Xentry_979_symbol: Boolean;
              signal Xexit_980_symbol: Boolean;
              signal rr_981_symbol : Boolean;
              signal ra_982_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_978_start <= Xentry_971_symbol; -- control passed to block
              Xentry_979_symbol  <= word_access_1_978_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_1/$entry
              rr_981_symbol <= Xentry_979_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_1/rr
              ptr_deref_197_load_1_req_0 <= rr_981_symbol; -- link to DP
              ra_982_symbol <= ptr_deref_197_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_1/ra
              Xexit_980_symbol <= ra_982_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_1/$exit
              word_access_1_978_symbol <= Xexit_980_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_1
            word_access_2_983: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_2 
              signal word_access_2_983_start: Boolean;
              signal Xentry_984_symbol: Boolean;
              signal Xexit_985_symbol: Boolean;
              signal rr_986_symbol : Boolean;
              signal ra_987_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_983_start <= Xentry_971_symbol; -- control passed to block
              Xentry_984_symbol  <= word_access_2_983_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_2/$entry
              rr_986_symbol <= Xentry_984_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_2/rr
              ptr_deref_197_load_2_req_0 <= rr_986_symbol; -- link to DP
              ra_987_symbol <= ptr_deref_197_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_2/ra
              Xexit_985_symbol <= ra_987_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_2/$exit
              word_access_2_983_symbol <= Xexit_985_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_2
            word_access_3_988: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_3 
              signal word_access_3_988_start: Boolean;
              signal Xentry_989_symbol: Boolean;
              signal Xexit_990_symbol: Boolean;
              signal rr_991_symbol : Boolean;
              signal ra_992_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_988_start <= Xentry_971_symbol; -- control passed to block
              Xentry_989_symbol  <= word_access_3_988_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_3/$entry
              rr_991_symbol <= Xentry_989_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_3/rr
              ptr_deref_197_load_3_req_0 <= rr_991_symbol; -- link to DP
              ra_992_symbol <= ptr_deref_197_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_3/ra
              Xexit_990_symbol <= ra_992_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_3/$exit
              word_access_3_988_symbol <= Xexit_990_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_3
            Xexit_972_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/$exit 
              signal Xexit_972_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_972_predecessors(0) <= word_access_0_973_symbol;
              Xexit_972_predecessors(1) <= word_access_1_978_symbol;
              Xexit_972_predecessors(2) <= word_access_2_983_symbol;
              Xexit_972_predecessors(3) <= word_access_3_988_symbol;
              Xexit_972_join: join -- 
                port map( -- 
                  preds => Xexit_972_predecessors,
                  symbol_out => Xexit_972_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/$exit
            word_access_970_symbol <= Xexit_972_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access
          Xexit_969_symbol <= word_access_970_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/$exit
          ptr_deref_197_request_967_symbol <= Xexit_969_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request
        ptr_deref_197_complete_993: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete 
          signal ptr_deref_197_complete_993_start: Boolean;
          signal Xentry_994_symbol: Boolean;
          signal Xexit_995_symbol: Boolean;
          signal word_access_996_symbol : Boolean;
          signal merge_req_1019_symbol : Boolean;
          signal merge_ack_1020_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_197_complete_993_start <= ptr_deref_197_active_x_x963_symbol; -- control passed to block
          Xentry_994_symbol  <= ptr_deref_197_complete_993_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/$entry
          word_access_996: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access 
            signal word_access_996_start: Boolean;
            signal Xentry_997_symbol: Boolean;
            signal Xexit_998_symbol: Boolean;
            signal word_access_0_999_symbol : Boolean;
            signal word_access_1_1004_symbol : Boolean;
            signal word_access_2_1009_symbol : Boolean;
            signal word_access_3_1014_symbol : Boolean;
            -- 
          begin -- 
            word_access_996_start <= Xentry_994_symbol; -- control passed to block
            Xentry_997_symbol  <= word_access_996_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/$entry
            word_access_0_999: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0 
              signal word_access_0_999_start: Boolean;
              signal Xentry_1000_symbol: Boolean;
              signal Xexit_1001_symbol: Boolean;
              signal cr_1002_symbol : Boolean;
              signal ca_1003_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_999_start <= Xentry_997_symbol; -- control passed to block
              Xentry_1000_symbol  <= word_access_0_999_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/$entry
              cr_1002_symbol <= Xentry_1000_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/cr
              ptr_deref_197_load_0_req_1 <= cr_1002_symbol; -- link to DP
              ca_1003_symbol <= ptr_deref_197_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/ca
              Xexit_1001_symbol <= ca_1003_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/$exit
              word_access_0_999_symbol <= Xexit_1001_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0
            word_access_1_1004: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_1 
              signal word_access_1_1004_start: Boolean;
              signal Xentry_1005_symbol: Boolean;
              signal Xexit_1006_symbol: Boolean;
              signal cr_1007_symbol : Boolean;
              signal ca_1008_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1004_start <= Xentry_997_symbol; -- control passed to block
              Xentry_1005_symbol  <= word_access_1_1004_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_1/$entry
              cr_1007_symbol <= Xentry_1005_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_1/cr
              ptr_deref_197_load_1_req_1 <= cr_1007_symbol; -- link to DP
              ca_1008_symbol <= ptr_deref_197_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_1/ca
              Xexit_1006_symbol <= ca_1008_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_1/$exit
              word_access_1_1004_symbol <= Xexit_1006_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_1
            word_access_2_1009: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_2 
              signal word_access_2_1009_start: Boolean;
              signal Xentry_1010_symbol: Boolean;
              signal Xexit_1011_symbol: Boolean;
              signal cr_1012_symbol : Boolean;
              signal ca_1013_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1009_start <= Xentry_997_symbol; -- control passed to block
              Xentry_1010_symbol  <= word_access_2_1009_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_2/$entry
              cr_1012_symbol <= Xentry_1010_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_2/cr
              ptr_deref_197_load_2_req_1 <= cr_1012_symbol; -- link to DP
              ca_1013_symbol <= ptr_deref_197_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_2/ca
              Xexit_1011_symbol <= ca_1013_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_2/$exit
              word_access_2_1009_symbol <= Xexit_1011_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_2
            word_access_3_1014: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_3 
              signal word_access_3_1014_start: Boolean;
              signal Xentry_1015_symbol: Boolean;
              signal Xexit_1016_symbol: Boolean;
              signal cr_1017_symbol : Boolean;
              signal ca_1018_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1014_start <= Xentry_997_symbol; -- control passed to block
              Xentry_1015_symbol  <= word_access_3_1014_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_3/$entry
              cr_1017_symbol <= Xentry_1015_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_3/cr
              ptr_deref_197_load_3_req_1 <= cr_1017_symbol; -- link to DP
              ca_1018_symbol <= ptr_deref_197_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_3/ca
              Xexit_1016_symbol <= ca_1018_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_3/$exit
              word_access_3_1014_symbol <= Xexit_1016_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_3
            Xexit_998_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/$exit 
              signal Xexit_998_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_998_predecessors(0) <= word_access_0_999_symbol;
              Xexit_998_predecessors(1) <= word_access_1_1004_symbol;
              Xexit_998_predecessors(2) <= word_access_2_1009_symbol;
              Xexit_998_predecessors(3) <= word_access_3_1014_symbol;
              Xexit_998_join: join -- 
                port map( -- 
                  preds => Xexit_998_predecessors,
                  symbol_out => Xexit_998_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/$exit
            word_access_996_symbol <= Xexit_998_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access
          merge_req_1019_symbol <= word_access_996_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/merge_req
          ptr_deref_197_gather_scatter_req_0 <= merge_req_1019_symbol; -- link to DP
          merge_ack_1020_symbol <= ptr_deref_197_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/merge_ack
          Xexit_995_symbol <= merge_ack_1020_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/$exit
          ptr_deref_197_complete_993_symbol <= Xexit_995_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete
        assign_stmt_203_active_x_x1021_symbol <= addr_of_202_complete_1053_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_203_active_
        assign_stmt_203_completed_x_x1022_symbol <= assign_stmt_203_active_x_x1021_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_203_completed_
        addr_of_202_active_x_x1023_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_active_ 
          signal addr_of_202_active_x_x1023_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          addr_of_202_active_x_x1023_predecessors(0) <= addr_of_202_trigger_x_x1024_symbol;
          addr_of_202_active_x_x1023_predecessors(1) <= array_obj_ref_201_root_address_calculated_1025_symbol;
          addr_of_202_active_x_x1023_join: join -- 
            port map( -- 
              preds => addr_of_202_active_x_x1023_predecessors,
              symbol_out => addr_of_202_active_x_x1023_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_active_
        addr_of_202_trigger_x_x1024_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_trigger_
        array_obj_ref_201_root_address_calculated_1025_symbol <= array_obj_ref_201_base_plus_offset_1048_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_root_address_calculated
        array_obj_ref_201_indices_scaled_1026_symbol <= array_obj_ref_201_index_scale_0_1036_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_indices_scaled
        array_obj_ref_201_offset_calculated_1027_symbol <= array_obj_ref_201_add_indices_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_offset_calculated
        array_obj_ref_201_index_computed_0_1028_symbol <= simple_obj_ref_200_complete_1030_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_computed_0
        array_obj_ref_201_index_resized_0_1029_symbol <= array_obj_ref_201_index_resize_0_1031_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resized_0
        simple_obj_ref_200_complete_1030_symbol <= assign_stmt_198_completed_x_x961_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_200_complete
        array_obj_ref_201_index_resize_0_1031: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0 
          signal array_obj_ref_201_index_resize_0_1031_start: Boolean;
          signal Xentry_1032_symbol: Boolean;
          signal Xexit_1033_symbol: Boolean;
          signal index_resize_req_1034_symbol : Boolean;
          signal index_resize_ack_1035_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_index_resize_0_1031_start <= array_obj_ref_201_index_computed_0_1028_symbol; -- control passed to block
          Xentry_1032_symbol  <= array_obj_ref_201_index_resize_0_1031_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/$entry
          index_resize_req_1034_symbol <= Xentry_1032_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/index_resize_req
          array_obj_ref_201_index_0_resize_req_0 <= index_resize_req_1034_symbol; -- link to DP
          index_resize_ack_1035_symbol <= array_obj_ref_201_index_0_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/index_resize_ack
          Xexit_1033_symbol <= index_resize_ack_1035_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/$exit
          array_obj_ref_201_index_resize_0_1031_symbol <= Xexit_1033_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0
        array_obj_ref_201_index_scale_0_1036: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0 
          signal array_obj_ref_201_index_scale_0_1036_start: Boolean;
          signal Xentry_1037_symbol: Boolean;
          signal Xexit_1038_symbol: Boolean;
          signal scale_rr_1039_symbol : Boolean;
          signal scale_ra_1040_symbol : Boolean;
          signal scale_cr_1041_symbol : Boolean;
          signal scale_ca_1042_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_index_scale_0_1036_start <= array_obj_ref_201_index_resized_0_1029_symbol; -- control passed to block
          Xentry_1037_symbol  <= array_obj_ref_201_index_scale_0_1036_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/$entry
          scale_rr_1039_symbol <= Xentry_1037_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_rr
          array_obj_ref_201_index_0_scale_req_0 <= scale_rr_1039_symbol; -- link to DP
          scale_ra_1040_symbol <= array_obj_ref_201_index_0_scale_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_ra
          scale_cr_1041_symbol <= scale_ra_1040_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_cr
          array_obj_ref_201_index_0_scale_req_1 <= scale_cr_1041_symbol; -- link to DP
          scale_ca_1042_symbol <= array_obj_ref_201_index_0_scale_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_ca
          Xexit_1038_symbol <= scale_ca_1042_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/$exit
          array_obj_ref_201_index_scale_0_1036_symbol <= Xexit_1038_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0
        array_obj_ref_201_add_indices_1043: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices 
          signal array_obj_ref_201_add_indices_1043_start: Boolean;
          signal Xentry_1044_symbol: Boolean;
          signal Xexit_1045_symbol: Boolean;
          signal final_index_req_1046_symbol : Boolean;
          signal final_index_ack_1047_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_add_indices_1043_start <= array_obj_ref_201_indices_scaled_1026_symbol; -- control passed to block
          Xentry_1044_symbol  <= array_obj_ref_201_add_indices_1043_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/$entry
          final_index_req_1046_symbol <= Xentry_1044_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/final_index_req
          array_obj_ref_201_offset_inst_req_0 <= final_index_req_1046_symbol; -- link to DP
          final_index_ack_1047_symbol <= array_obj_ref_201_offset_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/final_index_ack
          Xexit_1045_symbol <= final_index_ack_1047_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/$exit
          array_obj_ref_201_add_indices_1043_symbol <= Xexit_1045_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices
        array_obj_ref_201_base_plus_offset_1048: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset 
          signal array_obj_ref_201_base_plus_offset_1048_start: Boolean;
          signal Xentry_1049_symbol: Boolean;
          signal Xexit_1050_symbol: Boolean;
          signal sum_rename_req_1051_symbol : Boolean;
          signal sum_rename_ack_1052_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_base_plus_offset_1048_start <= array_obj_ref_201_offset_calculated_1027_symbol; -- control passed to block
          Xentry_1049_symbol  <= array_obj_ref_201_base_plus_offset_1048_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/$entry
          sum_rename_req_1051_symbol <= Xentry_1049_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/sum_rename_req
          array_obj_ref_201_root_address_inst_req_0 <= sum_rename_req_1051_symbol; -- link to DP
          sum_rename_ack_1052_symbol <= array_obj_ref_201_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/sum_rename_ack
          Xexit_1050_symbol <= sum_rename_ack_1052_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/$exit
          array_obj_ref_201_base_plus_offset_1048_symbol <= Xexit_1050_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset
        addr_of_202_complete_1053: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete 
          signal addr_of_202_complete_1053_start: Boolean;
          signal Xentry_1054_symbol: Boolean;
          signal Xexit_1055_symbol: Boolean;
          signal final_reg_req_1056_symbol : Boolean;
          signal final_reg_ack_1057_symbol : Boolean;
          -- 
        begin -- 
          addr_of_202_complete_1053_start <= addr_of_202_active_x_x1023_symbol; -- control passed to block
          Xentry_1054_symbol  <= addr_of_202_complete_1053_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/$entry
          final_reg_req_1056_symbol <= Xentry_1054_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/final_reg_req
          addr_of_202_final_reg_req_0 <= final_reg_req_1056_symbol; -- link to DP
          final_reg_ack_1057_symbol <= addr_of_202_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/final_reg_ack
          Xexit_1055_symbol <= final_reg_ack_1057_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/$exit
          addr_of_202_complete_1053_symbol <= Xexit_1055_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete
        assign_stmt_208_active_x_x1058_symbol <= array_obj_ref_207_complete_1075_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_208_active_
        assign_stmt_208_completed_x_x1059_symbol <= assign_stmt_208_active_x_x1058_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_208_completed_
        array_obj_ref_207_trigger_x_x1060_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_trigger_
        array_obj_ref_207_active_x_x1061_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_active_ 
          signal array_obj_ref_207_active_x_x1061_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_207_active_x_x1061_predecessors(0) <= array_obj_ref_207_trigger_x_x1060_symbol;
          array_obj_ref_207_active_x_x1061_predecessors(1) <= array_obj_ref_207_root_address_calculated_1063_symbol;
          array_obj_ref_207_active_x_x1061_join: join -- 
            port map( -- 
              preds => array_obj_ref_207_active_x_x1061_predecessors,
              symbol_out => array_obj_ref_207_active_x_x1061_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_active_
        array_obj_ref_207_base_address_calculated_1062_symbol <= assign_stmt_203_completed_x_x1022_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_address_calculated
        array_obj_ref_207_root_address_calculated_1063_symbol <= array_obj_ref_207_base_plus_offset_1070_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_root_address_calculated
        array_obj_ref_207_base_address_resized_1064_symbol <= array_obj_ref_207_base_addr_resize_1065_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_address_resized
        array_obj_ref_207_base_addr_resize_1065: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize 
          signal array_obj_ref_207_base_addr_resize_1065_start: Boolean;
          signal Xentry_1066_symbol: Boolean;
          signal Xexit_1067_symbol: Boolean;
          signal base_resize_req_1068_symbol : Boolean;
          signal base_resize_ack_1069_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_207_base_addr_resize_1065_start <= array_obj_ref_207_base_address_calculated_1062_symbol; -- control passed to block
          Xentry_1066_symbol  <= array_obj_ref_207_base_addr_resize_1065_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/$entry
          base_resize_req_1068_symbol <= Xentry_1066_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/base_resize_req
          array_obj_ref_207_base_resize_req_0 <= base_resize_req_1068_symbol; -- link to DP
          base_resize_ack_1069_symbol <= array_obj_ref_207_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/base_resize_ack
          Xexit_1067_symbol <= base_resize_ack_1069_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/$exit
          array_obj_ref_207_base_addr_resize_1065_symbol <= Xexit_1067_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize
        array_obj_ref_207_base_plus_offset_1070: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset 
          signal array_obj_ref_207_base_plus_offset_1070_start: Boolean;
          signal Xentry_1071_symbol: Boolean;
          signal Xexit_1072_symbol: Boolean;
          signal sum_rename_req_1073_symbol : Boolean;
          signal sum_rename_ack_1074_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_207_base_plus_offset_1070_start <= array_obj_ref_207_base_address_resized_1064_symbol; -- control passed to block
          Xentry_1071_symbol  <= array_obj_ref_207_base_plus_offset_1070_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/$entry
          sum_rename_req_1073_symbol <= Xentry_1071_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/sum_rename_req
          array_obj_ref_207_root_address_inst_req_0 <= sum_rename_req_1073_symbol; -- link to DP
          sum_rename_ack_1074_symbol <= array_obj_ref_207_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/sum_rename_ack
          Xexit_1072_symbol <= sum_rename_ack_1074_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/$exit
          array_obj_ref_207_base_plus_offset_1070_symbol <= Xexit_1072_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset
        array_obj_ref_207_complete_1075: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete 
          signal array_obj_ref_207_complete_1075_start: Boolean;
          signal Xentry_1076_symbol: Boolean;
          signal Xexit_1077_symbol: Boolean;
          signal final_reg_req_1078_symbol : Boolean;
          signal final_reg_ack_1079_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_207_complete_1075_start <= array_obj_ref_207_active_x_x1061_symbol; -- control passed to block
          Xentry_1076_symbol  <= array_obj_ref_207_complete_1075_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/$entry
          final_reg_req_1078_symbol <= Xentry_1076_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/final_reg_req
          array_obj_ref_207_final_reg_req_0 <= final_reg_req_1078_symbol; -- link to DP
          final_reg_ack_1079_symbol <= array_obj_ref_207_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/final_reg_ack
          Xexit_1077_symbol <= final_reg_ack_1079_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/$exit
          array_obj_ref_207_complete_1075_symbol <= Xexit_1077_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete
        assign_stmt_212_active_x_x1080_symbol <= simple_obj_ref_211_complete_1082_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_212_active_
        assign_stmt_212_completed_x_x1081_symbol <= ptr_deref_210_complete_1159_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_212_completed_
        simple_obj_ref_211_complete_1082_symbol <= assign_stmt_194_completed_x_x924_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_211_complete
        ptr_deref_210_trigger_x_x1083_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_trigger_ 
          signal ptr_deref_210_trigger_x_x1083_predecessors: BooleanArray(4 downto 0);
          -- 
        begin -- 
          ptr_deref_210_trigger_x_x1083_predecessors(0) <= ptr_deref_210_word_address_calculated_1088_symbol;
          ptr_deref_210_trigger_x_x1083_predecessors(1) <= ptr_deref_210_base_address_calculated_1085_symbol;
          ptr_deref_210_trigger_x_x1083_predecessors(2) <= assign_stmt_212_active_x_x1080_symbol;
          ptr_deref_210_trigger_x_x1083_predecessors(3) <= ptr_deref_183_active_x_x853_symbol;
          ptr_deref_210_trigger_x_x1083_predecessors(4) <= ptr_deref_197_active_x_x963_symbol;
          ptr_deref_210_trigger_x_x1083_join: join -- 
            port map( -- 
              preds => ptr_deref_210_trigger_x_x1083_predecessors,
              symbol_out => ptr_deref_210_trigger_x_x1083_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_trigger_
        ptr_deref_210_active_x_x1084_symbol <= ptr_deref_210_request_1131_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_active_
        ptr_deref_210_base_address_calculated_1085_symbol <= simple_obj_ref_209_complete_1086_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_address_calculated
        simple_obj_ref_209_complete_1086_symbol <= assign_stmt_208_completed_x_x1059_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_209_complete
        ptr_deref_210_root_address_calculated_1087_symbol <= ptr_deref_210_base_plus_offset_1095_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_root_address_calculated
        ptr_deref_210_word_address_calculated_1088_symbol <= ptr_deref_210_word_addrgen_1100_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_address_calculated
        ptr_deref_210_base_address_resized_1089_symbol <= ptr_deref_210_base_addr_resize_1090_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_address_resized
        ptr_deref_210_base_addr_resize_1090: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize 
          signal ptr_deref_210_base_addr_resize_1090_start: Boolean;
          signal Xentry_1091_symbol: Boolean;
          signal Xexit_1092_symbol: Boolean;
          signal base_resize_req_1093_symbol : Boolean;
          signal base_resize_ack_1094_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_base_addr_resize_1090_start <= ptr_deref_210_base_address_calculated_1085_symbol; -- control passed to block
          Xentry_1091_symbol  <= ptr_deref_210_base_addr_resize_1090_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/$entry
          base_resize_req_1093_symbol <= Xentry_1091_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/base_resize_req
          ptr_deref_210_base_resize_req_0 <= base_resize_req_1093_symbol; -- link to DP
          base_resize_ack_1094_symbol <= ptr_deref_210_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/base_resize_ack
          Xexit_1092_symbol <= base_resize_ack_1094_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/$exit
          ptr_deref_210_base_addr_resize_1090_symbol <= Xexit_1092_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize
        ptr_deref_210_base_plus_offset_1095: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset 
          signal ptr_deref_210_base_plus_offset_1095_start: Boolean;
          signal Xentry_1096_symbol: Boolean;
          signal Xexit_1097_symbol: Boolean;
          signal sum_rename_req_1098_symbol : Boolean;
          signal sum_rename_ack_1099_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_base_plus_offset_1095_start <= ptr_deref_210_base_address_resized_1089_symbol; -- control passed to block
          Xentry_1096_symbol  <= ptr_deref_210_base_plus_offset_1095_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/$entry
          sum_rename_req_1098_symbol <= Xentry_1096_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/sum_rename_req
          ptr_deref_210_root_address_inst_req_0 <= sum_rename_req_1098_symbol; -- link to DP
          sum_rename_ack_1099_symbol <= ptr_deref_210_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/sum_rename_ack
          Xexit_1097_symbol <= sum_rename_ack_1099_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/$exit
          ptr_deref_210_base_plus_offset_1095_symbol <= Xexit_1097_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset
        ptr_deref_210_word_addrgen_1100: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen 
          signal ptr_deref_210_word_addrgen_1100_start: Boolean;
          signal Xentry_1101_symbol: Boolean;
          signal Xexit_1102_symbol: Boolean;
          signal word_0_1103_symbol : Boolean;
          signal word_1_1110_symbol : Boolean;
          signal word_2_1117_symbol : Boolean;
          signal word_3_1124_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_word_addrgen_1100_start <= ptr_deref_210_root_address_calculated_1087_symbol; -- control passed to block
          Xentry_1101_symbol  <= ptr_deref_210_word_addrgen_1100_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/$entry
          word_0_1103: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0 
            signal word_0_1103_start: Boolean;
            signal Xentry_1104_symbol: Boolean;
            signal Xexit_1105_symbol: Boolean;
            signal rr_1106_symbol : Boolean;
            signal ra_1107_symbol : Boolean;
            signal cr_1108_symbol : Boolean;
            signal ca_1109_symbol : Boolean;
            -- 
          begin -- 
            word_0_1103_start <= Xentry_1101_symbol; -- control passed to block
            Xentry_1104_symbol  <= word_0_1103_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0/$entry
            rr_1106_symbol <= Xentry_1104_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0/rr
            ptr_deref_210_addr_0_req_0 <= rr_1106_symbol; -- link to DP
            ra_1107_symbol <= ptr_deref_210_addr_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0/ra
            cr_1108_symbol <= ra_1107_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0/cr
            ptr_deref_210_addr_0_req_1 <= cr_1108_symbol; -- link to DP
            ca_1109_symbol <= ptr_deref_210_addr_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0/ca
            Xexit_1105_symbol <= ca_1109_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0/$exit
            word_0_1103_symbol <= Xexit_1105_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_0
          word_1_1110: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1 
            signal word_1_1110_start: Boolean;
            signal Xentry_1111_symbol: Boolean;
            signal Xexit_1112_symbol: Boolean;
            signal rr_1113_symbol : Boolean;
            signal ra_1114_symbol : Boolean;
            signal cr_1115_symbol : Boolean;
            signal ca_1116_symbol : Boolean;
            -- 
          begin -- 
            word_1_1110_start <= Xentry_1101_symbol; -- control passed to block
            Xentry_1111_symbol  <= word_1_1110_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1/$entry
            rr_1113_symbol <= Xentry_1111_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1/rr
            ptr_deref_210_addr_1_req_0 <= rr_1113_symbol; -- link to DP
            ra_1114_symbol <= ptr_deref_210_addr_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1/ra
            cr_1115_symbol <= ra_1114_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1/cr
            ptr_deref_210_addr_1_req_1 <= cr_1115_symbol; -- link to DP
            ca_1116_symbol <= ptr_deref_210_addr_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1/ca
            Xexit_1112_symbol <= ca_1116_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1/$exit
            word_1_1110_symbol <= Xexit_1112_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_1
          word_2_1117: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2 
            signal word_2_1117_start: Boolean;
            signal Xentry_1118_symbol: Boolean;
            signal Xexit_1119_symbol: Boolean;
            signal rr_1120_symbol : Boolean;
            signal ra_1121_symbol : Boolean;
            signal cr_1122_symbol : Boolean;
            signal ca_1123_symbol : Boolean;
            -- 
          begin -- 
            word_2_1117_start <= Xentry_1101_symbol; -- control passed to block
            Xentry_1118_symbol  <= word_2_1117_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2/$entry
            rr_1120_symbol <= Xentry_1118_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2/rr
            ptr_deref_210_addr_2_req_0 <= rr_1120_symbol; -- link to DP
            ra_1121_symbol <= ptr_deref_210_addr_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2/ra
            cr_1122_symbol <= ra_1121_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2/cr
            ptr_deref_210_addr_2_req_1 <= cr_1122_symbol; -- link to DP
            ca_1123_symbol <= ptr_deref_210_addr_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2/ca
            Xexit_1119_symbol <= ca_1123_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2/$exit
            word_2_1117_symbol <= Xexit_1119_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_2
          word_3_1124: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3 
            signal word_3_1124_start: Boolean;
            signal Xentry_1125_symbol: Boolean;
            signal Xexit_1126_symbol: Boolean;
            signal rr_1127_symbol : Boolean;
            signal ra_1128_symbol : Boolean;
            signal cr_1129_symbol : Boolean;
            signal ca_1130_symbol : Boolean;
            -- 
          begin -- 
            word_3_1124_start <= Xentry_1101_symbol; -- control passed to block
            Xentry_1125_symbol  <= word_3_1124_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3/$entry
            rr_1127_symbol <= Xentry_1125_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3/rr
            ptr_deref_210_addr_3_req_0 <= rr_1127_symbol; -- link to DP
            ra_1128_symbol <= ptr_deref_210_addr_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3/ra
            cr_1129_symbol <= ra_1128_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3/cr
            ptr_deref_210_addr_3_req_1 <= cr_1129_symbol; -- link to DP
            ca_1130_symbol <= ptr_deref_210_addr_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3/ca
            Xexit_1126_symbol <= ca_1130_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3/$exit
            word_3_1124_symbol <= Xexit_1126_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/word_3
          Xexit_1102_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/$exit 
            signal Xexit_1102_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_1102_predecessors(0) <= word_0_1103_symbol;
            Xexit_1102_predecessors(1) <= word_1_1110_symbol;
            Xexit_1102_predecessors(2) <= word_2_1117_symbol;
            Xexit_1102_predecessors(3) <= word_3_1124_symbol;
            Xexit_1102_join: join -- 
              port map( -- 
                preds => Xexit_1102_predecessors,
                symbol_out => Xexit_1102_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/$exit
          ptr_deref_210_word_addrgen_1100_symbol <= Xexit_1102_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen
        ptr_deref_210_request_1131: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request 
          signal ptr_deref_210_request_1131_start: Boolean;
          signal Xentry_1132_symbol: Boolean;
          signal Xexit_1133_symbol: Boolean;
          signal split_req_1134_symbol : Boolean;
          signal split_ack_1135_symbol : Boolean;
          signal word_access_1136_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_request_1131_start <= ptr_deref_210_trigger_x_x1083_symbol; -- control passed to block
          Xentry_1132_symbol  <= ptr_deref_210_request_1131_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/$entry
          split_req_1134_symbol <= Xentry_1132_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/split_req
          ptr_deref_210_gather_scatter_req_0 <= split_req_1134_symbol; -- link to DP
          split_ack_1135_symbol <= ptr_deref_210_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/split_ack
          word_access_1136: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access 
            signal word_access_1136_start: Boolean;
            signal Xentry_1137_symbol: Boolean;
            signal Xexit_1138_symbol: Boolean;
            signal word_access_0_1139_symbol : Boolean;
            signal word_access_1_1144_symbol : Boolean;
            signal word_access_2_1149_symbol : Boolean;
            signal word_access_3_1154_symbol : Boolean;
            -- 
          begin -- 
            word_access_1136_start <= split_ack_1135_symbol; -- control passed to block
            Xentry_1137_symbol  <= word_access_1136_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/$entry
            word_access_0_1139: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0 
              signal word_access_0_1139_start: Boolean;
              signal Xentry_1140_symbol: Boolean;
              signal Xexit_1141_symbol: Boolean;
              signal rr_1142_symbol : Boolean;
              signal ra_1143_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1139_start <= Xentry_1137_symbol; -- control passed to block
              Xentry_1140_symbol  <= word_access_0_1139_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/$entry
              rr_1142_symbol <= Xentry_1140_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/rr
              ptr_deref_210_store_0_req_0 <= rr_1142_symbol; -- link to DP
              ra_1143_symbol <= ptr_deref_210_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/ra
              Xexit_1141_symbol <= ra_1143_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/$exit
              word_access_0_1139_symbol <= Xexit_1141_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0
            word_access_1_1144: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_1 
              signal word_access_1_1144_start: Boolean;
              signal Xentry_1145_symbol: Boolean;
              signal Xexit_1146_symbol: Boolean;
              signal rr_1147_symbol : Boolean;
              signal ra_1148_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1144_start <= Xentry_1137_symbol; -- control passed to block
              Xentry_1145_symbol  <= word_access_1_1144_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_1/$entry
              rr_1147_symbol <= Xentry_1145_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_1/rr
              ptr_deref_210_store_1_req_0 <= rr_1147_symbol; -- link to DP
              ra_1148_symbol <= ptr_deref_210_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_1/ra
              Xexit_1146_symbol <= ra_1148_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_1/$exit
              word_access_1_1144_symbol <= Xexit_1146_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_1
            word_access_2_1149: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_2 
              signal word_access_2_1149_start: Boolean;
              signal Xentry_1150_symbol: Boolean;
              signal Xexit_1151_symbol: Boolean;
              signal rr_1152_symbol : Boolean;
              signal ra_1153_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1149_start <= Xentry_1137_symbol; -- control passed to block
              Xentry_1150_symbol  <= word_access_2_1149_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_2/$entry
              rr_1152_symbol <= Xentry_1150_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_2/rr
              ptr_deref_210_store_2_req_0 <= rr_1152_symbol; -- link to DP
              ra_1153_symbol <= ptr_deref_210_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_2/ra
              Xexit_1151_symbol <= ra_1153_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_2/$exit
              word_access_2_1149_symbol <= Xexit_1151_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_2
            word_access_3_1154: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_3 
              signal word_access_3_1154_start: Boolean;
              signal Xentry_1155_symbol: Boolean;
              signal Xexit_1156_symbol: Boolean;
              signal rr_1157_symbol : Boolean;
              signal ra_1158_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1154_start <= Xentry_1137_symbol; -- control passed to block
              Xentry_1155_symbol  <= word_access_3_1154_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_3/$entry
              rr_1157_symbol <= Xentry_1155_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_3/rr
              ptr_deref_210_store_3_req_0 <= rr_1157_symbol; -- link to DP
              ra_1158_symbol <= ptr_deref_210_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_3/ra
              Xexit_1156_symbol <= ra_1158_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_3/$exit
              word_access_3_1154_symbol <= Xexit_1156_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_3
            Xexit_1138_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/$exit 
              signal Xexit_1138_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1138_predecessors(0) <= word_access_0_1139_symbol;
              Xexit_1138_predecessors(1) <= word_access_1_1144_symbol;
              Xexit_1138_predecessors(2) <= word_access_2_1149_symbol;
              Xexit_1138_predecessors(3) <= word_access_3_1154_symbol;
              Xexit_1138_join: join -- 
                port map( -- 
                  preds => Xexit_1138_predecessors,
                  symbol_out => Xexit_1138_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/$exit
            word_access_1136_symbol <= Xexit_1138_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access
          Xexit_1133_symbol <= word_access_1136_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/$exit
          ptr_deref_210_request_1131_symbol <= Xexit_1133_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request
        ptr_deref_210_complete_1159: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete 
          signal ptr_deref_210_complete_1159_start: Boolean;
          signal Xentry_1160_symbol: Boolean;
          signal Xexit_1161_symbol: Boolean;
          signal word_access_1162_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_complete_1159_start <= ptr_deref_210_active_x_x1084_symbol; -- control passed to block
          Xentry_1160_symbol  <= ptr_deref_210_complete_1159_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/$entry
          word_access_1162: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access 
            signal word_access_1162_start: Boolean;
            signal Xentry_1163_symbol: Boolean;
            signal Xexit_1164_symbol: Boolean;
            signal word_access_0_1165_symbol : Boolean;
            signal word_access_1_1170_symbol : Boolean;
            signal word_access_2_1175_symbol : Boolean;
            signal word_access_3_1180_symbol : Boolean;
            -- 
          begin -- 
            word_access_1162_start <= Xentry_1160_symbol; -- control passed to block
            Xentry_1163_symbol  <= word_access_1162_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/$entry
            word_access_0_1165: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0 
              signal word_access_0_1165_start: Boolean;
              signal Xentry_1166_symbol: Boolean;
              signal Xexit_1167_symbol: Boolean;
              signal cr_1168_symbol : Boolean;
              signal ca_1169_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1165_start <= Xentry_1163_symbol; -- control passed to block
              Xentry_1166_symbol  <= word_access_0_1165_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/$entry
              cr_1168_symbol <= Xentry_1166_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/cr
              ptr_deref_210_store_0_req_1 <= cr_1168_symbol; -- link to DP
              ca_1169_symbol <= ptr_deref_210_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/ca
              Xexit_1167_symbol <= ca_1169_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/$exit
              word_access_0_1165_symbol <= Xexit_1167_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0
            word_access_1_1170: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_1 
              signal word_access_1_1170_start: Boolean;
              signal Xentry_1171_symbol: Boolean;
              signal Xexit_1172_symbol: Boolean;
              signal cr_1173_symbol : Boolean;
              signal ca_1174_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1170_start <= Xentry_1163_symbol; -- control passed to block
              Xentry_1171_symbol  <= word_access_1_1170_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_1/$entry
              cr_1173_symbol <= Xentry_1171_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_1/cr
              ptr_deref_210_store_1_req_1 <= cr_1173_symbol; -- link to DP
              ca_1174_symbol <= ptr_deref_210_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_1/ca
              Xexit_1172_symbol <= ca_1174_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_1/$exit
              word_access_1_1170_symbol <= Xexit_1172_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_1
            word_access_2_1175: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_2 
              signal word_access_2_1175_start: Boolean;
              signal Xentry_1176_symbol: Boolean;
              signal Xexit_1177_symbol: Boolean;
              signal cr_1178_symbol : Boolean;
              signal ca_1179_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1175_start <= Xentry_1163_symbol; -- control passed to block
              Xentry_1176_symbol  <= word_access_2_1175_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_2/$entry
              cr_1178_symbol <= Xentry_1176_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_2/cr
              ptr_deref_210_store_2_req_1 <= cr_1178_symbol; -- link to DP
              ca_1179_symbol <= ptr_deref_210_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_2/ca
              Xexit_1177_symbol <= ca_1179_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_2/$exit
              word_access_2_1175_symbol <= Xexit_1177_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_2
            word_access_3_1180: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_3 
              signal word_access_3_1180_start: Boolean;
              signal Xentry_1181_symbol: Boolean;
              signal Xexit_1182_symbol: Boolean;
              signal cr_1183_symbol : Boolean;
              signal ca_1184_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1180_start <= Xentry_1163_symbol; -- control passed to block
              Xentry_1181_symbol  <= word_access_3_1180_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_3/$entry
              cr_1183_symbol <= Xentry_1181_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_3/cr
              ptr_deref_210_store_3_req_1 <= cr_1183_symbol; -- link to DP
              ca_1184_symbol <= ptr_deref_210_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_3/ca
              Xexit_1182_symbol <= ca_1184_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_3/$exit
              word_access_3_1180_symbol <= Xexit_1182_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_3
            Xexit_1164_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/$exit 
              signal Xexit_1164_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1164_predecessors(0) <= word_access_0_1165_symbol;
              Xexit_1164_predecessors(1) <= word_access_1_1170_symbol;
              Xexit_1164_predecessors(2) <= word_access_2_1175_symbol;
              Xexit_1164_predecessors(3) <= word_access_3_1180_symbol;
              Xexit_1164_join: join -- 
                port map( -- 
                  preds => Xexit_1164_predecessors,
                  symbol_out => Xexit_1164_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/$exit
            word_access_1162_symbol <= Xexit_1164_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access
          Xexit_1161_symbol <= word_access_1162_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/$exit
          ptr_deref_210_complete_1159_symbol <= Xexit_1161_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete
        assign_stmt_216_active_x_x1185_symbol <= ptr_deref_215_complete_1218_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_216_active_
        assign_stmt_216_completed_x_x1186_symbol <= assign_stmt_216_active_x_x1185_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_216_completed_
        ptr_deref_215_trigger_x_x1187_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_trigger_ 
          signal ptr_deref_215_trigger_x_x1187_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_215_trigger_x_x1187_predecessors(0) <= ptr_deref_215_word_address_calculated_1191_symbol;
          ptr_deref_215_trigger_x_x1187_predecessors(1) <= ptr_deref_210_active_x_x1084_symbol;
          ptr_deref_215_trigger_x_x1187_join: join -- 
            port map( -- 
              preds => ptr_deref_215_trigger_x_x1187_predecessors,
              symbol_out => ptr_deref_215_trigger_x_x1187_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_trigger_
        ptr_deref_215_active_x_x1188_symbol <= ptr_deref_215_request_1192_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_active_
        ptr_deref_215_base_address_calculated_1189_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_base_address_calculated
        ptr_deref_215_root_address_calculated_1190_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_root_address_calculated
        ptr_deref_215_word_address_calculated_1191_symbol <= ptr_deref_215_root_address_calculated_1190_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_word_address_calculated
        ptr_deref_215_request_1192: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request 
          signal ptr_deref_215_request_1192_start: Boolean;
          signal Xentry_1193_symbol: Boolean;
          signal Xexit_1194_symbol: Boolean;
          signal word_access_1195_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_215_request_1192_start <= ptr_deref_215_trigger_x_x1187_symbol; -- control passed to block
          Xentry_1193_symbol  <= ptr_deref_215_request_1192_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/$entry
          word_access_1195: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access 
            signal word_access_1195_start: Boolean;
            signal Xentry_1196_symbol: Boolean;
            signal Xexit_1197_symbol: Boolean;
            signal word_access_0_1198_symbol : Boolean;
            signal word_access_1_1203_symbol : Boolean;
            signal word_access_2_1208_symbol : Boolean;
            signal word_access_3_1213_symbol : Boolean;
            -- 
          begin -- 
            word_access_1195_start <= Xentry_1193_symbol; -- control passed to block
            Xentry_1196_symbol  <= word_access_1195_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/$entry
            word_access_0_1198: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0 
              signal word_access_0_1198_start: Boolean;
              signal Xentry_1199_symbol: Boolean;
              signal Xexit_1200_symbol: Boolean;
              signal rr_1201_symbol : Boolean;
              signal ra_1202_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1198_start <= Xentry_1196_symbol; -- control passed to block
              Xentry_1199_symbol  <= word_access_0_1198_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/$entry
              rr_1201_symbol <= Xentry_1199_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/rr
              ptr_deref_215_load_0_req_0 <= rr_1201_symbol; -- link to DP
              ra_1202_symbol <= ptr_deref_215_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/ra
              Xexit_1200_symbol <= ra_1202_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/$exit
              word_access_0_1198_symbol <= Xexit_1200_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0
            word_access_1_1203: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_1 
              signal word_access_1_1203_start: Boolean;
              signal Xentry_1204_symbol: Boolean;
              signal Xexit_1205_symbol: Boolean;
              signal rr_1206_symbol : Boolean;
              signal ra_1207_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1203_start <= Xentry_1196_symbol; -- control passed to block
              Xentry_1204_symbol  <= word_access_1_1203_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_1/$entry
              rr_1206_symbol <= Xentry_1204_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_1/rr
              ptr_deref_215_load_1_req_0 <= rr_1206_symbol; -- link to DP
              ra_1207_symbol <= ptr_deref_215_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_1/ra
              Xexit_1205_symbol <= ra_1207_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_1/$exit
              word_access_1_1203_symbol <= Xexit_1205_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_1
            word_access_2_1208: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_2 
              signal word_access_2_1208_start: Boolean;
              signal Xentry_1209_symbol: Boolean;
              signal Xexit_1210_symbol: Boolean;
              signal rr_1211_symbol : Boolean;
              signal ra_1212_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1208_start <= Xentry_1196_symbol; -- control passed to block
              Xentry_1209_symbol  <= word_access_2_1208_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_2/$entry
              rr_1211_symbol <= Xentry_1209_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_2/rr
              ptr_deref_215_load_2_req_0 <= rr_1211_symbol; -- link to DP
              ra_1212_symbol <= ptr_deref_215_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_2/ra
              Xexit_1210_symbol <= ra_1212_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_2/$exit
              word_access_2_1208_symbol <= Xexit_1210_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_2
            word_access_3_1213: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_3 
              signal word_access_3_1213_start: Boolean;
              signal Xentry_1214_symbol: Boolean;
              signal Xexit_1215_symbol: Boolean;
              signal rr_1216_symbol : Boolean;
              signal ra_1217_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1213_start <= Xentry_1196_symbol; -- control passed to block
              Xentry_1214_symbol  <= word_access_3_1213_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_3/$entry
              rr_1216_symbol <= Xentry_1214_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_3/rr
              ptr_deref_215_load_3_req_0 <= rr_1216_symbol; -- link to DP
              ra_1217_symbol <= ptr_deref_215_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_3/ra
              Xexit_1215_symbol <= ra_1217_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_3/$exit
              word_access_3_1213_symbol <= Xexit_1215_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_3
            Xexit_1197_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/$exit 
              signal Xexit_1197_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1197_predecessors(0) <= word_access_0_1198_symbol;
              Xexit_1197_predecessors(1) <= word_access_1_1203_symbol;
              Xexit_1197_predecessors(2) <= word_access_2_1208_symbol;
              Xexit_1197_predecessors(3) <= word_access_3_1213_symbol;
              Xexit_1197_join: join -- 
                port map( -- 
                  preds => Xexit_1197_predecessors,
                  symbol_out => Xexit_1197_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/$exit
            word_access_1195_symbol <= Xexit_1197_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access
          Xexit_1194_symbol <= word_access_1195_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/$exit
          ptr_deref_215_request_1192_symbol <= Xexit_1194_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request
        ptr_deref_215_complete_1218: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete 
          signal ptr_deref_215_complete_1218_start: Boolean;
          signal Xentry_1219_symbol: Boolean;
          signal Xexit_1220_symbol: Boolean;
          signal word_access_1221_symbol : Boolean;
          signal merge_req_1244_symbol : Boolean;
          signal merge_ack_1245_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_215_complete_1218_start <= ptr_deref_215_active_x_x1188_symbol; -- control passed to block
          Xentry_1219_symbol  <= ptr_deref_215_complete_1218_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/$entry
          word_access_1221: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access 
            signal word_access_1221_start: Boolean;
            signal Xentry_1222_symbol: Boolean;
            signal Xexit_1223_symbol: Boolean;
            signal word_access_0_1224_symbol : Boolean;
            signal word_access_1_1229_symbol : Boolean;
            signal word_access_2_1234_symbol : Boolean;
            signal word_access_3_1239_symbol : Boolean;
            -- 
          begin -- 
            word_access_1221_start <= Xentry_1219_symbol; -- control passed to block
            Xentry_1222_symbol  <= word_access_1221_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/$entry
            word_access_0_1224: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0 
              signal word_access_0_1224_start: Boolean;
              signal Xentry_1225_symbol: Boolean;
              signal Xexit_1226_symbol: Boolean;
              signal cr_1227_symbol : Boolean;
              signal ca_1228_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1224_start <= Xentry_1222_symbol; -- control passed to block
              Xentry_1225_symbol  <= word_access_0_1224_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/$entry
              cr_1227_symbol <= Xentry_1225_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/cr
              ptr_deref_215_load_0_req_1 <= cr_1227_symbol; -- link to DP
              ca_1228_symbol <= ptr_deref_215_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/ca
              Xexit_1226_symbol <= ca_1228_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/$exit
              word_access_0_1224_symbol <= Xexit_1226_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0
            word_access_1_1229: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_1 
              signal word_access_1_1229_start: Boolean;
              signal Xentry_1230_symbol: Boolean;
              signal Xexit_1231_symbol: Boolean;
              signal cr_1232_symbol : Boolean;
              signal ca_1233_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1229_start <= Xentry_1222_symbol; -- control passed to block
              Xentry_1230_symbol  <= word_access_1_1229_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_1/$entry
              cr_1232_symbol <= Xentry_1230_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_1/cr
              ptr_deref_215_load_1_req_1 <= cr_1232_symbol; -- link to DP
              ca_1233_symbol <= ptr_deref_215_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_1/ca
              Xexit_1231_symbol <= ca_1233_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_1/$exit
              word_access_1_1229_symbol <= Xexit_1231_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_1
            word_access_2_1234: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_2 
              signal word_access_2_1234_start: Boolean;
              signal Xentry_1235_symbol: Boolean;
              signal Xexit_1236_symbol: Boolean;
              signal cr_1237_symbol : Boolean;
              signal ca_1238_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1234_start <= Xentry_1222_symbol; -- control passed to block
              Xentry_1235_symbol  <= word_access_2_1234_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_2/$entry
              cr_1237_symbol <= Xentry_1235_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_2/cr
              ptr_deref_215_load_2_req_1 <= cr_1237_symbol; -- link to DP
              ca_1238_symbol <= ptr_deref_215_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_2/ca
              Xexit_1236_symbol <= ca_1238_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_2/$exit
              word_access_2_1234_symbol <= Xexit_1236_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_2
            word_access_3_1239: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_3 
              signal word_access_3_1239_start: Boolean;
              signal Xentry_1240_symbol: Boolean;
              signal Xexit_1241_symbol: Boolean;
              signal cr_1242_symbol : Boolean;
              signal ca_1243_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1239_start <= Xentry_1222_symbol; -- control passed to block
              Xentry_1240_symbol  <= word_access_3_1239_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_3/$entry
              cr_1242_symbol <= Xentry_1240_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_3/cr
              ptr_deref_215_load_3_req_1 <= cr_1242_symbol; -- link to DP
              ca_1243_symbol <= ptr_deref_215_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_3/ca
              Xexit_1241_symbol <= ca_1243_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_3/$exit
              word_access_3_1239_symbol <= Xexit_1241_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_3
            Xexit_1223_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/$exit 
              signal Xexit_1223_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1223_predecessors(0) <= word_access_0_1224_symbol;
              Xexit_1223_predecessors(1) <= word_access_1_1229_symbol;
              Xexit_1223_predecessors(2) <= word_access_2_1234_symbol;
              Xexit_1223_predecessors(3) <= word_access_3_1239_symbol;
              Xexit_1223_join: join -- 
                port map( -- 
                  preds => Xexit_1223_predecessors,
                  symbol_out => Xexit_1223_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/$exit
            word_access_1221_symbol <= Xexit_1223_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access
          merge_req_1244_symbol <= word_access_1221_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/merge_req
          ptr_deref_215_gather_scatter_req_0 <= merge_req_1244_symbol; -- link to DP
          merge_ack_1245_symbol <= ptr_deref_215_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/merge_ack
          Xexit_1220_symbol <= merge_ack_1245_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/$exit
          ptr_deref_215_complete_1218_symbol <= Xexit_1220_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete
        assign_stmt_221_active_x_x1246_symbol <= binary_220_complete_1251_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_221_active_
        assign_stmt_221_completed_x_x1247_symbol <= assign_stmt_221_active_x_x1246_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_221_completed_
        binary_220_active_x_x1248_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_active_ 
          signal binary_220_active_x_x1248_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_220_active_x_x1248_predecessors(0) <= binary_220_trigger_x_x1249_symbol;
          binary_220_active_x_x1248_predecessors(1) <= simple_obj_ref_218_complete_1250_symbol;
          binary_220_active_x_x1248_join: join -- 
            port map( -- 
              preds => binary_220_active_x_x1248_predecessors,
              symbol_out => binary_220_active_x_x1248_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_active_
        binary_220_trigger_x_x1249_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_trigger_
        simple_obj_ref_218_complete_1250_symbol <= assign_stmt_216_completed_x_x1186_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_218_complete
        binary_220_complete_1251: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete 
          signal binary_220_complete_1251_start: Boolean;
          signal Xentry_1252_symbol: Boolean;
          signal Xexit_1253_symbol: Boolean;
          signal rr_1254_symbol : Boolean;
          signal ra_1255_symbol : Boolean;
          signal cr_1256_symbol : Boolean;
          signal ca_1257_symbol : Boolean;
          -- 
        begin -- 
          binary_220_complete_1251_start <= binary_220_active_x_x1248_symbol; -- control passed to block
          Xentry_1252_symbol  <= binary_220_complete_1251_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/$entry
          rr_1254_symbol <= Xentry_1252_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/rr
          binary_220_inst_req_0 <= rr_1254_symbol; -- link to DP
          ra_1255_symbol <= binary_220_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/ra
          cr_1256_symbol <= ra_1255_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/cr
          binary_220_inst_req_1 <= cr_1256_symbol; -- link to DP
          ca_1257_symbol <= binary_220_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/ca
          Xexit_1253_symbol <= ca_1257_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/$exit
          binary_220_complete_1251_symbol <= Xexit_1253_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete
        assign_stmt_225_active_x_x1258_symbol <= simple_obj_ref_224_complete_1260_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_225_active_
        assign_stmt_225_completed_x_x1259_symbol <= ptr_deref_223_complete_1294_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_225_completed_
        simple_obj_ref_224_complete_1260_symbol <= assign_stmt_221_completed_x_x1247_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_224_complete
        ptr_deref_223_trigger_x_x1261_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_trigger_ 
          signal ptr_deref_223_trigger_x_x1261_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          ptr_deref_223_trigger_x_x1261_predecessors(0) <= ptr_deref_223_word_address_calculated_1265_symbol;
          ptr_deref_223_trigger_x_x1261_predecessors(1) <= assign_stmt_225_active_x_x1258_symbol;
          ptr_deref_223_trigger_x_x1261_predecessors(2) <= ptr_deref_215_active_x_x1188_symbol;
          ptr_deref_223_trigger_x_x1261_join: join -- 
            port map( -- 
              preds => ptr_deref_223_trigger_x_x1261_predecessors,
              symbol_out => ptr_deref_223_trigger_x_x1261_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_trigger_
        ptr_deref_223_active_x_x1262_symbol <= ptr_deref_223_request_1266_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_active_
        ptr_deref_223_base_address_calculated_1263_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_base_address_calculated
        ptr_deref_223_root_address_calculated_1264_symbol <= Xentry_848_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_root_address_calculated
        ptr_deref_223_word_address_calculated_1265_symbol <= ptr_deref_223_root_address_calculated_1264_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_word_address_calculated
        ptr_deref_223_request_1266: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request 
          signal ptr_deref_223_request_1266_start: Boolean;
          signal Xentry_1267_symbol: Boolean;
          signal Xexit_1268_symbol: Boolean;
          signal split_req_1269_symbol : Boolean;
          signal split_ack_1270_symbol : Boolean;
          signal word_access_1271_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_223_request_1266_start <= ptr_deref_223_trigger_x_x1261_symbol; -- control passed to block
          Xentry_1267_symbol  <= ptr_deref_223_request_1266_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/$entry
          split_req_1269_symbol <= Xentry_1267_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/split_req
          ptr_deref_223_gather_scatter_req_0 <= split_req_1269_symbol; -- link to DP
          split_ack_1270_symbol <= ptr_deref_223_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/split_ack
          word_access_1271: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access 
            signal word_access_1271_start: Boolean;
            signal Xentry_1272_symbol: Boolean;
            signal Xexit_1273_symbol: Boolean;
            signal word_access_0_1274_symbol : Boolean;
            signal word_access_1_1279_symbol : Boolean;
            signal word_access_2_1284_symbol : Boolean;
            signal word_access_3_1289_symbol : Boolean;
            -- 
          begin -- 
            word_access_1271_start <= split_ack_1270_symbol; -- control passed to block
            Xentry_1272_symbol  <= word_access_1271_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/$entry
            word_access_0_1274: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0 
              signal word_access_0_1274_start: Boolean;
              signal Xentry_1275_symbol: Boolean;
              signal Xexit_1276_symbol: Boolean;
              signal rr_1277_symbol : Boolean;
              signal ra_1278_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1274_start <= Xentry_1272_symbol; -- control passed to block
              Xentry_1275_symbol  <= word_access_0_1274_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/$entry
              rr_1277_symbol <= Xentry_1275_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/rr
              ptr_deref_223_store_0_req_0 <= rr_1277_symbol; -- link to DP
              ra_1278_symbol <= ptr_deref_223_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/ra
              Xexit_1276_symbol <= ra_1278_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/$exit
              word_access_0_1274_symbol <= Xexit_1276_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0
            word_access_1_1279: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_1 
              signal word_access_1_1279_start: Boolean;
              signal Xentry_1280_symbol: Boolean;
              signal Xexit_1281_symbol: Boolean;
              signal rr_1282_symbol : Boolean;
              signal ra_1283_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1279_start <= Xentry_1272_symbol; -- control passed to block
              Xentry_1280_symbol  <= word_access_1_1279_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_1/$entry
              rr_1282_symbol <= Xentry_1280_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_1/rr
              ptr_deref_223_store_1_req_0 <= rr_1282_symbol; -- link to DP
              ra_1283_symbol <= ptr_deref_223_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_1/ra
              Xexit_1281_symbol <= ra_1283_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_1/$exit
              word_access_1_1279_symbol <= Xexit_1281_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_1
            word_access_2_1284: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_2 
              signal word_access_2_1284_start: Boolean;
              signal Xentry_1285_symbol: Boolean;
              signal Xexit_1286_symbol: Boolean;
              signal rr_1287_symbol : Boolean;
              signal ra_1288_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1284_start <= Xentry_1272_symbol; -- control passed to block
              Xentry_1285_symbol  <= word_access_2_1284_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_2/$entry
              rr_1287_symbol <= Xentry_1285_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_2/rr
              ptr_deref_223_store_2_req_0 <= rr_1287_symbol; -- link to DP
              ra_1288_symbol <= ptr_deref_223_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_2/ra
              Xexit_1286_symbol <= ra_1288_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_2/$exit
              word_access_2_1284_symbol <= Xexit_1286_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_2
            word_access_3_1289: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_3 
              signal word_access_3_1289_start: Boolean;
              signal Xentry_1290_symbol: Boolean;
              signal Xexit_1291_symbol: Boolean;
              signal rr_1292_symbol : Boolean;
              signal ra_1293_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1289_start <= Xentry_1272_symbol; -- control passed to block
              Xentry_1290_symbol  <= word_access_3_1289_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_3/$entry
              rr_1292_symbol <= Xentry_1290_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_3/rr
              ptr_deref_223_store_3_req_0 <= rr_1292_symbol; -- link to DP
              ra_1293_symbol <= ptr_deref_223_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_3/ra
              Xexit_1291_symbol <= ra_1293_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_3/$exit
              word_access_3_1289_symbol <= Xexit_1291_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_3
            Xexit_1273_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/$exit 
              signal Xexit_1273_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1273_predecessors(0) <= word_access_0_1274_symbol;
              Xexit_1273_predecessors(1) <= word_access_1_1279_symbol;
              Xexit_1273_predecessors(2) <= word_access_2_1284_symbol;
              Xexit_1273_predecessors(3) <= word_access_3_1289_symbol;
              Xexit_1273_join: join -- 
                port map( -- 
                  preds => Xexit_1273_predecessors,
                  symbol_out => Xexit_1273_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/$exit
            word_access_1271_symbol <= Xexit_1273_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access
          Xexit_1268_symbol <= word_access_1271_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/$exit
          ptr_deref_223_request_1266_symbol <= Xexit_1268_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request
        ptr_deref_223_complete_1294: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete 
          signal ptr_deref_223_complete_1294_start: Boolean;
          signal Xentry_1295_symbol: Boolean;
          signal Xexit_1296_symbol: Boolean;
          signal word_access_1297_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_223_complete_1294_start <= ptr_deref_223_active_x_x1262_symbol; -- control passed to block
          Xentry_1295_symbol  <= ptr_deref_223_complete_1294_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/$entry
          word_access_1297: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access 
            signal word_access_1297_start: Boolean;
            signal Xentry_1298_symbol: Boolean;
            signal Xexit_1299_symbol: Boolean;
            signal word_access_0_1300_symbol : Boolean;
            signal word_access_1_1305_symbol : Boolean;
            signal word_access_2_1310_symbol : Boolean;
            signal word_access_3_1315_symbol : Boolean;
            -- 
          begin -- 
            word_access_1297_start <= Xentry_1295_symbol; -- control passed to block
            Xentry_1298_symbol  <= word_access_1297_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/$entry
            word_access_0_1300: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0 
              signal word_access_0_1300_start: Boolean;
              signal Xentry_1301_symbol: Boolean;
              signal Xexit_1302_symbol: Boolean;
              signal cr_1303_symbol : Boolean;
              signal ca_1304_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1300_start <= Xentry_1298_symbol; -- control passed to block
              Xentry_1301_symbol  <= word_access_0_1300_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/$entry
              cr_1303_symbol <= Xentry_1301_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/cr
              ptr_deref_223_store_0_req_1 <= cr_1303_symbol; -- link to DP
              ca_1304_symbol <= ptr_deref_223_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/ca
              Xexit_1302_symbol <= ca_1304_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/$exit
              word_access_0_1300_symbol <= Xexit_1302_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0
            word_access_1_1305: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_1 
              signal word_access_1_1305_start: Boolean;
              signal Xentry_1306_symbol: Boolean;
              signal Xexit_1307_symbol: Boolean;
              signal cr_1308_symbol : Boolean;
              signal ca_1309_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1305_start <= Xentry_1298_symbol; -- control passed to block
              Xentry_1306_symbol  <= word_access_1_1305_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_1/$entry
              cr_1308_symbol <= Xentry_1306_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_1/cr
              ptr_deref_223_store_1_req_1 <= cr_1308_symbol; -- link to DP
              ca_1309_symbol <= ptr_deref_223_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_1/ca
              Xexit_1307_symbol <= ca_1309_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_1/$exit
              word_access_1_1305_symbol <= Xexit_1307_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_1
            word_access_2_1310: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_2 
              signal word_access_2_1310_start: Boolean;
              signal Xentry_1311_symbol: Boolean;
              signal Xexit_1312_symbol: Boolean;
              signal cr_1313_symbol : Boolean;
              signal ca_1314_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1310_start <= Xentry_1298_symbol; -- control passed to block
              Xentry_1311_symbol  <= word_access_2_1310_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_2/$entry
              cr_1313_symbol <= Xentry_1311_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_2/cr
              ptr_deref_223_store_2_req_1 <= cr_1313_symbol; -- link to DP
              ca_1314_symbol <= ptr_deref_223_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_2/ca
              Xexit_1312_symbol <= ca_1314_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_2/$exit
              word_access_2_1310_symbol <= Xexit_1312_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_2
            word_access_3_1315: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_3 
              signal word_access_3_1315_start: Boolean;
              signal Xentry_1316_symbol: Boolean;
              signal Xexit_1317_symbol: Boolean;
              signal cr_1318_symbol : Boolean;
              signal ca_1319_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1315_start <= Xentry_1298_symbol; -- control passed to block
              Xentry_1316_symbol  <= word_access_3_1315_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_3/$entry
              cr_1318_symbol <= Xentry_1316_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_3/cr
              ptr_deref_223_store_3_req_1 <= cr_1318_symbol; -- link to DP
              ca_1319_symbol <= ptr_deref_223_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_3/ca
              Xexit_1317_symbol <= ca_1319_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_3/$exit
              word_access_3_1315_symbol <= Xexit_1317_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_3
            Xexit_1299_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/$exit 
              signal Xexit_1299_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1299_predecessors(0) <= word_access_0_1300_symbol;
              Xexit_1299_predecessors(1) <= word_access_1_1305_symbol;
              Xexit_1299_predecessors(2) <= word_access_2_1310_symbol;
              Xexit_1299_predecessors(3) <= word_access_3_1315_symbol;
              Xexit_1299_join: join -- 
                port map( -- 
                  preds => Xexit_1299_predecessors,
                  symbol_out => Xexit_1299_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/$exit
            word_access_1297_symbol <= Xexit_1299_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access
          Xexit_1296_symbol <= word_access_1297_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/$exit
          ptr_deref_223_complete_1294_symbol <= Xexit_1296_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete
        Xexit_849_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/$exit 
          signal Xexit_849_predecessors: BooleanArray(5 downto 0);
          -- 
        begin -- 
          Xexit_849_predecessors(0) <= ptr_deref_183_base_address_calculated_854_symbol;
          Xexit_849_predecessors(1) <= ptr_deref_197_base_address_calculated_964_symbol;
          Xexit_849_predecessors(2) <= assign_stmt_212_completed_x_x1081_symbol;
          Xexit_849_predecessors(3) <= ptr_deref_215_base_address_calculated_1189_symbol;
          Xexit_849_predecessors(4) <= assign_stmt_225_completed_x_x1259_symbol;
          Xexit_849_predecessors(5) <= ptr_deref_223_base_address_calculated_1263_symbol;
          Xexit_849_join: join -- 
            port map( -- 
              preds => Xexit_849_predecessors,
              symbol_out => Xexit_849_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/$exit
        assign_stmt_184_to_assign_stmt_225_847_symbol <= Xexit_849_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225
      assign_stmt_233_to_assign_stmt_245_1320: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245 
        signal assign_stmt_233_to_assign_stmt_245_1320_start: Boolean;
        signal Xentry_1321_symbol: Boolean;
        signal Xexit_1322_symbol: Boolean;
        signal assign_stmt_237_active_x_x1323_symbol : Boolean;
        signal assign_stmt_237_completed_x_x1324_symbol : Boolean;
        signal ptr_deref_235_trigger_x_x1325_symbol : Boolean;
        signal ptr_deref_235_active_x_x1326_symbol : Boolean;
        signal ptr_deref_235_base_address_calculated_1327_symbol : Boolean;
        signal ptr_deref_235_root_address_calculated_1328_symbol : Boolean;
        signal ptr_deref_235_word_address_calculated_1329_symbol : Boolean;
        signal ptr_deref_235_request_1330_symbol : Boolean;
        signal ptr_deref_235_complete_1358_symbol : Boolean;
        signal assign_stmt_245_active_x_x1384_symbol : Boolean;
        signal assign_stmt_245_completed_x_x1385_symbol : Boolean;
        signal simple_obj_ref_243_trigger_x_x1386_symbol : Boolean;
        signal simple_obj_ref_243_active_x_x1387_symbol : Boolean;
        signal simple_obj_ref_243_root_address_calculated_1388_symbol : Boolean;
        signal simple_obj_ref_243_word_address_calculated_1389_symbol : Boolean;
        signal simple_obj_ref_243_request_1390_symbol : Boolean;
        signal simple_obj_ref_243_complete_1403_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_233_to_assign_stmt_245_1320_start <= assign_stmt_233_to_assign_stmt_245_x_xentry_x_xx_x636_symbol; -- control passed to block
        Xentry_1321_symbol  <= assign_stmt_233_to_assign_stmt_245_1320_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/$entry
        assign_stmt_237_active_x_x1323_symbol <= Xentry_1321_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_237_active_
        assign_stmt_237_completed_x_x1324_symbol <= ptr_deref_235_complete_1358_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_237_completed_
        ptr_deref_235_trigger_x_x1325_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_trigger_ 
          signal ptr_deref_235_trigger_x_x1325_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_235_trigger_x_x1325_predecessors(0) <= ptr_deref_235_word_address_calculated_1329_symbol;
          ptr_deref_235_trigger_x_x1325_predecessors(1) <= assign_stmt_237_active_x_x1323_symbol;
          ptr_deref_235_trigger_x_x1325_join: join -- 
            port map( -- 
              preds => ptr_deref_235_trigger_x_x1325_predecessors,
              symbol_out => ptr_deref_235_trigger_x_x1325_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_trigger_
        ptr_deref_235_active_x_x1326_symbol <= ptr_deref_235_request_1330_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_active_
        ptr_deref_235_base_address_calculated_1327_symbol <= Xentry_1321_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_base_address_calculated
        ptr_deref_235_root_address_calculated_1328_symbol <= Xentry_1321_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_root_address_calculated
        ptr_deref_235_word_address_calculated_1329_symbol <= ptr_deref_235_root_address_calculated_1328_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_word_address_calculated
        ptr_deref_235_request_1330: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request 
          signal ptr_deref_235_request_1330_start: Boolean;
          signal Xentry_1331_symbol: Boolean;
          signal Xexit_1332_symbol: Boolean;
          signal split_req_1333_symbol : Boolean;
          signal split_ack_1334_symbol : Boolean;
          signal word_access_1335_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_235_request_1330_start <= ptr_deref_235_trigger_x_x1325_symbol; -- control passed to block
          Xentry_1331_symbol  <= ptr_deref_235_request_1330_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/$entry
          split_req_1333_symbol <= Xentry_1331_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/split_req
          ptr_deref_235_gather_scatter_req_0 <= split_req_1333_symbol; -- link to DP
          split_ack_1334_symbol <= ptr_deref_235_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/split_ack
          word_access_1335: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access 
            signal word_access_1335_start: Boolean;
            signal Xentry_1336_symbol: Boolean;
            signal Xexit_1337_symbol: Boolean;
            signal word_access_0_1338_symbol : Boolean;
            signal word_access_1_1343_symbol : Boolean;
            signal word_access_2_1348_symbol : Boolean;
            signal word_access_3_1353_symbol : Boolean;
            -- 
          begin -- 
            word_access_1335_start <= split_ack_1334_symbol; -- control passed to block
            Xentry_1336_symbol  <= word_access_1335_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/$entry
            word_access_0_1338: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0 
              signal word_access_0_1338_start: Boolean;
              signal Xentry_1339_symbol: Boolean;
              signal Xexit_1340_symbol: Boolean;
              signal rr_1341_symbol : Boolean;
              signal ra_1342_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1338_start <= Xentry_1336_symbol; -- control passed to block
              Xentry_1339_symbol  <= word_access_0_1338_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/$entry
              rr_1341_symbol <= Xentry_1339_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/rr
              ptr_deref_235_store_0_req_0 <= rr_1341_symbol; -- link to DP
              ra_1342_symbol <= ptr_deref_235_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/ra
              Xexit_1340_symbol <= ra_1342_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/$exit
              word_access_0_1338_symbol <= Xexit_1340_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0
            word_access_1_1343: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_1 
              signal word_access_1_1343_start: Boolean;
              signal Xentry_1344_symbol: Boolean;
              signal Xexit_1345_symbol: Boolean;
              signal rr_1346_symbol : Boolean;
              signal ra_1347_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1343_start <= Xentry_1336_symbol; -- control passed to block
              Xentry_1344_symbol  <= word_access_1_1343_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_1/$entry
              rr_1346_symbol <= Xentry_1344_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_1/rr
              ptr_deref_235_store_1_req_0 <= rr_1346_symbol; -- link to DP
              ra_1347_symbol <= ptr_deref_235_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_1/ra
              Xexit_1345_symbol <= ra_1347_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_1/$exit
              word_access_1_1343_symbol <= Xexit_1345_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_1
            word_access_2_1348: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_2 
              signal word_access_2_1348_start: Boolean;
              signal Xentry_1349_symbol: Boolean;
              signal Xexit_1350_symbol: Boolean;
              signal rr_1351_symbol : Boolean;
              signal ra_1352_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1348_start <= Xentry_1336_symbol; -- control passed to block
              Xentry_1349_symbol  <= word_access_2_1348_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_2/$entry
              rr_1351_symbol <= Xentry_1349_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_2/rr
              ptr_deref_235_store_2_req_0 <= rr_1351_symbol; -- link to DP
              ra_1352_symbol <= ptr_deref_235_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_2/ra
              Xexit_1350_symbol <= ra_1352_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_2/$exit
              word_access_2_1348_symbol <= Xexit_1350_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_2
            word_access_3_1353: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_3 
              signal word_access_3_1353_start: Boolean;
              signal Xentry_1354_symbol: Boolean;
              signal Xexit_1355_symbol: Boolean;
              signal rr_1356_symbol : Boolean;
              signal ra_1357_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1353_start <= Xentry_1336_symbol; -- control passed to block
              Xentry_1354_symbol  <= word_access_3_1353_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_3/$entry
              rr_1356_symbol <= Xentry_1354_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_3/rr
              ptr_deref_235_store_3_req_0 <= rr_1356_symbol; -- link to DP
              ra_1357_symbol <= ptr_deref_235_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_3/ra
              Xexit_1355_symbol <= ra_1357_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_3/$exit
              word_access_3_1353_symbol <= Xexit_1355_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_3
            Xexit_1337_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/$exit 
              signal Xexit_1337_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1337_predecessors(0) <= word_access_0_1338_symbol;
              Xexit_1337_predecessors(1) <= word_access_1_1343_symbol;
              Xexit_1337_predecessors(2) <= word_access_2_1348_symbol;
              Xexit_1337_predecessors(3) <= word_access_3_1353_symbol;
              Xexit_1337_join: join -- 
                port map( -- 
                  preds => Xexit_1337_predecessors,
                  symbol_out => Xexit_1337_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/$exit
            word_access_1335_symbol <= Xexit_1337_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access
          Xexit_1332_symbol <= word_access_1335_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/$exit
          ptr_deref_235_request_1330_symbol <= Xexit_1332_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request
        ptr_deref_235_complete_1358: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete 
          signal ptr_deref_235_complete_1358_start: Boolean;
          signal Xentry_1359_symbol: Boolean;
          signal Xexit_1360_symbol: Boolean;
          signal word_access_1361_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_235_complete_1358_start <= ptr_deref_235_active_x_x1326_symbol; -- control passed to block
          Xentry_1359_symbol  <= ptr_deref_235_complete_1358_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/$entry
          word_access_1361: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access 
            signal word_access_1361_start: Boolean;
            signal Xentry_1362_symbol: Boolean;
            signal Xexit_1363_symbol: Boolean;
            signal word_access_0_1364_symbol : Boolean;
            signal word_access_1_1369_symbol : Boolean;
            signal word_access_2_1374_symbol : Boolean;
            signal word_access_3_1379_symbol : Boolean;
            -- 
          begin -- 
            word_access_1361_start <= Xentry_1359_symbol; -- control passed to block
            Xentry_1362_symbol  <= word_access_1361_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/$entry
            word_access_0_1364: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0 
              signal word_access_0_1364_start: Boolean;
              signal Xentry_1365_symbol: Boolean;
              signal Xexit_1366_symbol: Boolean;
              signal cr_1367_symbol : Boolean;
              signal ca_1368_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1364_start <= Xentry_1362_symbol; -- control passed to block
              Xentry_1365_symbol  <= word_access_0_1364_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/$entry
              cr_1367_symbol <= Xentry_1365_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/cr
              ptr_deref_235_store_0_req_1 <= cr_1367_symbol; -- link to DP
              ca_1368_symbol <= ptr_deref_235_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/ca
              Xexit_1366_symbol <= ca_1368_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/$exit
              word_access_0_1364_symbol <= Xexit_1366_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0
            word_access_1_1369: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_1 
              signal word_access_1_1369_start: Boolean;
              signal Xentry_1370_symbol: Boolean;
              signal Xexit_1371_symbol: Boolean;
              signal cr_1372_symbol : Boolean;
              signal ca_1373_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1369_start <= Xentry_1362_symbol; -- control passed to block
              Xentry_1370_symbol  <= word_access_1_1369_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_1/$entry
              cr_1372_symbol <= Xentry_1370_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_1/cr
              ptr_deref_235_store_1_req_1 <= cr_1372_symbol; -- link to DP
              ca_1373_symbol <= ptr_deref_235_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_1/ca
              Xexit_1371_symbol <= ca_1373_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_1/$exit
              word_access_1_1369_symbol <= Xexit_1371_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_1
            word_access_2_1374: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_2 
              signal word_access_2_1374_start: Boolean;
              signal Xentry_1375_symbol: Boolean;
              signal Xexit_1376_symbol: Boolean;
              signal cr_1377_symbol : Boolean;
              signal ca_1378_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1374_start <= Xentry_1362_symbol; -- control passed to block
              Xentry_1375_symbol  <= word_access_2_1374_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_2/$entry
              cr_1377_symbol <= Xentry_1375_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_2/cr
              ptr_deref_235_store_2_req_1 <= cr_1377_symbol; -- link to DP
              ca_1378_symbol <= ptr_deref_235_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_2/ca
              Xexit_1376_symbol <= ca_1378_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_2/$exit
              word_access_2_1374_symbol <= Xexit_1376_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_2
            word_access_3_1379: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_3 
              signal word_access_3_1379_start: Boolean;
              signal Xentry_1380_symbol: Boolean;
              signal Xexit_1381_symbol: Boolean;
              signal cr_1382_symbol : Boolean;
              signal ca_1383_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1379_start <= Xentry_1362_symbol; -- control passed to block
              Xentry_1380_symbol  <= word_access_3_1379_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_3/$entry
              cr_1382_symbol <= Xentry_1380_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_3/cr
              ptr_deref_235_store_3_req_1 <= cr_1382_symbol; -- link to DP
              ca_1383_symbol <= ptr_deref_235_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_3/ca
              Xexit_1381_symbol <= ca_1383_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_3/$exit
              word_access_3_1379_symbol <= Xexit_1381_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_3
            Xexit_1363_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/$exit 
              signal Xexit_1363_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1363_predecessors(0) <= word_access_0_1364_symbol;
              Xexit_1363_predecessors(1) <= word_access_1_1369_symbol;
              Xexit_1363_predecessors(2) <= word_access_2_1374_symbol;
              Xexit_1363_predecessors(3) <= word_access_3_1379_symbol;
              Xexit_1363_join: join -- 
                port map( -- 
                  preds => Xexit_1363_predecessors,
                  symbol_out => Xexit_1363_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/$exit
            word_access_1361_symbol <= Xexit_1363_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access
          Xexit_1360_symbol <= word_access_1361_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/$exit
          ptr_deref_235_complete_1358_symbol <= Xexit_1360_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete
        assign_stmt_245_active_x_x1384_symbol <= Xentry_1321_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_245_active_
        assign_stmt_245_completed_x_x1385_symbol <= simple_obj_ref_243_complete_1403_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_245_completed_
        simple_obj_ref_243_trigger_x_x1386_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_trigger_ 
          signal simple_obj_ref_243_trigger_x_x1386_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          simple_obj_ref_243_trigger_x_x1386_predecessors(0) <= simple_obj_ref_243_word_address_calculated_1389_symbol;
          simple_obj_ref_243_trigger_x_x1386_predecessors(1) <= assign_stmt_245_active_x_x1384_symbol;
          simple_obj_ref_243_trigger_x_x1386_join: join -- 
            port map( -- 
              preds => simple_obj_ref_243_trigger_x_x1386_predecessors,
              symbol_out => simple_obj_ref_243_trigger_x_x1386_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_trigger_
        simple_obj_ref_243_active_x_x1387_symbol <= simple_obj_ref_243_request_1390_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_active_
        simple_obj_ref_243_root_address_calculated_1388_symbol <= Xentry_1321_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_root_address_calculated
        simple_obj_ref_243_word_address_calculated_1389_symbol <= simple_obj_ref_243_root_address_calculated_1388_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_word_address_calculated
        simple_obj_ref_243_request_1390: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request 
          signal simple_obj_ref_243_request_1390_start: Boolean;
          signal Xentry_1391_symbol: Boolean;
          signal Xexit_1392_symbol: Boolean;
          signal split_req_1393_symbol : Boolean;
          signal split_ack_1394_symbol : Boolean;
          signal word_access_1395_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_243_request_1390_start <= simple_obj_ref_243_trigger_x_x1386_symbol; -- control passed to block
          Xentry_1391_symbol  <= simple_obj_ref_243_request_1390_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/$entry
          split_req_1393_symbol <= Xentry_1391_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/split_req
          simple_obj_ref_243_gather_scatter_req_0 <= split_req_1393_symbol; -- link to DP
          split_ack_1394_symbol <= simple_obj_ref_243_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/split_ack
          word_access_1395: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access 
            signal word_access_1395_start: Boolean;
            signal Xentry_1396_symbol: Boolean;
            signal Xexit_1397_symbol: Boolean;
            signal word_access_0_1398_symbol : Boolean;
            -- 
          begin -- 
            word_access_1395_start <= split_ack_1394_symbol; -- control passed to block
            Xentry_1396_symbol  <= word_access_1395_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/$entry
            word_access_0_1398: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0 
              signal word_access_0_1398_start: Boolean;
              signal Xentry_1399_symbol: Boolean;
              signal Xexit_1400_symbol: Boolean;
              signal rr_1401_symbol : Boolean;
              signal ra_1402_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1398_start <= Xentry_1396_symbol; -- control passed to block
              Xentry_1399_symbol  <= word_access_0_1398_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/$entry
              rr_1401_symbol <= Xentry_1399_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/rr
              simple_obj_ref_243_store_0_req_0 <= rr_1401_symbol; -- link to DP
              ra_1402_symbol <= simple_obj_ref_243_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/ra
              Xexit_1400_symbol <= ra_1402_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/$exit
              word_access_0_1398_symbol <= Xexit_1400_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0
            Xexit_1397_symbol <= word_access_0_1398_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/$exit
            word_access_1395_symbol <= Xexit_1397_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access
          Xexit_1392_symbol <= word_access_1395_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/$exit
          simple_obj_ref_243_request_1390_symbol <= Xexit_1392_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request
        simple_obj_ref_243_complete_1403: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete 
          signal simple_obj_ref_243_complete_1403_start: Boolean;
          signal Xentry_1404_symbol: Boolean;
          signal Xexit_1405_symbol: Boolean;
          signal word_access_1406_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_243_complete_1403_start <= simple_obj_ref_243_active_x_x1387_symbol; -- control passed to block
          Xentry_1404_symbol  <= simple_obj_ref_243_complete_1403_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/$entry
          word_access_1406: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access 
            signal word_access_1406_start: Boolean;
            signal Xentry_1407_symbol: Boolean;
            signal Xexit_1408_symbol: Boolean;
            signal word_access_0_1409_symbol : Boolean;
            -- 
          begin -- 
            word_access_1406_start <= Xentry_1404_symbol; -- control passed to block
            Xentry_1407_symbol  <= word_access_1406_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/$entry
            word_access_0_1409: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0 
              signal word_access_0_1409_start: Boolean;
              signal Xentry_1410_symbol: Boolean;
              signal Xexit_1411_symbol: Boolean;
              signal cr_1412_symbol : Boolean;
              signal ca_1413_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1409_start <= Xentry_1407_symbol; -- control passed to block
              Xentry_1410_symbol  <= word_access_0_1409_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/$entry
              cr_1412_symbol <= Xentry_1410_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/cr
              simple_obj_ref_243_store_0_req_1 <= cr_1412_symbol; -- link to DP
              ca_1413_symbol <= simple_obj_ref_243_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/ca
              Xexit_1411_symbol <= ca_1413_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/$exit
              word_access_0_1409_symbol <= Xexit_1411_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0
            Xexit_1408_symbol <= word_access_0_1409_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/$exit
            word_access_1406_symbol <= Xexit_1408_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access
          Xexit_1405_symbol <= word_access_1406_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/$exit
          simple_obj_ref_243_complete_1403_symbol <= Xexit_1405_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete
        Xexit_1322_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/$exit 
          signal Xexit_1322_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          Xexit_1322_predecessors(0) <= assign_stmt_237_completed_x_x1324_symbol;
          Xexit_1322_predecessors(1) <= ptr_deref_235_base_address_calculated_1327_symbol;
          Xexit_1322_predecessors(2) <= assign_stmt_245_completed_x_x1385_symbol;
          Xexit_1322_join: join -- 
            port map( -- 
              preds => Xexit_1322_predecessors,
              symbol_out => Xexit_1322_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/$exit
        assign_stmt_233_to_assign_stmt_245_1320_symbol <= Xexit_1322_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245
      assign_stmt_252_1414: Block -- branch_block_stmt_134/assign_stmt_252 
        signal assign_stmt_252_1414_start: Boolean;
        signal Xentry_1415_symbol: Boolean;
        signal Xexit_1416_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_252_1414_start <= assign_stmt_252_x_xentry_x_xx_x640_symbol; -- control passed to block
        Xentry_1415_symbol  <= assign_stmt_252_1414_start; -- transition branch_block_stmt_134/assign_stmt_252/$entry
        Xexit_1416_symbol <= Xentry_1415_symbol; -- transition branch_block_stmt_134/assign_stmt_252/$exit
        assign_stmt_252_1414_symbol <= Xexit_1416_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_252
      assign_stmt_256_1417: Block -- branch_block_stmt_134/assign_stmt_256 
        signal assign_stmt_256_1417_start: Boolean;
        signal Xentry_1418_symbol: Boolean;
        signal Xexit_1419_symbol: Boolean;
        signal assign_stmt_256_active_x_x1420_symbol : Boolean;
        signal assign_stmt_256_completed_x_x1421_symbol : Boolean;
        signal type_cast_255_active_x_x1422_symbol : Boolean;
        signal type_cast_255_trigger_x_x1423_symbol : Boolean;
        signal simple_obj_ref_254_trigger_x_x1424_symbol : Boolean;
        signal simple_obj_ref_254_complete_1425_symbol : Boolean;
        signal type_cast_255_complete_1430_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_256_1417_start <= assign_stmt_256_x_xentry_x_xx_x642_symbol; -- control passed to block
        Xentry_1418_symbol  <= assign_stmt_256_1417_start; -- transition branch_block_stmt_134/assign_stmt_256/$entry
        assign_stmt_256_active_x_x1420_symbol <= type_cast_255_complete_1430_symbol; -- transition branch_block_stmt_134/assign_stmt_256/assign_stmt_256_active_
        assign_stmt_256_completed_x_x1421_symbol <= assign_stmt_256_active_x_x1420_symbol; -- transition branch_block_stmt_134/assign_stmt_256/assign_stmt_256_completed_
        type_cast_255_active_x_x1422_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_256/type_cast_255_active_ 
          signal type_cast_255_active_x_x1422_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_255_active_x_x1422_predecessors(0) <= type_cast_255_trigger_x_x1423_symbol;
          type_cast_255_active_x_x1422_predecessors(1) <= simple_obj_ref_254_complete_1425_symbol;
          type_cast_255_active_x_x1422_join: join -- 
            port map( -- 
              preds => type_cast_255_active_x_x1422_predecessors,
              symbol_out => type_cast_255_active_x_x1422_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_256/type_cast_255_active_
        type_cast_255_trigger_x_x1423_symbol <= Xentry_1418_symbol; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_trigger_
        simple_obj_ref_254_trigger_x_x1424_symbol <= Xentry_1418_symbol; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_trigger_
        simple_obj_ref_254_complete_1425: Block -- branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete 
          signal simple_obj_ref_254_complete_1425_start: Boolean;
          signal Xentry_1426_symbol: Boolean;
          signal Xexit_1427_symbol: Boolean;
          signal req_1428_symbol : Boolean;
          signal ack_1429_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_254_complete_1425_start <= simple_obj_ref_254_trigger_x_x1424_symbol; -- control passed to block
          Xentry_1426_symbol  <= simple_obj_ref_254_complete_1425_start; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/$entry
          req_1428_symbol <= Xentry_1426_symbol; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/req
          simple_obj_ref_254_inst_req_0 <= req_1428_symbol; -- link to DP
          ack_1429_symbol <= simple_obj_ref_254_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/ack
          Xexit_1427_symbol <= ack_1429_symbol; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/$exit
          simple_obj_ref_254_complete_1425_symbol <= Xexit_1427_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete
        type_cast_255_complete_1430: Block -- branch_block_stmt_134/assign_stmt_256/type_cast_255_complete 
          signal type_cast_255_complete_1430_start: Boolean;
          signal Xentry_1431_symbol: Boolean;
          signal Xexit_1432_symbol: Boolean;
          signal req_1433_symbol : Boolean;
          signal ack_1434_symbol : Boolean;
          -- 
        begin -- 
          type_cast_255_complete_1430_start <= type_cast_255_active_x_x1422_symbol; -- control passed to block
          Xentry_1431_symbol  <= type_cast_255_complete_1430_start; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/$entry
          req_1433_symbol <= Xentry_1431_symbol; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/req
          type_cast_255_inst_req_0 <= req_1433_symbol; -- link to DP
          ack_1434_symbol <= type_cast_255_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/ack
          Xexit_1432_symbol <= ack_1434_symbol; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/$exit
          type_cast_255_complete_1430_symbol <= Xexit_1432_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_256/type_cast_255_complete
        Xexit_1419_symbol <= assign_stmt_256_completed_x_x1421_symbol; -- transition branch_block_stmt_134/assign_stmt_256/$exit
        assign_stmt_256_1417_symbol <= Xexit_1419_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_256
      assign_stmt_260_to_assign_stmt_273_1435: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273 
        signal assign_stmt_260_to_assign_stmt_273_1435_start: Boolean;
        signal Xentry_1436_symbol: Boolean;
        signal Xexit_1437_symbol: Boolean;
        signal assign_stmt_260_active_x_x1438_symbol : Boolean;
        signal assign_stmt_260_completed_x_x1439_symbol : Boolean;
        signal simple_obj_ref_259_complete_1440_symbol : Boolean;
        signal ptr_deref_258_trigger_x_x1441_symbol : Boolean;
        signal ptr_deref_258_active_x_x1442_symbol : Boolean;
        signal ptr_deref_258_base_address_calculated_1443_symbol : Boolean;
        signal ptr_deref_258_root_address_calculated_1444_symbol : Boolean;
        signal ptr_deref_258_word_address_calculated_1445_symbol : Boolean;
        signal ptr_deref_258_request_1446_symbol : Boolean;
        signal ptr_deref_258_complete_1459_symbol : Boolean;
        signal assign_stmt_264_active_x_x1470_symbol : Boolean;
        signal assign_stmt_264_completed_x_x1471_symbol : Boolean;
        signal ptr_deref_263_trigger_x_x1472_symbol : Boolean;
        signal ptr_deref_263_active_x_x1473_symbol : Boolean;
        signal ptr_deref_263_base_address_calculated_1474_symbol : Boolean;
        signal ptr_deref_263_root_address_calculated_1475_symbol : Boolean;
        signal ptr_deref_263_word_address_calculated_1476_symbol : Boolean;
        signal ptr_deref_263_request_1477_symbol : Boolean;
        signal ptr_deref_263_complete_1488_symbol : Boolean;
        signal assign_stmt_268_active_x_x1501_symbol : Boolean;
        signal assign_stmt_268_completed_x_x1502_symbol : Boolean;
        signal type_cast_267_active_x_x1503_symbol : Boolean;
        signal type_cast_267_trigger_x_x1504_symbol : Boolean;
        signal simple_obj_ref_266_complete_1505_symbol : Boolean;
        signal type_cast_267_complete_1506_symbol : Boolean;
        signal assign_stmt_273_active_x_x1511_symbol : Boolean;
        signal assign_stmt_273_completed_x_x1512_symbol : Boolean;
        signal binary_272_active_x_x1513_symbol : Boolean;
        signal binary_272_trigger_x_x1514_symbol : Boolean;
        signal simple_obj_ref_270_complete_1515_symbol : Boolean;
        signal binary_272_complete_1516_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_260_to_assign_stmt_273_1435_start <= assign_stmt_260_to_assign_stmt_273_x_xentry_x_xx_x644_symbol; -- control passed to block
        Xentry_1436_symbol  <= assign_stmt_260_to_assign_stmt_273_1435_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/$entry
        assign_stmt_260_active_x_x1438_symbol <= simple_obj_ref_259_complete_1440_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_260_active_
        assign_stmt_260_completed_x_x1439_symbol <= ptr_deref_258_complete_1459_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_260_completed_
        simple_obj_ref_259_complete_1440_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/simple_obj_ref_259_complete
        ptr_deref_258_trigger_x_x1441_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_trigger_ 
          signal ptr_deref_258_trigger_x_x1441_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_258_trigger_x_x1441_predecessors(0) <= ptr_deref_258_word_address_calculated_1445_symbol;
          ptr_deref_258_trigger_x_x1441_predecessors(1) <= assign_stmt_260_active_x_x1438_symbol;
          ptr_deref_258_trigger_x_x1441_join: join -- 
            port map( -- 
              preds => ptr_deref_258_trigger_x_x1441_predecessors,
              symbol_out => ptr_deref_258_trigger_x_x1441_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_trigger_
        ptr_deref_258_active_x_x1442_symbol <= ptr_deref_258_request_1446_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_active_
        ptr_deref_258_base_address_calculated_1443_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_base_address_calculated
        ptr_deref_258_root_address_calculated_1444_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_root_address_calculated
        ptr_deref_258_word_address_calculated_1445_symbol <= ptr_deref_258_root_address_calculated_1444_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_word_address_calculated
        ptr_deref_258_request_1446: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request 
          signal ptr_deref_258_request_1446_start: Boolean;
          signal Xentry_1447_symbol: Boolean;
          signal Xexit_1448_symbol: Boolean;
          signal split_req_1449_symbol : Boolean;
          signal split_ack_1450_symbol : Boolean;
          signal word_access_1451_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_258_request_1446_start <= ptr_deref_258_trigger_x_x1441_symbol; -- control passed to block
          Xentry_1447_symbol  <= ptr_deref_258_request_1446_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/$entry
          split_req_1449_symbol <= Xentry_1447_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/split_req
          ptr_deref_258_gather_scatter_req_0 <= split_req_1449_symbol; -- link to DP
          split_ack_1450_symbol <= ptr_deref_258_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/split_ack
          word_access_1451: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access 
            signal word_access_1451_start: Boolean;
            signal Xentry_1452_symbol: Boolean;
            signal Xexit_1453_symbol: Boolean;
            signal word_access_0_1454_symbol : Boolean;
            -- 
          begin -- 
            word_access_1451_start <= split_ack_1450_symbol; -- control passed to block
            Xentry_1452_symbol  <= word_access_1451_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/$entry
            word_access_0_1454: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0 
              signal word_access_0_1454_start: Boolean;
              signal Xentry_1455_symbol: Boolean;
              signal Xexit_1456_symbol: Boolean;
              signal rr_1457_symbol : Boolean;
              signal ra_1458_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1454_start <= Xentry_1452_symbol; -- control passed to block
              Xentry_1455_symbol  <= word_access_0_1454_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/$entry
              rr_1457_symbol <= Xentry_1455_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/rr
              ptr_deref_258_store_0_req_0 <= rr_1457_symbol; -- link to DP
              ra_1458_symbol <= ptr_deref_258_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/ra
              Xexit_1456_symbol <= ra_1458_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/$exit
              word_access_0_1454_symbol <= Xexit_1456_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0
            Xexit_1453_symbol <= word_access_0_1454_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/$exit
            word_access_1451_symbol <= Xexit_1453_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access
          Xexit_1448_symbol <= word_access_1451_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/$exit
          ptr_deref_258_request_1446_symbol <= Xexit_1448_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request
        ptr_deref_258_complete_1459: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete 
          signal ptr_deref_258_complete_1459_start: Boolean;
          signal Xentry_1460_symbol: Boolean;
          signal Xexit_1461_symbol: Boolean;
          signal word_access_1462_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_258_complete_1459_start <= ptr_deref_258_active_x_x1442_symbol; -- control passed to block
          Xentry_1460_symbol  <= ptr_deref_258_complete_1459_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/$entry
          word_access_1462: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access 
            signal word_access_1462_start: Boolean;
            signal Xentry_1463_symbol: Boolean;
            signal Xexit_1464_symbol: Boolean;
            signal word_access_0_1465_symbol : Boolean;
            -- 
          begin -- 
            word_access_1462_start <= Xentry_1460_symbol; -- control passed to block
            Xentry_1463_symbol  <= word_access_1462_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/$entry
            word_access_0_1465: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0 
              signal word_access_0_1465_start: Boolean;
              signal Xentry_1466_symbol: Boolean;
              signal Xexit_1467_symbol: Boolean;
              signal cr_1468_symbol : Boolean;
              signal ca_1469_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1465_start <= Xentry_1463_symbol; -- control passed to block
              Xentry_1466_symbol  <= word_access_0_1465_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/$entry
              cr_1468_symbol <= Xentry_1466_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/cr
              ptr_deref_258_store_0_req_1 <= cr_1468_symbol; -- link to DP
              ca_1469_symbol <= ptr_deref_258_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/ca
              Xexit_1467_symbol <= ca_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/$exit
              word_access_0_1465_symbol <= Xexit_1467_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0
            Xexit_1464_symbol <= word_access_0_1465_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/$exit
            word_access_1462_symbol <= Xexit_1464_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access
          Xexit_1461_symbol <= word_access_1462_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/$exit
          ptr_deref_258_complete_1459_symbol <= Xexit_1461_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete
        assign_stmt_264_active_x_x1470_symbol <= ptr_deref_263_complete_1488_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_264_active_
        assign_stmt_264_completed_x_x1471_symbol <= assign_stmt_264_active_x_x1470_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_264_completed_
        ptr_deref_263_trigger_x_x1472_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_trigger_ 
          signal ptr_deref_263_trigger_x_x1472_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_263_trigger_x_x1472_predecessors(0) <= ptr_deref_263_word_address_calculated_1476_symbol;
          ptr_deref_263_trigger_x_x1472_predecessors(1) <= ptr_deref_258_active_x_x1442_symbol;
          ptr_deref_263_trigger_x_x1472_join: join -- 
            port map( -- 
              preds => ptr_deref_263_trigger_x_x1472_predecessors,
              symbol_out => ptr_deref_263_trigger_x_x1472_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_trigger_
        ptr_deref_263_active_x_x1473_symbol <= ptr_deref_263_request_1477_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_active_
        ptr_deref_263_base_address_calculated_1474_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_base_address_calculated
        ptr_deref_263_root_address_calculated_1475_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_root_address_calculated
        ptr_deref_263_word_address_calculated_1476_symbol <= ptr_deref_263_root_address_calculated_1475_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_word_address_calculated
        ptr_deref_263_request_1477: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request 
          signal ptr_deref_263_request_1477_start: Boolean;
          signal Xentry_1478_symbol: Boolean;
          signal Xexit_1479_symbol: Boolean;
          signal word_access_1480_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_263_request_1477_start <= ptr_deref_263_trigger_x_x1472_symbol; -- control passed to block
          Xentry_1478_symbol  <= ptr_deref_263_request_1477_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/$entry
          word_access_1480: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access 
            signal word_access_1480_start: Boolean;
            signal Xentry_1481_symbol: Boolean;
            signal Xexit_1482_symbol: Boolean;
            signal word_access_0_1483_symbol : Boolean;
            -- 
          begin -- 
            word_access_1480_start <= Xentry_1478_symbol; -- control passed to block
            Xentry_1481_symbol  <= word_access_1480_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/$entry
            word_access_0_1483: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0 
              signal word_access_0_1483_start: Boolean;
              signal Xentry_1484_symbol: Boolean;
              signal Xexit_1485_symbol: Boolean;
              signal rr_1486_symbol : Boolean;
              signal ra_1487_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1483_start <= Xentry_1481_symbol; -- control passed to block
              Xentry_1484_symbol  <= word_access_0_1483_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/$entry
              rr_1486_symbol <= Xentry_1484_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/rr
              ptr_deref_263_load_0_req_0 <= rr_1486_symbol; -- link to DP
              ra_1487_symbol <= ptr_deref_263_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/ra
              Xexit_1485_symbol <= ra_1487_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/$exit
              word_access_0_1483_symbol <= Xexit_1485_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0
            Xexit_1482_symbol <= word_access_0_1483_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/$exit
            word_access_1480_symbol <= Xexit_1482_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access
          Xexit_1479_symbol <= word_access_1480_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/$exit
          ptr_deref_263_request_1477_symbol <= Xexit_1479_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request
        ptr_deref_263_complete_1488: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete 
          signal ptr_deref_263_complete_1488_start: Boolean;
          signal Xentry_1489_symbol: Boolean;
          signal Xexit_1490_symbol: Boolean;
          signal word_access_1491_symbol : Boolean;
          signal merge_req_1499_symbol : Boolean;
          signal merge_ack_1500_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_263_complete_1488_start <= ptr_deref_263_active_x_x1473_symbol; -- control passed to block
          Xentry_1489_symbol  <= ptr_deref_263_complete_1488_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/$entry
          word_access_1491: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access 
            signal word_access_1491_start: Boolean;
            signal Xentry_1492_symbol: Boolean;
            signal Xexit_1493_symbol: Boolean;
            signal word_access_0_1494_symbol : Boolean;
            -- 
          begin -- 
            word_access_1491_start <= Xentry_1489_symbol; -- control passed to block
            Xentry_1492_symbol  <= word_access_1491_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/$entry
            word_access_0_1494: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0 
              signal word_access_0_1494_start: Boolean;
              signal Xentry_1495_symbol: Boolean;
              signal Xexit_1496_symbol: Boolean;
              signal cr_1497_symbol : Boolean;
              signal ca_1498_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1494_start <= Xentry_1492_symbol; -- control passed to block
              Xentry_1495_symbol  <= word_access_0_1494_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/$entry
              cr_1497_symbol <= Xentry_1495_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/cr
              ptr_deref_263_load_0_req_1 <= cr_1497_symbol; -- link to DP
              ca_1498_symbol <= ptr_deref_263_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/ca
              Xexit_1496_symbol <= ca_1498_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/$exit
              word_access_0_1494_symbol <= Xexit_1496_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0
            Xexit_1493_symbol <= word_access_0_1494_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/$exit
            word_access_1491_symbol <= Xexit_1493_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access
          merge_req_1499_symbol <= word_access_1491_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/merge_req
          ptr_deref_263_gather_scatter_req_0 <= merge_req_1499_symbol; -- link to DP
          merge_ack_1500_symbol <= ptr_deref_263_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/merge_ack
          Xexit_1490_symbol <= merge_ack_1500_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/$exit
          ptr_deref_263_complete_1488_symbol <= Xexit_1490_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete
        assign_stmt_268_active_x_x1501_symbol <= type_cast_267_complete_1506_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_268_active_
        assign_stmt_268_completed_x_x1502_symbol <= assign_stmt_268_active_x_x1501_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_268_completed_
        type_cast_267_active_x_x1503_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_active_ 
          signal type_cast_267_active_x_x1503_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_267_active_x_x1503_predecessors(0) <= type_cast_267_trigger_x_x1504_symbol;
          type_cast_267_active_x_x1503_predecessors(1) <= simple_obj_ref_266_complete_1505_symbol;
          type_cast_267_active_x_x1503_join: join -- 
            port map( -- 
              preds => type_cast_267_active_x_x1503_predecessors,
              symbol_out => type_cast_267_active_x_x1503_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_active_
        type_cast_267_trigger_x_x1504_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_trigger_
        simple_obj_ref_266_complete_1505_symbol <= assign_stmt_264_completed_x_x1471_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/simple_obj_ref_266_complete
        type_cast_267_complete_1506: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete 
          signal type_cast_267_complete_1506_start: Boolean;
          signal Xentry_1507_symbol: Boolean;
          signal Xexit_1508_symbol: Boolean;
          signal req_1509_symbol : Boolean;
          signal ack_1510_symbol : Boolean;
          -- 
        begin -- 
          type_cast_267_complete_1506_start <= type_cast_267_active_x_x1503_symbol; -- control passed to block
          Xentry_1507_symbol  <= type_cast_267_complete_1506_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/$entry
          req_1509_symbol <= Xentry_1507_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/req
          type_cast_267_inst_req_0 <= req_1509_symbol; -- link to DP
          ack_1510_symbol <= type_cast_267_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/ack
          Xexit_1508_symbol <= ack_1510_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/$exit
          type_cast_267_complete_1506_symbol <= Xexit_1508_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete
        assign_stmt_273_active_x_x1511_symbol <= binary_272_complete_1516_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_273_active_
        assign_stmt_273_completed_x_x1512_symbol <= assign_stmt_273_active_x_x1511_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_273_completed_
        binary_272_active_x_x1513_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_active_ 
          signal binary_272_active_x_x1513_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_272_active_x_x1513_predecessors(0) <= binary_272_trigger_x_x1514_symbol;
          binary_272_active_x_x1513_predecessors(1) <= simple_obj_ref_270_complete_1515_symbol;
          binary_272_active_x_x1513_join: join -- 
            port map( -- 
              preds => binary_272_active_x_x1513_predecessors,
              symbol_out => binary_272_active_x_x1513_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_active_
        binary_272_trigger_x_x1514_symbol <= Xentry_1436_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_trigger_
        simple_obj_ref_270_complete_1515_symbol <= assign_stmt_268_completed_x_x1502_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/simple_obj_ref_270_complete
        binary_272_complete_1516: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete 
          signal binary_272_complete_1516_start: Boolean;
          signal Xentry_1517_symbol: Boolean;
          signal Xexit_1518_symbol: Boolean;
          signal rr_1519_symbol : Boolean;
          signal ra_1520_symbol : Boolean;
          signal cr_1521_symbol : Boolean;
          signal ca_1522_symbol : Boolean;
          -- 
        begin -- 
          binary_272_complete_1516_start <= binary_272_active_x_x1513_symbol; -- control passed to block
          Xentry_1517_symbol  <= binary_272_complete_1516_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/$entry
          rr_1519_symbol <= Xentry_1517_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/rr
          binary_272_inst_req_0 <= rr_1519_symbol; -- link to DP
          ra_1520_symbol <= binary_272_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/ra
          cr_1521_symbol <= ra_1520_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/cr
          binary_272_inst_req_1 <= cr_1521_symbol; -- link to DP
          ca_1522_symbol <= binary_272_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/ca
          Xexit_1518_symbol <= ca_1522_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/$exit
          binary_272_complete_1516_symbol <= Xexit_1518_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete
        Xexit_1437_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/$exit 
          signal Xexit_1437_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          Xexit_1437_predecessors(0) <= assign_stmt_260_completed_x_x1439_symbol;
          Xexit_1437_predecessors(1) <= ptr_deref_258_base_address_calculated_1443_symbol;
          Xexit_1437_predecessors(2) <= ptr_deref_263_base_address_calculated_1474_symbol;
          Xexit_1437_predecessors(3) <= assign_stmt_273_completed_x_x1512_symbol;
          Xexit_1437_join: join -- 
            port map( -- 
              preds => Xexit_1437_predecessors,
              symbol_out => Xexit_1437_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/$exit
        assign_stmt_260_to_assign_stmt_273_1435_symbol <= Xexit_1437_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273
      if_stmt_274_dead_link_1523: Block -- branch_block_stmt_134/if_stmt_274_dead_link 
        signal if_stmt_274_dead_link_1523_start: Boolean;
        signal Xentry_1524_symbol: Boolean;
        signal Xexit_1525_symbol: Boolean;
        signal dead_transition_1526_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_dead_link_1523_start <= if_stmt_274_x_xentry_x_xx_x646_symbol; -- control passed to block
        Xentry_1524_symbol  <= if_stmt_274_dead_link_1523_start; -- transition branch_block_stmt_134/if_stmt_274_dead_link/$entry
        dead_transition_1526_symbol <= false;
        Xexit_1525_symbol <= dead_transition_1526_symbol; -- transition branch_block_stmt_134/if_stmt_274_dead_link/$exit
        if_stmt_274_dead_link_1523_symbol <= Xexit_1525_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_dead_link
      if_stmt_274_eval_test_1527: Block -- branch_block_stmt_134/if_stmt_274_eval_test 
        signal if_stmt_274_eval_test_1527_start: Boolean;
        signal Xentry_1528_symbol: Boolean;
        signal Xexit_1529_symbol: Boolean;
        signal branch_req_1530_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_eval_test_1527_start <= if_stmt_274_x_xentry_x_xx_x646_symbol; -- control passed to block
        Xentry_1528_symbol  <= if_stmt_274_eval_test_1527_start; -- transition branch_block_stmt_134/if_stmt_274_eval_test/$entry
        branch_req_1530_symbol <= Xentry_1528_symbol; -- transition branch_block_stmt_134/if_stmt_274_eval_test/branch_req
        if_stmt_274_branch_req_0 <= branch_req_1530_symbol; -- link to DP
        Xexit_1529_symbol <= branch_req_1530_symbol; -- transition branch_block_stmt_134/if_stmt_274_eval_test/$exit
        if_stmt_274_eval_test_1527_symbol <= Xexit_1529_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_eval_test
      simple_obj_ref_275_place_1531_symbol  <=  if_stmt_274_eval_test_1527_symbol; -- place branch_block_stmt_134/simple_obj_ref_275_place (optimized away) 
      if_stmt_274_if_link_1532: Block -- branch_block_stmt_134/if_stmt_274_if_link 
        signal if_stmt_274_if_link_1532_start: Boolean;
        signal Xentry_1533_symbol: Boolean;
        signal Xexit_1534_symbol: Boolean;
        signal if_choice_transition_1535_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_if_link_1532_start <= simple_obj_ref_275_place_1531_symbol; -- control passed to block
        Xentry_1533_symbol  <= if_stmt_274_if_link_1532_start; -- transition branch_block_stmt_134/if_stmt_274_if_link/$entry
        if_choice_transition_1535_symbol <= if_stmt_274_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_274_if_link/if_choice_transition
        Xexit_1534_symbol <= if_choice_transition_1535_symbol; -- transition branch_block_stmt_134/if_stmt_274_if_link/$exit
        if_stmt_274_if_link_1532_symbol <= Xexit_1534_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_if_link
      if_stmt_274_else_link_1536: Block -- branch_block_stmt_134/if_stmt_274_else_link 
        signal if_stmt_274_else_link_1536_start: Boolean;
        signal Xentry_1537_symbol: Boolean;
        signal Xexit_1538_symbol: Boolean;
        signal else_choice_transition_1539_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_else_link_1536_start <= simple_obj_ref_275_place_1531_symbol; -- control passed to block
        Xentry_1537_symbol  <= if_stmt_274_else_link_1536_start; -- transition branch_block_stmt_134/if_stmt_274_else_link/$entry
        else_choice_transition_1539_symbol <= if_stmt_274_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_274_else_link/else_choice_transition
        Xexit_1538_symbol <= else_choice_transition_1539_symbol; -- transition branch_block_stmt_134/if_stmt_274_else_link/$exit
        if_stmt_274_else_link_1536_symbol <= Xexit_1538_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_else_link
      bb_4_bb_5_1540_symbol  <=  if_stmt_274_if_link_1532_symbol; -- place branch_block_stmt_134/bb_4_bb_5 (optimized away) 
      bb_4_bb_8_1541_symbol  <=  if_stmt_274_else_link_1536_symbol; -- place branch_block_stmt_134/bb_4_bb_8 (optimized away) 
      assign_stmt_283_to_assign_stmt_297_1542: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297 
        signal assign_stmt_283_to_assign_stmt_297_1542_start: Boolean;
        signal Xentry_1543_symbol: Boolean;
        signal Xexit_1544_symbol: Boolean;
        signal assign_stmt_283_active_x_x1545_symbol : Boolean;
        signal assign_stmt_283_completed_x_x1546_symbol : Boolean;
        signal simple_obj_ref_282_trigger_x_x1547_symbol : Boolean;
        signal simple_obj_ref_282_active_x_x1548_symbol : Boolean;
        signal simple_obj_ref_282_root_address_calculated_1549_symbol : Boolean;
        signal simple_obj_ref_282_word_address_calculated_1550_symbol : Boolean;
        signal simple_obj_ref_282_request_1551_symbol : Boolean;
        signal simple_obj_ref_282_complete_1562_symbol : Boolean;
        signal assign_stmt_287_active_x_x1575_symbol : Boolean;
        signal assign_stmt_287_completed_x_x1576_symbol : Boolean;
        signal simple_obj_ref_286_complete_1577_symbol : Boolean;
        signal ptr_deref_285_trigger_x_x1578_symbol : Boolean;
        signal ptr_deref_285_active_x_x1579_symbol : Boolean;
        signal ptr_deref_285_base_address_calculated_1580_symbol : Boolean;
        signal ptr_deref_285_root_address_calculated_1581_symbol : Boolean;
        signal ptr_deref_285_word_address_calculated_1582_symbol : Boolean;
        signal ptr_deref_285_request_1583_symbol : Boolean;
        signal ptr_deref_285_complete_1611_symbol : Boolean;
        signal assign_stmt_290_active_x_x1637_symbol : Boolean;
        signal assign_stmt_290_completed_x_x1638_symbol : Boolean;
        signal simple_obj_ref_289_trigger_x_x1639_symbol : Boolean;
        signal simple_obj_ref_289_active_x_x1640_symbol : Boolean;
        signal simple_obj_ref_289_root_address_calculated_1641_symbol : Boolean;
        signal simple_obj_ref_289_word_address_calculated_1642_symbol : Boolean;
        signal simple_obj_ref_289_request_1643_symbol : Boolean;
        signal simple_obj_ref_289_complete_1654_symbol : Boolean;
        signal assign_stmt_297_active_x_x1667_symbol : Boolean;
        signal assign_stmt_297_completed_x_x1668_symbol : Boolean;
        signal binary_296_active_x_x1669_symbol : Boolean;
        signal binary_296_trigger_x_x1670_symbol : Boolean;
        signal type_cast_293_active_x_x1671_symbol : Boolean;
        signal type_cast_293_trigger_x_x1672_symbol : Boolean;
        signal simple_obj_ref_292_complete_1673_symbol : Boolean;
        signal type_cast_293_complete_1674_symbol : Boolean;
        signal binary_296_complete_1681_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_283_to_assign_stmt_297_1542_start <= assign_stmt_283_to_assign_stmt_297_x_xentry_x_xx_x650_symbol; -- control passed to block
        Xentry_1543_symbol  <= assign_stmt_283_to_assign_stmt_297_1542_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/$entry
        assign_stmt_283_active_x_x1545_symbol <= simple_obj_ref_282_complete_1562_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_283_active_
        assign_stmt_283_completed_x_x1546_symbol <= assign_stmt_283_active_x_x1545_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_283_completed_
        simple_obj_ref_282_trigger_x_x1547_symbol <= simple_obj_ref_282_word_address_calculated_1550_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_trigger_
        simple_obj_ref_282_active_x_x1548_symbol <= simple_obj_ref_282_request_1551_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_active_
        simple_obj_ref_282_root_address_calculated_1549_symbol <= Xentry_1543_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_root_address_calculated
        simple_obj_ref_282_word_address_calculated_1550_symbol <= simple_obj_ref_282_root_address_calculated_1549_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_word_address_calculated
        simple_obj_ref_282_request_1551: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request 
          signal simple_obj_ref_282_request_1551_start: Boolean;
          signal Xentry_1552_symbol: Boolean;
          signal Xexit_1553_symbol: Boolean;
          signal word_access_1554_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_282_request_1551_start <= simple_obj_ref_282_trigger_x_x1547_symbol; -- control passed to block
          Xentry_1552_symbol  <= simple_obj_ref_282_request_1551_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/$entry
          word_access_1554: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access 
            signal word_access_1554_start: Boolean;
            signal Xentry_1555_symbol: Boolean;
            signal Xexit_1556_symbol: Boolean;
            signal word_access_0_1557_symbol : Boolean;
            -- 
          begin -- 
            word_access_1554_start <= Xentry_1552_symbol; -- control passed to block
            Xentry_1555_symbol  <= word_access_1554_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/$entry
            word_access_0_1557: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0 
              signal word_access_0_1557_start: Boolean;
              signal Xentry_1558_symbol: Boolean;
              signal Xexit_1559_symbol: Boolean;
              signal rr_1560_symbol : Boolean;
              signal ra_1561_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1557_start <= Xentry_1555_symbol; -- control passed to block
              Xentry_1558_symbol  <= word_access_0_1557_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/$entry
              rr_1560_symbol <= Xentry_1558_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/rr
              simple_obj_ref_282_load_0_req_0 <= rr_1560_symbol; -- link to DP
              ra_1561_symbol <= simple_obj_ref_282_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/ra
              Xexit_1559_symbol <= ra_1561_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/$exit
              word_access_0_1557_symbol <= Xexit_1559_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0
            Xexit_1556_symbol <= word_access_0_1557_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/$exit
            word_access_1554_symbol <= Xexit_1556_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access
          Xexit_1553_symbol <= word_access_1554_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/$exit
          simple_obj_ref_282_request_1551_symbol <= Xexit_1553_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request
        simple_obj_ref_282_complete_1562: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete 
          signal simple_obj_ref_282_complete_1562_start: Boolean;
          signal Xentry_1563_symbol: Boolean;
          signal Xexit_1564_symbol: Boolean;
          signal word_access_1565_symbol : Boolean;
          signal merge_req_1573_symbol : Boolean;
          signal merge_ack_1574_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_282_complete_1562_start <= simple_obj_ref_282_active_x_x1548_symbol; -- control passed to block
          Xentry_1563_symbol  <= simple_obj_ref_282_complete_1562_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/$entry
          word_access_1565: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access 
            signal word_access_1565_start: Boolean;
            signal Xentry_1566_symbol: Boolean;
            signal Xexit_1567_symbol: Boolean;
            signal word_access_0_1568_symbol : Boolean;
            -- 
          begin -- 
            word_access_1565_start <= Xentry_1563_symbol; -- control passed to block
            Xentry_1566_symbol  <= word_access_1565_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/$entry
            word_access_0_1568: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0 
              signal word_access_0_1568_start: Boolean;
              signal Xentry_1569_symbol: Boolean;
              signal Xexit_1570_symbol: Boolean;
              signal cr_1571_symbol : Boolean;
              signal ca_1572_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1568_start <= Xentry_1566_symbol; -- control passed to block
              Xentry_1569_symbol  <= word_access_0_1568_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/$entry
              cr_1571_symbol <= Xentry_1569_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/cr
              simple_obj_ref_282_load_0_req_1 <= cr_1571_symbol; -- link to DP
              ca_1572_symbol <= simple_obj_ref_282_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/ca
              Xexit_1570_symbol <= ca_1572_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/$exit
              word_access_0_1568_symbol <= Xexit_1570_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0
            Xexit_1567_symbol <= word_access_0_1568_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/$exit
            word_access_1565_symbol <= Xexit_1567_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access
          merge_req_1573_symbol <= word_access_1565_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/merge_req
          simple_obj_ref_282_gather_scatter_req_0 <= merge_req_1573_symbol; -- link to DP
          merge_ack_1574_symbol <= simple_obj_ref_282_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/merge_ack
          Xexit_1564_symbol <= merge_ack_1574_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/$exit
          simple_obj_ref_282_complete_1562_symbol <= Xexit_1564_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete
        assign_stmt_287_active_x_x1575_symbol <= simple_obj_ref_286_complete_1577_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_287_active_
        assign_stmt_287_completed_x_x1576_symbol <= ptr_deref_285_complete_1611_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_287_completed_
        simple_obj_ref_286_complete_1577_symbol <= assign_stmt_283_completed_x_x1546_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_286_complete
        ptr_deref_285_trigger_x_x1578_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_trigger_ 
          signal ptr_deref_285_trigger_x_x1578_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_285_trigger_x_x1578_predecessors(0) <= ptr_deref_285_word_address_calculated_1582_symbol;
          ptr_deref_285_trigger_x_x1578_predecessors(1) <= assign_stmt_287_active_x_x1575_symbol;
          ptr_deref_285_trigger_x_x1578_join: join -- 
            port map( -- 
              preds => ptr_deref_285_trigger_x_x1578_predecessors,
              symbol_out => ptr_deref_285_trigger_x_x1578_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_trigger_
        ptr_deref_285_active_x_x1579_symbol <= ptr_deref_285_request_1583_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_active_
        ptr_deref_285_base_address_calculated_1580_symbol <= Xentry_1543_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_base_address_calculated
        ptr_deref_285_root_address_calculated_1581_symbol <= Xentry_1543_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_root_address_calculated
        ptr_deref_285_word_address_calculated_1582_symbol <= ptr_deref_285_root_address_calculated_1581_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_word_address_calculated
        ptr_deref_285_request_1583: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request 
          signal ptr_deref_285_request_1583_start: Boolean;
          signal Xentry_1584_symbol: Boolean;
          signal Xexit_1585_symbol: Boolean;
          signal split_req_1586_symbol : Boolean;
          signal split_ack_1587_symbol : Boolean;
          signal word_access_1588_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_285_request_1583_start <= ptr_deref_285_trigger_x_x1578_symbol; -- control passed to block
          Xentry_1584_symbol  <= ptr_deref_285_request_1583_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/$entry
          split_req_1586_symbol <= Xentry_1584_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/split_req
          ptr_deref_285_gather_scatter_req_0 <= split_req_1586_symbol; -- link to DP
          split_ack_1587_symbol <= ptr_deref_285_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/split_ack
          word_access_1588: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access 
            signal word_access_1588_start: Boolean;
            signal Xentry_1589_symbol: Boolean;
            signal Xexit_1590_symbol: Boolean;
            signal word_access_0_1591_symbol : Boolean;
            signal word_access_1_1596_symbol : Boolean;
            signal word_access_2_1601_symbol : Boolean;
            signal word_access_3_1606_symbol : Boolean;
            -- 
          begin -- 
            word_access_1588_start <= split_ack_1587_symbol; -- control passed to block
            Xentry_1589_symbol  <= word_access_1588_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/$entry
            word_access_0_1591: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0 
              signal word_access_0_1591_start: Boolean;
              signal Xentry_1592_symbol: Boolean;
              signal Xexit_1593_symbol: Boolean;
              signal rr_1594_symbol : Boolean;
              signal ra_1595_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1591_start <= Xentry_1589_symbol; -- control passed to block
              Xentry_1592_symbol  <= word_access_0_1591_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/$entry
              rr_1594_symbol <= Xentry_1592_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/rr
              ptr_deref_285_store_0_req_0 <= rr_1594_symbol; -- link to DP
              ra_1595_symbol <= ptr_deref_285_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/ra
              Xexit_1593_symbol <= ra_1595_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/$exit
              word_access_0_1591_symbol <= Xexit_1593_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0
            word_access_1_1596: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_1 
              signal word_access_1_1596_start: Boolean;
              signal Xentry_1597_symbol: Boolean;
              signal Xexit_1598_symbol: Boolean;
              signal rr_1599_symbol : Boolean;
              signal ra_1600_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1596_start <= Xentry_1589_symbol; -- control passed to block
              Xentry_1597_symbol  <= word_access_1_1596_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_1/$entry
              rr_1599_symbol <= Xentry_1597_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_1/rr
              ptr_deref_285_store_1_req_0 <= rr_1599_symbol; -- link to DP
              ra_1600_symbol <= ptr_deref_285_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_1/ra
              Xexit_1598_symbol <= ra_1600_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_1/$exit
              word_access_1_1596_symbol <= Xexit_1598_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_1
            word_access_2_1601: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_2 
              signal word_access_2_1601_start: Boolean;
              signal Xentry_1602_symbol: Boolean;
              signal Xexit_1603_symbol: Boolean;
              signal rr_1604_symbol : Boolean;
              signal ra_1605_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1601_start <= Xentry_1589_symbol; -- control passed to block
              Xentry_1602_symbol  <= word_access_2_1601_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_2/$entry
              rr_1604_symbol <= Xentry_1602_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_2/rr
              ptr_deref_285_store_2_req_0 <= rr_1604_symbol; -- link to DP
              ra_1605_symbol <= ptr_deref_285_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_2/ra
              Xexit_1603_symbol <= ra_1605_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_2/$exit
              word_access_2_1601_symbol <= Xexit_1603_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_2
            word_access_3_1606: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_3 
              signal word_access_3_1606_start: Boolean;
              signal Xentry_1607_symbol: Boolean;
              signal Xexit_1608_symbol: Boolean;
              signal rr_1609_symbol : Boolean;
              signal ra_1610_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1606_start <= Xentry_1589_symbol; -- control passed to block
              Xentry_1607_symbol  <= word_access_3_1606_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_3/$entry
              rr_1609_symbol <= Xentry_1607_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_3/rr
              ptr_deref_285_store_3_req_0 <= rr_1609_symbol; -- link to DP
              ra_1610_symbol <= ptr_deref_285_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_3/ra
              Xexit_1608_symbol <= ra_1610_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_3/$exit
              word_access_3_1606_symbol <= Xexit_1608_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_3
            Xexit_1590_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/$exit 
              signal Xexit_1590_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1590_predecessors(0) <= word_access_0_1591_symbol;
              Xexit_1590_predecessors(1) <= word_access_1_1596_symbol;
              Xexit_1590_predecessors(2) <= word_access_2_1601_symbol;
              Xexit_1590_predecessors(3) <= word_access_3_1606_symbol;
              Xexit_1590_join: join -- 
                port map( -- 
                  preds => Xexit_1590_predecessors,
                  symbol_out => Xexit_1590_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/$exit
            word_access_1588_symbol <= Xexit_1590_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access
          Xexit_1585_symbol <= word_access_1588_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/$exit
          ptr_deref_285_request_1583_symbol <= Xexit_1585_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request
        ptr_deref_285_complete_1611: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete 
          signal ptr_deref_285_complete_1611_start: Boolean;
          signal Xentry_1612_symbol: Boolean;
          signal Xexit_1613_symbol: Boolean;
          signal word_access_1614_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_285_complete_1611_start <= ptr_deref_285_active_x_x1579_symbol; -- control passed to block
          Xentry_1612_symbol  <= ptr_deref_285_complete_1611_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/$entry
          word_access_1614: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access 
            signal word_access_1614_start: Boolean;
            signal Xentry_1615_symbol: Boolean;
            signal Xexit_1616_symbol: Boolean;
            signal word_access_0_1617_symbol : Boolean;
            signal word_access_1_1622_symbol : Boolean;
            signal word_access_2_1627_symbol : Boolean;
            signal word_access_3_1632_symbol : Boolean;
            -- 
          begin -- 
            word_access_1614_start <= Xentry_1612_symbol; -- control passed to block
            Xentry_1615_symbol  <= word_access_1614_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/$entry
            word_access_0_1617: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0 
              signal word_access_0_1617_start: Boolean;
              signal Xentry_1618_symbol: Boolean;
              signal Xexit_1619_symbol: Boolean;
              signal cr_1620_symbol : Boolean;
              signal ca_1621_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1617_start <= Xentry_1615_symbol; -- control passed to block
              Xentry_1618_symbol  <= word_access_0_1617_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/$entry
              cr_1620_symbol <= Xentry_1618_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/cr
              ptr_deref_285_store_0_req_1 <= cr_1620_symbol; -- link to DP
              ca_1621_symbol <= ptr_deref_285_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/ca
              Xexit_1619_symbol <= ca_1621_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/$exit
              word_access_0_1617_symbol <= Xexit_1619_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0
            word_access_1_1622: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_1 
              signal word_access_1_1622_start: Boolean;
              signal Xentry_1623_symbol: Boolean;
              signal Xexit_1624_symbol: Boolean;
              signal cr_1625_symbol : Boolean;
              signal ca_1626_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1622_start <= Xentry_1615_symbol; -- control passed to block
              Xentry_1623_symbol  <= word_access_1_1622_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_1/$entry
              cr_1625_symbol <= Xentry_1623_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_1/cr
              ptr_deref_285_store_1_req_1 <= cr_1625_symbol; -- link to DP
              ca_1626_symbol <= ptr_deref_285_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_1/ca
              Xexit_1624_symbol <= ca_1626_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_1/$exit
              word_access_1_1622_symbol <= Xexit_1624_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_1
            word_access_2_1627: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_2 
              signal word_access_2_1627_start: Boolean;
              signal Xentry_1628_symbol: Boolean;
              signal Xexit_1629_symbol: Boolean;
              signal cr_1630_symbol : Boolean;
              signal ca_1631_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1627_start <= Xentry_1615_symbol; -- control passed to block
              Xentry_1628_symbol  <= word_access_2_1627_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_2/$entry
              cr_1630_symbol <= Xentry_1628_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_2/cr
              ptr_deref_285_store_2_req_1 <= cr_1630_symbol; -- link to DP
              ca_1631_symbol <= ptr_deref_285_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_2/ca
              Xexit_1629_symbol <= ca_1631_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_2/$exit
              word_access_2_1627_symbol <= Xexit_1629_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_2
            word_access_3_1632: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_3 
              signal word_access_3_1632_start: Boolean;
              signal Xentry_1633_symbol: Boolean;
              signal Xexit_1634_symbol: Boolean;
              signal cr_1635_symbol : Boolean;
              signal ca_1636_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1632_start <= Xentry_1615_symbol; -- control passed to block
              Xentry_1633_symbol  <= word_access_3_1632_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_3/$entry
              cr_1635_symbol <= Xentry_1633_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_3/cr
              ptr_deref_285_store_3_req_1 <= cr_1635_symbol; -- link to DP
              ca_1636_symbol <= ptr_deref_285_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_3/ca
              Xexit_1634_symbol <= ca_1636_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_3/$exit
              word_access_3_1632_symbol <= Xexit_1634_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_3
            Xexit_1616_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/$exit 
              signal Xexit_1616_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1616_predecessors(0) <= word_access_0_1617_symbol;
              Xexit_1616_predecessors(1) <= word_access_1_1622_symbol;
              Xexit_1616_predecessors(2) <= word_access_2_1627_symbol;
              Xexit_1616_predecessors(3) <= word_access_3_1632_symbol;
              Xexit_1616_join: join -- 
                port map( -- 
                  preds => Xexit_1616_predecessors,
                  symbol_out => Xexit_1616_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/$exit
            word_access_1614_symbol <= Xexit_1616_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access
          Xexit_1613_symbol <= word_access_1614_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/$exit
          ptr_deref_285_complete_1611_symbol <= Xexit_1613_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete
        assign_stmt_290_active_x_x1637_symbol <= simple_obj_ref_289_complete_1654_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_290_active_
        assign_stmt_290_completed_x_x1638_symbol <= assign_stmt_290_active_x_x1637_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_290_completed_
        simple_obj_ref_289_trigger_x_x1639_symbol <= simple_obj_ref_289_word_address_calculated_1642_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_trigger_
        simple_obj_ref_289_active_x_x1640_symbol <= simple_obj_ref_289_request_1643_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_active_
        simple_obj_ref_289_root_address_calculated_1641_symbol <= Xentry_1543_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_root_address_calculated
        simple_obj_ref_289_word_address_calculated_1642_symbol <= simple_obj_ref_289_root_address_calculated_1641_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_word_address_calculated
        simple_obj_ref_289_request_1643: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request 
          signal simple_obj_ref_289_request_1643_start: Boolean;
          signal Xentry_1644_symbol: Boolean;
          signal Xexit_1645_symbol: Boolean;
          signal word_access_1646_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_289_request_1643_start <= simple_obj_ref_289_trigger_x_x1639_symbol; -- control passed to block
          Xentry_1644_symbol  <= simple_obj_ref_289_request_1643_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/$entry
          word_access_1646: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access 
            signal word_access_1646_start: Boolean;
            signal Xentry_1647_symbol: Boolean;
            signal Xexit_1648_symbol: Boolean;
            signal word_access_0_1649_symbol : Boolean;
            -- 
          begin -- 
            word_access_1646_start <= Xentry_1644_symbol; -- control passed to block
            Xentry_1647_symbol  <= word_access_1646_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/$entry
            word_access_0_1649: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0 
              signal word_access_0_1649_start: Boolean;
              signal Xentry_1650_symbol: Boolean;
              signal Xexit_1651_symbol: Boolean;
              signal rr_1652_symbol : Boolean;
              signal ra_1653_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1649_start <= Xentry_1647_symbol; -- control passed to block
              Xentry_1650_symbol  <= word_access_0_1649_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/$entry
              rr_1652_symbol <= Xentry_1650_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/rr
              simple_obj_ref_289_load_0_req_0 <= rr_1652_symbol; -- link to DP
              ra_1653_symbol <= simple_obj_ref_289_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/ra
              Xexit_1651_symbol <= ra_1653_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/$exit
              word_access_0_1649_symbol <= Xexit_1651_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0
            Xexit_1648_symbol <= word_access_0_1649_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/$exit
            word_access_1646_symbol <= Xexit_1648_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access
          Xexit_1645_symbol <= word_access_1646_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/$exit
          simple_obj_ref_289_request_1643_symbol <= Xexit_1645_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request
        simple_obj_ref_289_complete_1654: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete 
          signal simple_obj_ref_289_complete_1654_start: Boolean;
          signal Xentry_1655_symbol: Boolean;
          signal Xexit_1656_symbol: Boolean;
          signal word_access_1657_symbol : Boolean;
          signal merge_req_1665_symbol : Boolean;
          signal merge_ack_1666_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_289_complete_1654_start <= simple_obj_ref_289_active_x_x1640_symbol; -- control passed to block
          Xentry_1655_symbol  <= simple_obj_ref_289_complete_1654_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/$entry
          word_access_1657: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access 
            signal word_access_1657_start: Boolean;
            signal Xentry_1658_symbol: Boolean;
            signal Xexit_1659_symbol: Boolean;
            signal word_access_0_1660_symbol : Boolean;
            -- 
          begin -- 
            word_access_1657_start <= Xentry_1655_symbol; -- control passed to block
            Xentry_1658_symbol  <= word_access_1657_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/$entry
            word_access_0_1660: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0 
              signal word_access_0_1660_start: Boolean;
              signal Xentry_1661_symbol: Boolean;
              signal Xexit_1662_symbol: Boolean;
              signal cr_1663_symbol : Boolean;
              signal ca_1664_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1660_start <= Xentry_1658_symbol; -- control passed to block
              Xentry_1661_symbol  <= word_access_0_1660_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/$entry
              cr_1663_symbol <= Xentry_1661_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/cr
              simple_obj_ref_289_load_0_req_1 <= cr_1663_symbol; -- link to DP
              ca_1664_symbol <= simple_obj_ref_289_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/ca
              Xexit_1662_symbol <= ca_1664_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/$exit
              word_access_0_1660_symbol <= Xexit_1662_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0
            Xexit_1659_symbol <= word_access_0_1660_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/$exit
            word_access_1657_symbol <= Xexit_1659_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access
          merge_req_1665_symbol <= word_access_1657_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/merge_req
          simple_obj_ref_289_gather_scatter_req_0 <= merge_req_1665_symbol; -- link to DP
          merge_ack_1666_symbol <= simple_obj_ref_289_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/merge_ack
          Xexit_1656_symbol <= merge_ack_1666_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/$exit
          simple_obj_ref_289_complete_1654_symbol <= Xexit_1656_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete
        assign_stmt_297_active_x_x1667_symbol <= binary_296_complete_1681_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_297_active_
        assign_stmt_297_completed_x_x1668_symbol <= assign_stmt_297_active_x_x1667_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_297_completed_
        binary_296_active_x_x1669_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_active_ 
          signal binary_296_active_x_x1669_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_296_active_x_x1669_predecessors(0) <= binary_296_trigger_x_x1670_symbol;
          binary_296_active_x_x1669_predecessors(1) <= type_cast_293_complete_1674_symbol;
          binary_296_active_x_x1669_join: join -- 
            port map( -- 
              preds => binary_296_active_x_x1669_predecessors,
              symbol_out => binary_296_active_x_x1669_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_active_
        binary_296_trigger_x_x1670_symbol <= Xentry_1543_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_trigger_
        type_cast_293_active_x_x1671_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_active_ 
          signal type_cast_293_active_x_x1671_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_293_active_x_x1671_predecessors(0) <= type_cast_293_trigger_x_x1672_symbol;
          type_cast_293_active_x_x1671_predecessors(1) <= simple_obj_ref_292_complete_1673_symbol;
          type_cast_293_active_x_x1671_join: join -- 
            port map( -- 
              preds => type_cast_293_active_x_x1671_predecessors,
              symbol_out => type_cast_293_active_x_x1671_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_active_
        type_cast_293_trigger_x_x1672_symbol <= Xentry_1543_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_trigger_
        simple_obj_ref_292_complete_1673_symbol <= assign_stmt_290_completed_x_x1638_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_292_complete
        type_cast_293_complete_1674: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete 
          signal type_cast_293_complete_1674_start: Boolean;
          signal Xentry_1675_symbol: Boolean;
          signal Xexit_1676_symbol: Boolean;
          signal rr_1677_symbol : Boolean;
          signal ra_1678_symbol : Boolean;
          signal cr_1679_symbol : Boolean;
          signal ca_1680_symbol : Boolean;
          -- 
        begin -- 
          type_cast_293_complete_1674_start <= type_cast_293_active_x_x1671_symbol; -- control passed to block
          Xentry_1675_symbol  <= type_cast_293_complete_1674_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/$entry
          rr_1677_symbol <= Xentry_1675_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/rr
          type_cast_293_inst_req_0 <= rr_1677_symbol; -- link to DP
          ra_1678_symbol <= type_cast_293_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/ra
          cr_1679_symbol <= ra_1678_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/cr
          type_cast_293_inst_req_1 <= cr_1679_symbol; -- link to DP
          ca_1680_symbol <= type_cast_293_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/ca
          Xexit_1676_symbol <= ca_1680_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/$exit
          type_cast_293_complete_1674_symbol <= Xexit_1676_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete
        binary_296_complete_1681: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete 
          signal binary_296_complete_1681_start: Boolean;
          signal Xentry_1682_symbol: Boolean;
          signal Xexit_1683_symbol: Boolean;
          signal rr_1684_symbol : Boolean;
          signal ra_1685_symbol : Boolean;
          signal cr_1686_symbol : Boolean;
          signal ca_1687_symbol : Boolean;
          -- 
        begin -- 
          binary_296_complete_1681_start <= binary_296_active_x_x1669_symbol; -- control passed to block
          Xentry_1682_symbol  <= binary_296_complete_1681_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/$entry
          rr_1684_symbol <= Xentry_1682_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/rr
          binary_296_inst_req_0 <= rr_1684_symbol; -- link to DP
          ra_1685_symbol <= binary_296_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/ra
          cr_1686_symbol <= ra_1685_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/cr
          binary_296_inst_req_1 <= cr_1686_symbol; -- link to DP
          ca_1687_symbol <= binary_296_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/ca
          Xexit_1683_symbol <= ca_1687_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/$exit
          binary_296_complete_1681_symbol <= Xexit_1683_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete
        Xexit_1544_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/$exit 
          signal Xexit_1544_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          Xexit_1544_predecessors(0) <= assign_stmt_287_completed_x_x1576_symbol;
          Xexit_1544_predecessors(1) <= ptr_deref_285_base_address_calculated_1580_symbol;
          Xexit_1544_predecessors(2) <= assign_stmt_297_completed_x_x1668_symbol;
          Xexit_1544_join: join -- 
            port map( -- 
              preds => Xexit_1544_predecessors,
              symbol_out => Xexit_1544_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/$exit
        assign_stmt_283_to_assign_stmt_297_1542_symbol <= Xexit_1544_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297
      if_stmt_298_dead_link_1688: Block -- branch_block_stmt_134/if_stmt_298_dead_link 
        signal if_stmt_298_dead_link_1688_start: Boolean;
        signal Xentry_1689_symbol: Boolean;
        signal Xexit_1690_symbol: Boolean;
        signal dead_transition_1691_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_dead_link_1688_start <= if_stmt_298_x_xentry_x_xx_x652_symbol; -- control passed to block
        Xentry_1689_symbol  <= if_stmt_298_dead_link_1688_start; -- transition branch_block_stmt_134/if_stmt_298_dead_link/$entry
        dead_transition_1691_symbol <= false;
        Xexit_1690_symbol <= dead_transition_1691_symbol; -- transition branch_block_stmt_134/if_stmt_298_dead_link/$exit
        if_stmt_298_dead_link_1688_symbol <= Xexit_1690_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_dead_link
      if_stmt_298_eval_test_1692: Block -- branch_block_stmt_134/if_stmt_298_eval_test 
        signal if_stmt_298_eval_test_1692_start: Boolean;
        signal Xentry_1693_symbol: Boolean;
        signal Xexit_1694_symbol: Boolean;
        signal branch_req_1695_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_eval_test_1692_start <= if_stmt_298_x_xentry_x_xx_x652_symbol; -- control passed to block
        Xentry_1693_symbol  <= if_stmt_298_eval_test_1692_start; -- transition branch_block_stmt_134/if_stmt_298_eval_test/$entry
        branch_req_1695_symbol <= Xentry_1693_symbol; -- transition branch_block_stmt_134/if_stmt_298_eval_test/branch_req
        if_stmt_298_branch_req_0 <= branch_req_1695_symbol; -- link to DP
        Xexit_1694_symbol <= branch_req_1695_symbol; -- transition branch_block_stmt_134/if_stmt_298_eval_test/$exit
        if_stmt_298_eval_test_1692_symbol <= Xexit_1694_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_eval_test
      simple_obj_ref_299_place_1696_symbol  <=  if_stmt_298_eval_test_1692_symbol; -- place branch_block_stmt_134/simple_obj_ref_299_place (optimized away) 
      if_stmt_298_if_link_1697: Block -- branch_block_stmt_134/if_stmt_298_if_link 
        signal if_stmt_298_if_link_1697_start: Boolean;
        signal Xentry_1698_symbol: Boolean;
        signal Xexit_1699_symbol: Boolean;
        signal if_choice_transition_1700_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_if_link_1697_start <= simple_obj_ref_299_place_1696_symbol; -- control passed to block
        Xentry_1698_symbol  <= if_stmt_298_if_link_1697_start; -- transition branch_block_stmt_134/if_stmt_298_if_link/$entry
        if_choice_transition_1700_symbol <= if_stmt_298_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_298_if_link/if_choice_transition
        Xexit_1699_symbol <= if_choice_transition_1700_symbol; -- transition branch_block_stmt_134/if_stmt_298_if_link/$exit
        if_stmt_298_if_link_1697_symbol <= Xexit_1699_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_if_link
      if_stmt_298_else_link_1701: Block -- branch_block_stmt_134/if_stmt_298_else_link 
        signal if_stmt_298_else_link_1701_start: Boolean;
        signal Xentry_1702_symbol: Boolean;
        signal Xexit_1703_symbol: Boolean;
        signal else_choice_transition_1704_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_else_link_1701_start <= simple_obj_ref_299_place_1696_symbol; -- control passed to block
        Xentry_1702_symbol  <= if_stmt_298_else_link_1701_start; -- transition branch_block_stmt_134/if_stmt_298_else_link/$entry
        else_choice_transition_1704_symbol <= if_stmt_298_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_298_else_link/else_choice_transition
        Xexit_1703_symbol <= else_choice_transition_1704_symbol; -- transition branch_block_stmt_134/if_stmt_298_else_link/$exit
        if_stmt_298_else_link_1701_symbol <= Xexit_1703_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_else_link
      bb_5_bb_6_1705_symbol  <=  if_stmt_298_if_link_1697_symbol; -- place branch_block_stmt_134/bb_5_bb_6 (optimized away) 
      bb_5_bb_7_1706_symbol  <=  if_stmt_298_else_link_1701_symbol; -- place branch_block_stmt_134/bb_5_bb_7 (optimized away) 
      assign_stmt_307_to_assign_stmt_319_1707: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319 
        signal assign_stmt_307_to_assign_stmt_319_1707_start: Boolean;
        signal Xentry_1708_symbol: Boolean;
        signal Xexit_1709_symbol: Boolean;
        signal assign_stmt_307_active_x_x1710_symbol : Boolean;
        signal assign_stmt_307_completed_x_x1711_symbol : Boolean;
        signal simple_obj_ref_306_trigger_x_x1712_symbol : Boolean;
        signal simple_obj_ref_306_active_x_x1713_symbol : Boolean;
        signal simple_obj_ref_306_root_address_calculated_1714_symbol : Boolean;
        signal simple_obj_ref_306_word_address_calculated_1715_symbol : Boolean;
        signal simple_obj_ref_306_request_1716_symbol : Boolean;
        signal simple_obj_ref_306_complete_1727_symbol : Boolean;
        signal assign_stmt_312_active_x_x1740_symbol : Boolean;
        signal assign_stmt_312_completed_x_x1741_symbol : Boolean;
        signal array_obj_ref_311_trigger_x_x1742_symbol : Boolean;
        signal array_obj_ref_311_active_x_x1743_symbol : Boolean;
        signal array_obj_ref_311_base_address_calculated_1744_symbol : Boolean;
        signal array_obj_ref_311_root_address_calculated_1745_symbol : Boolean;
        signal array_obj_ref_311_base_address_resized_1746_symbol : Boolean;
        signal array_obj_ref_311_base_addr_resize_1747_symbol : Boolean;
        signal array_obj_ref_311_base_plus_offset_1752_symbol : Boolean;
        signal array_obj_ref_311_complete_1757_symbol : Boolean;
        signal assign_stmt_316_active_x_x1762_symbol : Boolean;
        signal assign_stmt_316_completed_x_x1763_symbol : Boolean;
        signal ptr_deref_315_trigger_x_x1764_symbol : Boolean;
        signal ptr_deref_315_active_x_x1765_symbol : Boolean;
        signal ptr_deref_315_base_address_calculated_1766_symbol : Boolean;
        signal simple_obj_ref_314_complete_1767_symbol : Boolean;
        signal ptr_deref_315_root_address_calculated_1768_symbol : Boolean;
        signal ptr_deref_315_word_address_calculated_1769_symbol : Boolean;
        signal ptr_deref_315_base_address_resized_1770_symbol : Boolean;
        signal ptr_deref_315_base_addr_resize_1771_symbol : Boolean;
        signal ptr_deref_315_base_plus_offset_1776_symbol : Boolean;
        signal ptr_deref_315_word_addrgen_1781_symbol : Boolean;
        signal ptr_deref_315_request_1812_symbol : Boolean;
        signal ptr_deref_315_complete_1838_symbol : Boolean;
        signal assign_stmt_319_active_x_x1866_symbol : Boolean;
        signal assign_stmt_319_completed_x_x1867_symbol : Boolean;
        signal simple_obj_ref_318_complete_1868_symbol : Boolean;
        signal simple_obj_ref_317_trigger_x_x1869_symbol : Boolean;
        signal simple_obj_ref_317_active_x_x1870_symbol : Boolean;
        signal simple_obj_ref_317_root_address_calculated_1871_symbol : Boolean;
        signal simple_obj_ref_317_word_address_calculated_1872_symbol : Boolean;
        signal simple_obj_ref_317_request_1873_symbol : Boolean;
        signal simple_obj_ref_317_complete_1886_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_307_to_assign_stmt_319_1707_start <= assign_stmt_307_to_assign_stmt_319_x_xentry_x_xx_x656_symbol; -- control passed to block
        Xentry_1708_symbol  <= assign_stmt_307_to_assign_stmt_319_1707_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/$entry
        assign_stmt_307_active_x_x1710_symbol <= simple_obj_ref_306_complete_1727_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_307_active_
        assign_stmt_307_completed_x_x1711_symbol <= assign_stmt_307_active_x_x1710_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_307_completed_
        simple_obj_ref_306_trigger_x_x1712_symbol <= simple_obj_ref_306_word_address_calculated_1715_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_trigger_
        simple_obj_ref_306_active_x_x1713_symbol <= simple_obj_ref_306_request_1716_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_active_
        simple_obj_ref_306_root_address_calculated_1714_symbol <= Xentry_1708_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_root_address_calculated
        simple_obj_ref_306_word_address_calculated_1715_symbol <= simple_obj_ref_306_root_address_calculated_1714_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_word_address_calculated
        simple_obj_ref_306_request_1716: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request 
          signal simple_obj_ref_306_request_1716_start: Boolean;
          signal Xentry_1717_symbol: Boolean;
          signal Xexit_1718_symbol: Boolean;
          signal word_access_1719_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_306_request_1716_start <= simple_obj_ref_306_trigger_x_x1712_symbol; -- control passed to block
          Xentry_1717_symbol  <= simple_obj_ref_306_request_1716_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/$entry
          word_access_1719: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access 
            signal word_access_1719_start: Boolean;
            signal Xentry_1720_symbol: Boolean;
            signal Xexit_1721_symbol: Boolean;
            signal word_access_0_1722_symbol : Boolean;
            -- 
          begin -- 
            word_access_1719_start <= Xentry_1717_symbol; -- control passed to block
            Xentry_1720_symbol  <= word_access_1719_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/$entry
            word_access_0_1722: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0 
              signal word_access_0_1722_start: Boolean;
              signal Xentry_1723_symbol: Boolean;
              signal Xexit_1724_symbol: Boolean;
              signal rr_1725_symbol : Boolean;
              signal ra_1726_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1722_start <= Xentry_1720_symbol; -- control passed to block
              Xentry_1723_symbol  <= word_access_0_1722_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/$entry
              rr_1725_symbol <= Xentry_1723_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/rr
              simple_obj_ref_306_load_0_req_0 <= rr_1725_symbol; -- link to DP
              ra_1726_symbol <= simple_obj_ref_306_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/ra
              Xexit_1724_symbol <= ra_1726_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/$exit
              word_access_0_1722_symbol <= Xexit_1724_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0
            Xexit_1721_symbol <= word_access_0_1722_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/$exit
            word_access_1719_symbol <= Xexit_1721_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access
          Xexit_1718_symbol <= word_access_1719_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/$exit
          simple_obj_ref_306_request_1716_symbol <= Xexit_1718_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request
        simple_obj_ref_306_complete_1727: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete 
          signal simple_obj_ref_306_complete_1727_start: Boolean;
          signal Xentry_1728_symbol: Boolean;
          signal Xexit_1729_symbol: Boolean;
          signal word_access_1730_symbol : Boolean;
          signal merge_req_1738_symbol : Boolean;
          signal merge_ack_1739_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_306_complete_1727_start <= simple_obj_ref_306_active_x_x1713_symbol; -- control passed to block
          Xentry_1728_symbol  <= simple_obj_ref_306_complete_1727_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/$entry
          word_access_1730: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access 
            signal word_access_1730_start: Boolean;
            signal Xentry_1731_symbol: Boolean;
            signal Xexit_1732_symbol: Boolean;
            signal word_access_0_1733_symbol : Boolean;
            -- 
          begin -- 
            word_access_1730_start <= Xentry_1728_symbol; -- control passed to block
            Xentry_1731_symbol  <= word_access_1730_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/$entry
            word_access_0_1733: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0 
              signal word_access_0_1733_start: Boolean;
              signal Xentry_1734_symbol: Boolean;
              signal Xexit_1735_symbol: Boolean;
              signal cr_1736_symbol : Boolean;
              signal ca_1737_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1733_start <= Xentry_1731_symbol; -- control passed to block
              Xentry_1734_symbol  <= word_access_0_1733_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/$entry
              cr_1736_symbol <= Xentry_1734_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/cr
              simple_obj_ref_306_load_0_req_1 <= cr_1736_symbol; -- link to DP
              ca_1737_symbol <= simple_obj_ref_306_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/ca
              Xexit_1735_symbol <= ca_1737_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/$exit
              word_access_0_1733_symbol <= Xexit_1735_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0
            Xexit_1732_symbol <= word_access_0_1733_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/$exit
            word_access_1730_symbol <= Xexit_1732_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access
          merge_req_1738_symbol <= word_access_1730_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/merge_req
          simple_obj_ref_306_gather_scatter_req_0 <= merge_req_1738_symbol; -- link to DP
          merge_ack_1739_symbol <= simple_obj_ref_306_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/merge_ack
          Xexit_1729_symbol <= merge_ack_1739_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/$exit
          simple_obj_ref_306_complete_1727_symbol <= Xexit_1729_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete
        assign_stmt_312_active_x_x1740_symbol <= array_obj_ref_311_complete_1757_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_312_active_
        assign_stmt_312_completed_x_x1741_symbol <= assign_stmt_312_active_x_x1740_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_312_completed_
        array_obj_ref_311_trigger_x_x1742_symbol <= Xentry_1708_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_trigger_
        array_obj_ref_311_active_x_x1743_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_active_ 
          signal array_obj_ref_311_active_x_x1743_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_311_active_x_x1743_predecessors(0) <= array_obj_ref_311_trigger_x_x1742_symbol;
          array_obj_ref_311_active_x_x1743_predecessors(1) <= array_obj_ref_311_root_address_calculated_1745_symbol;
          array_obj_ref_311_active_x_x1743_join: join -- 
            port map( -- 
              preds => array_obj_ref_311_active_x_x1743_predecessors,
              symbol_out => array_obj_ref_311_active_x_x1743_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_active_
        array_obj_ref_311_base_address_calculated_1744_symbol <= assign_stmt_307_completed_x_x1711_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_address_calculated
        array_obj_ref_311_root_address_calculated_1745_symbol <= array_obj_ref_311_base_plus_offset_1752_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_root_address_calculated
        array_obj_ref_311_base_address_resized_1746_symbol <= array_obj_ref_311_base_addr_resize_1747_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_address_resized
        array_obj_ref_311_base_addr_resize_1747: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize 
          signal array_obj_ref_311_base_addr_resize_1747_start: Boolean;
          signal Xentry_1748_symbol: Boolean;
          signal Xexit_1749_symbol: Boolean;
          signal base_resize_req_1750_symbol : Boolean;
          signal base_resize_ack_1751_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_311_base_addr_resize_1747_start <= array_obj_ref_311_base_address_calculated_1744_symbol; -- control passed to block
          Xentry_1748_symbol  <= array_obj_ref_311_base_addr_resize_1747_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/$entry
          base_resize_req_1750_symbol <= Xentry_1748_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/base_resize_req
          array_obj_ref_311_base_resize_req_0 <= base_resize_req_1750_symbol; -- link to DP
          base_resize_ack_1751_symbol <= array_obj_ref_311_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/base_resize_ack
          Xexit_1749_symbol <= base_resize_ack_1751_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/$exit
          array_obj_ref_311_base_addr_resize_1747_symbol <= Xexit_1749_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize
        array_obj_ref_311_base_plus_offset_1752: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset 
          signal array_obj_ref_311_base_plus_offset_1752_start: Boolean;
          signal Xentry_1753_symbol: Boolean;
          signal Xexit_1754_symbol: Boolean;
          signal sum_rename_req_1755_symbol : Boolean;
          signal sum_rename_ack_1756_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_311_base_plus_offset_1752_start <= array_obj_ref_311_base_address_resized_1746_symbol; -- control passed to block
          Xentry_1753_symbol  <= array_obj_ref_311_base_plus_offset_1752_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/$entry
          sum_rename_req_1755_symbol <= Xentry_1753_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/sum_rename_req
          array_obj_ref_311_root_address_inst_req_0 <= sum_rename_req_1755_symbol; -- link to DP
          sum_rename_ack_1756_symbol <= array_obj_ref_311_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/sum_rename_ack
          Xexit_1754_symbol <= sum_rename_ack_1756_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/$exit
          array_obj_ref_311_base_plus_offset_1752_symbol <= Xexit_1754_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset
        array_obj_ref_311_complete_1757: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete 
          signal array_obj_ref_311_complete_1757_start: Boolean;
          signal Xentry_1758_symbol: Boolean;
          signal Xexit_1759_symbol: Boolean;
          signal final_reg_req_1760_symbol : Boolean;
          signal final_reg_ack_1761_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_311_complete_1757_start <= array_obj_ref_311_active_x_x1743_symbol; -- control passed to block
          Xentry_1758_symbol  <= array_obj_ref_311_complete_1757_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/$entry
          final_reg_req_1760_symbol <= Xentry_1758_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/final_reg_req
          array_obj_ref_311_final_reg_req_0 <= final_reg_req_1760_symbol; -- link to DP
          final_reg_ack_1761_symbol <= array_obj_ref_311_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/final_reg_ack
          Xexit_1759_symbol <= final_reg_ack_1761_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/$exit
          array_obj_ref_311_complete_1757_symbol <= Xexit_1759_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete
        assign_stmt_316_active_x_x1762_symbol <= ptr_deref_315_complete_1838_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_316_active_
        assign_stmt_316_completed_x_x1763_symbol <= assign_stmt_316_active_x_x1762_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_316_completed_
        ptr_deref_315_trigger_x_x1764_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_trigger_ 
          signal ptr_deref_315_trigger_x_x1764_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_315_trigger_x_x1764_predecessors(0) <= ptr_deref_315_word_address_calculated_1769_symbol;
          ptr_deref_315_trigger_x_x1764_predecessors(1) <= ptr_deref_315_base_address_calculated_1766_symbol;
          ptr_deref_315_trigger_x_x1764_join: join -- 
            port map( -- 
              preds => ptr_deref_315_trigger_x_x1764_predecessors,
              symbol_out => ptr_deref_315_trigger_x_x1764_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_trigger_
        ptr_deref_315_active_x_x1765_symbol <= ptr_deref_315_request_1812_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_active_
        ptr_deref_315_base_address_calculated_1766_symbol <= simple_obj_ref_314_complete_1767_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_address_calculated
        simple_obj_ref_314_complete_1767_symbol <= assign_stmt_312_completed_x_x1741_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_314_complete
        ptr_deref_315_root_address_calculated_1768_symbol <= ptr_deref_315_base_plus_offset_1776_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_root_address_calculated
        ptr_deref_315_word_address_calculated_1769_symbol <= ptr_deref_315_word_addrgen_1781_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_address_calculated
        ptr_deref_315_base_address_resized_1770_symbol <= ptr_deref_315_base_addr_resize_1771_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_address_resized
        ptr_deref_315_base_addr_resize_1771: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize 
          signal ptr_deref_315_base_addr_resize_1771_start: Boolean;
          signal Xentry_1772_symbol: Boolean;
          signal Xexit_1773_symbol: Boolean;
          signal base_resize_req_1774_symbol : Boolean;
          signal base_resize_ack_1775_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_base_addr_resize_1771_start <= ptr_deref_315_base_address_calculated_1766_symbol; -- control passed to block
          Xentry_1772_symbol  <= ptr_deref_315_base_addr_resize_1771_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/$entry
          base_resize_req_1774_symbol <= Xentry_1772_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/base_resize_req
          ptr_deref_315_base_resize_req_0 <= base_resize_req_1774_symbol; -- link to DP
          base_resize_ack_1775_symbol <= ptr_deref_315_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/base_resize_ack
          Xexit_1773_symbol <= base_resize_ack_1775_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/$exit
          ptr_deref_315_base_addr_resize_1771_symbol <= Xexit_1773_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize
        ptr_deref_315_base_plus_offset_1776: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset 
          signal ptr_deref_315_base_plus_offset_1776_start: Boolean;
          signal Xentry_1777_symbol: Boolean;
          signal Xexit_1778_symbol: Boolean;
          signal sum_rename_req_1779_symbol : Boolean;
          signal sum_rename_ack_1780_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_base_plus_offset_1776_start <= ptr_deref_315_base_address_resized_1770_symbol; -- control passed to block
          Xentry_1777_symbol  <= ptr_deref_315_base_plus_offset_1776_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/$entry
          sum_rename_req_1779_symbol <= Xentry_1777_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/sum_rename_req
          ptr_deref_315_root_address_inst_req_0 <= sum_rename_req_1779_symbol; -- link to DP
          sum_rename_ack_1780_symbol <= ptr_deref_315_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/sum_rename_ack
          Xexit_1778_symbol <= sum_rename_ack_1780_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/$exit
          ptr_deref_315_base_plus_offset_1776_symbol <= Xexit_1778_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset
        ptr_deref_315_word_addrgen_1781: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen 
          signal ptr_deref_315_word_addrgen_1781_start: Boolean;
          signal Xentry_1782_symbol: Boolean;
          signal Xexit_1783_symbol: Boolean;
          signal word_0_1784_symbol : Boolean;
          signal word_1_1791_symbol : Boolean;
          signal word_2_1798_symbol : Boolean;
          signal word_3_1805_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_word_addrgen_1781_start <= ptr_deref_315_root_address_calculated_1768_symbol; -- control passed to block
          Xentry_1782_symbol  <= ptr_deref_315_word_addrgen_1781_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/$entry
          word_0_1784: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0 
            signal word_0_1784_start: Boolean;
            signal Xentry_1785_symbol: Boolean;
            signal Xexit_1786_symbol: Boolean;
            signal rr_1787_symbol : Boolean;
            signal ra_1788_symbol : Boolean;
            signal cr_1789_symbol : Boolean;
            signal ca_1790_symbol : Boolean;
            -- 
          begin -- 
            word_0_1784_start <= Xentry_1782_symbol; -- control passed to block
            Xentry_1785_symbol  <= word_0_1784_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0/$entry
            rr_1787_symbol <= Xentry_1785_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0/rr
            ptr_deref_315_addr_0_req_0 <= rr_1787_symbol; -- link to DP
            ra_1788_symbol <= ptr_deref_315_addr_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0/ra
            cr_1789_symbol <= ra_1788_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0/cr
            ptr_deref_315_addr_0_req_1 <= cr_1789_symbol; -- link to DP
            ca_1790_symbol <= ptr_deref_315_addr_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0/ca
            Xexit_1786_symbol <= ca_1790_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0/$exit
            word_0_1784_symbol <= Xexit_1786_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_0
          word_1_1791: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1 
            signal word_1_1791_start: Boolean;
            signal Xentry_1792_symbol: Boolean;
            signal Xexit_1793_symbol: Boolean;
            signal rr_1794_symbol : Boolean;
            signal ra_1795_symbol : Boolean;
            signal cr_1796_symbol : Boolean;
            signal ca_1797_symbol : Boolean;
            -- 
          begin -- 
            word_1_1791_start <= Xentry_1782_symbol; -- control passed to block
            Xentry_1792_symbol  <= word_1_1791_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1/$entry
            rr_1794_symbol <= Xentry_1792_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1/rr
            ptr_deref_315_addr_1_req_0 <= rr_1794_symbol; -- link to DP
            ra_1795_symbol <= ptr_deref_315_addr_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1/ra
            cr_1796_symbol <= ra_1795_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1/cr
            ptr_deref_315_addr_1_req_1 <= cr_1796_symbol; -- link to DP
            ca_1797_symbol <= ptr_deref_315_addr_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1/ca
            Xexit_1793_symbol <= ca_1797_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1/$exit
            word_1_1791_symbol <= Xexit_1793_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_1
          word_2_1798: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2 
            signal word_2_1798_start: Boolean;
            signal Xentry_1799_symbol: Boolean;
            signal Xexit_1800_symbol: Boolean;
            signal rr_1801_symbol : Boolean;
            signal ra_1802_symbol : Boolean;
            signal cr_1803_symbol : Boolean;
            signal ca_1804_symbol : Boolean;
            -- 
          begin -- 
            word_2_1798_start <= Xentry_1782_symbol; -- control passed to block
            Xentry_1799_symbol  <= word_2_1798_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2/$entry
            rr_1801_symbol <= Xentry_1799_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2/rr
            ptr_deref_315_addr_2_req_0 <= rr_1801_symbol; -- link to DP
            ra_1802_symbol <= ptr_deref_315_addr_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2/ra
            cr_1803_symbol <= ra_1802_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2/cr
            ptr_deref_315_addr_2_req_1 <= cr_1803_symbol; -- link to DP
            ca_1804_symbol <= ptr_deref_315_addr_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2/ca
            Xexit_1800_symbol <= ca_1804_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2/$exit
            word_2_1798_symbol <= Xexit_1800_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_2
          word_3_1805: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3 
            signal word_3_1805_start: Boolean;
            signal Xentry_1806_symbol: Boolean;
            signal Xexit_1807_symbol: Boolean;
            signal rr_1808_symbol : Boolean;
            signal ra_1809_symbol : Boolean;
            signal cr_1810_symbol : Boolean;
            signal ca_1811_symbol : Boolean;
            -- 
          begin -- 
            word_3_1805_start <= Xentry_1782_symbol; -- control passed to block
            Xentry_1806_symbol  <= word_3_1805_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3/$entry
            rr_1808_symbol <= Xentry_1806_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3/rr
            ptr_deref_315_addr_3_req_0 <= rr_1808_symbol; -- link to DP
            ra_1809_symbol <= ptr_deref_315_addr_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3/ra
            cr_1810_symbol <= ra_1809_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3/cr
            ptr_deref_315_addr_3_req_1 <= cr_1810_symbol; -- link to DP
            ca_1811_symbol <= ptr_deref_315_addr_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3/ca
            Xexit_1807_symbol <= ca_1811_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3/$exit
            word_3_1805_symbol <= Xexit_1807_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/word_3
          Xexit_1783_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/$exit 
            signal Xexit_1783_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_1783_predecessors(0) <= word_0_1784_symbol;
            Xexit_1783_predecessors(1) <= word_1_1791_symbol;
            Xexit_1783_predecessors(2) <= word_2_1798_symbol;
            Xexit_1783_predecessors(3) <= word_3_1805_symbol;
            Xexit_1783_join: join -- 
              port map( -- 
                preds => Xexit_1783_predecessors,
                symbol_out => Xexit_1783_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/$exit
          ptr_deref_315_word_addrgen_1781_symbol <= Xexit_1783_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen
        ptr_deref_315_request_1812: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request 
          signal ptr_deref_315_request_1812_start: Boolean;
          signal Xentry_1813_symbol: Boolean;
          signal Xexit_1814_symbol: Boolean;
          signal word_access_1815_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_request_1812_start <= ptr_deref_315_trigger_x_x1764_symbol; -- control passed to block
          Xentry_1813_symbol  <= ptr_deref_315_request_1812_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/$entry
          word_access_1815: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access 
            signal word_access_1815_start: Boolean;
            signal Xentry_1816_symbol: Boolean;
            signal Xexit_1817_symbol: Boolean;
            signal word_access_0_1818_symbol : Boolean;
            signal word_access_1_1823_symbol : Boolean;
            signal word_access_2_1828_symbol : Boolean;
            signal word_access_3_1833_symbol : Boolean;
            -- 
          begin -- 
            word_access_1815_start <= Xentry_1813_symbol; -- control passed to block
            Xentry_1816_symbol  <= word_access_1815_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/$entry
            word_access_0_1818: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0 
              signal word_access_0_1818_start: Boolean;
              signal Xentry_1819_symbol: Boolean;
              signal Xexit_1820_symbol: Boolean;
              signal rr_1821_symbol : Boolean;
              signal ra_1822_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1818_start <= Xentry_1816_symbol; -- control passed to block
              Xentry_1819_symbol  <= word_access_0_1818_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/$entry
              rr_1821_symbol <= Xentry_1819_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/rr
              ptr_deref_315_load_0_req_0 <= rr_1821_symbol; -- link to DP
              ra_1822_symbol <= ptr_deref_315_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/ra
              Xexit_1820_symbol <= ra_1822_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/$exit
              word_access_0_1818_symbol <= Xexit_1820_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0
            word_access_1_1823: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_1 
              signal word_access_1_1823_start: Boolean;
              signal Xentry_1824_symbol: Boolean;
              signal Xexit_1825_symbol: Boolean;
              signal rr_1826_symbol : Boolean;
              signal ra_1827_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1823_start <= Xentry_1816_symbol; -- control passed to block
              Xentry_1824_symbol  <= word_access_1_1823_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_1/$entry
              rr_1826_symbol <= Xentry_1824_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_1/rr
              ptr_deref_315_load_1_req_0 <= rr_1826_symbol; -- link to DP
              ra_1827_symbol <= ptr_deref_315_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_1/ra
              Xexit_1825_symbol <= ra_1827_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_1/$exit
              word_access_1_1823_symbol <= Xexit_1825_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_1
            word_access_2_1828: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_2 
              signal word_access_2_1828_start: Boolean;
              signal Xentry_1829_symbol: Boolean;
              signal Xexit_1830_symbol: Boolean;
              signal rr_1831_symbol : Boolean;
              signal ra_1832_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1828_start <= Xentry_1816_symbol; -- control passed to block
              Xentry_1829_symbol  <= word_access_2_1828_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_2/$entry
              rr_1831_symbol <= Xentry_1829_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_2/rr
              ptr_deref_315_load_2_req_0 <= rr_1831_symbol; -- link to DP
              ra_1832_symbol <= ptr_deref_315_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_2/ra
              Xexit_1830_symbol <= ra_1832_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_2/$exit
              word_access_2_1828_symbol <= Xexit_1830_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_2
            word_access_3_1833: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_3 
              signal word_access_3_1833_start: Boolean;
              signal Xentry_1834_symbol: Boolean;
              signal Xexit_1835_symbol: Boolean;
              signal rr_1836_symbol : Boolean;
              signal ra_1837_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1833_start <= Xentry_1816_symbol; -- control passed to block
              Xentry_1834_symbol  <= word_access_3_1833_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_3/$entry
              rr_1836_symbol <= Xentry_1834_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_3/rr
              ptr_deref_315_load_3_req_0 <= rr_1836_symbol; -- link to DP
              ra_1837_symbol <= ptr_deref_315_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_3/ra
              Xexit_1835_symbol <= ra_1837_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_3/$exit
              word_access_3_1833_symbol <= Xexit_1835_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_3
            Xexit_1817_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/$exit 
              signal Xexit_1817_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1817_predecessors(0) <= word_access_0_1818_symbol;
              Xexit_1817_predecessors(1) <= word_access_1_1823_symbol;
              Xexit_1817_predecessors(2) <= word_access_2_1828_symbol;
              Xexit_1817_predecessors(3) <= word_access_3_1833_symbol;
              Xexit_1817_join: join -- 
                port map( -- 
                  preds => Xexit_1817_predecessors,
                  symbol_out => Xexit_1817_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/$exit
            word_access_1815_symbol <= Xexit_1817_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access
          Xexit_1814_symbol <= word_access_1815_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/$exit
          ptr_deref_315_request_1812_symbol <= Xexit_1814_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request
        ptr_deref_315_complete_1838: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete 
          signal ptr_deref_315_complete_1838_start: Boolean;
          signal Xentry_1839_symbol: Boolean;
          signal Xexit_1840_symbol: Boolean;
          signal word_access_1841_symbol : Boolean;
          signal merge_req_1864_symbol : Boolean;
          signal merge_ack_1865_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_complete_1838_start <= ptr_deref_315_active_x_x1765_symbol; -- control passed to block
          Xentry_1839_symbol  <= ptr_deref_315_complete_1838_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/$entry
          word_access_1841: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access 
            signal word_access_1841_start: Boolean;
            signal Xentry_1842_symbol: Boolean;
            signal Xexit_1843_symbol: Boolean;
            signal word_access_0_1844_symbol : Boolean;
            signal word_access_1_1849_symbol : Boolean;
            signal word_access_2_1854_symbol : Boolean;
            signal word_access_3_1859_symbol : Boolean;
            -- 
          begin -- 
            word_access_1841_start <= Xentry_1839_symbol; -- control passed to block
            Xentry_1842_symbol  <= word_access_1841_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/$entry
            word_access_0_1844: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0 
              signal word_access_0_1844_start: Boolean;
              signal Xentry_1845_symbol: Boolean;
              signal Xexit_1846_symbol: Boolean;
              signal cr_1847_symbol : Boolean;
              signal ca_1848_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1844_start <= Xentry_1842_symbol; -- control passed to block
              Xentry_1845_symbol  <= word_access_0_1844_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/$entry
              cr_1847_symbol <= Xentry_1845_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/cr
              ptr_deref_315_load_0_req_1 <= cr_1847_symbol; -- link to DP
              ca_1848_symbol <= ptr_deref_315_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/ca
              Xexit_1846_symbol <= ca_1848_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/$exit
              word_access_0_1844_symbol <= Xexit_1846_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0
            word_access_1_1849: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_1 
              signal word_access_1_1849_start: Boolean;
              signal Xentry_1850_symbol: Boolean;
              signal Xexit_1851_symbol: Boolean;
              signal cr_1852_symbol : Boolean;
              signal ca_1853_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1849_start <= Xentry_1842_symbol; -- control passed to block
              Xentry_1850_symbol  <= word_access_1_1849_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_1/$entry
              cr_1852_symbol <= Xentry_1850_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_1/cr
              ptr_deref_315_load_1_req_1 <= cr_1852_symbol; -- link to DP
              ca_1853_symbol <= ptr_deref_315_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_1/ca
              Xexit_1851_symbol <= ca_1853_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_1/$exit
              word_access_1_1849_symbol <= Xexit_1851_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_1
            word_access_2_1854: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_2 
              signal word_access_2_1854_start: Boolean;
              signal Xentry_1855_symbol: Boolean;
              signal Xexit_1856_symbol: Boolean;
              signal cr_1857_symbol : Boolean;
              signal ca_1858_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1854_start <= Xentry_1842_symbol; -- control passed to block
              Xentry_1855_symbol  <= word_access_2_1854_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_2/$entry
              cr_1857_symbol <= Xentry_1855_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_2/cr
              ptr_deref_315_load_2_req_1 <= cr_1857_symbol; -- link to DP
              ca_1858_symbol <= ptr_deref_315_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_2/ca
              Xexit_1856_symbol <= ca_1858_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_2/$exit
              word_access_2_1854_symbol <= Xexit_1856_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_2
            word_access_3_1859: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_3 
              signal word_access_3_1859_start: Boolean;
              signal Xentry_1860_symbol: Boolean;
              signal Xexit_1861_symbol: Boolean;
              signal cr_1862_symbol : Boolean;
              signal ca_1863_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1859_start <= Xentry_1842_symbol; -- control passed to block
              Xentry_1860_symbol  <= word_access_3_1859_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_3/$entry
              cr_1862_symbol <= Xentry_1860_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_3/cr
              ptr_deref_315_load_3_req_1 <= cr_1862_symbol; -- link to DP
              ca_1863_symbol <= ptr_deref_315_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_3/ca
              Xexit_1861_symbol <= ca_1863_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_3/$exit
              word_access_3_1859_symbol <= Xexit_1861_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_3
            Xexit_1843_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/$exit 
              signal Xexit_1843_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1843_predecessors(0) <= word_access_0_1844_symbol;
              Xexit_1843_predecessors(1) <= word_access_1_1849_symbol;
              Xexit_1843_predecessors(2) <= word_access_2_1854_symbol;
              Xexit_1843_predecessors(3) <= word_access_3_1859_symbol;
              Xexit_1843_join: join -- 
                port map( -- 
                  preds => Xexit_1843_predecessors,
                  symbol_out => Xexit_1843_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/$exit
            word_access_1841_symbol <= Xexit_1843_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access
          merge_req_1864_symbol <= word_access_1841_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/merge_req
          ptr_deref_315_gather_scatter_req_0 <= merge_req_1864_symbol; -- link to DP
          merge_ack_1865_symbol <= ptr_deref_315_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/merge_ack
          Xexit_1840_symbol <= merge_ack_1865_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/$exit
          ptr_deref_315_complete_1838_symbol <= Xexit_1840_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete
        assign_stmt_319_active_x_x1866_symbol <= simple_obj_ref_318_complete_1868_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_319_active_
        assign_stmt_319_completed_x_x1867_symbol <= simple_obj_ref_317_complete_1886_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_319_completed_
        simple_obj_ref_318_complete_1868_symbol <= assign_stmt_316_completed_x_x1763_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_318_complete
        simple_obj_ref_317_trigger_x_x1869_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_trigger_ 
          signal simple_obj_ref_317_trigger_x_x1869_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          simple_obj_ref_317_trigger_x_x1869_predecessors(0) <= simple_obj_ref_317_word_address_calculated_1872_symbol;
          simple_obj_ref_317_trigger_x_x1869_predecessors(1) <= assign_stmt_319_active_x_x1866_symbol;
          simple_obj_ref_317_trigger_x_x1869_predecessors(2) <= simple_obj_ref_306_active_x_x1713_symbol;
          simple_obj_ref_317_trigger_x_x1869_join: join -- 
            port map( -- 
              preds => simple_obj_ref_317_trigger_x_x1869_predecessors,
              symbol_out => simple_obj_ref_317_trigger_x_x1869_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_trigger_
        simple_obj_ref_317_active_x_x1870_symbol <= simple_obj_ref_317_request_1873_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_active_
        simple_obj_ref_317_root_address_calculated_1871_symbol <= Xentry_1708_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_root_address_calculated
        simple_obj_ref_317_word_address_calculated_1872_symbol <= simple_obj_ref_317_root_address_calculated_1871_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_word_address_calculated
        simple_obj_ref_317_request_1873: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request 
          signal simple_obj_ref_317_request_1873_start: Boolean;
          signal Xentry_1874_symbol: Boolean;
          signal Xexit_1875_symbol: Boolean;
          signal split_req_1876_symbol : Boolean;
          signal split_ack_1877_symbol : Boolean;
          signal word_access_1878_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_317_request_1873_start <= simple_obj_ref_317_trigger_x_x1869_symbol; -- control passed to block
          Xentry_1874_symbol  <= simple_obj_ref_317_request_1873_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/$entry
          split_req_1876_symbol <= Xentry_1874_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/split_req
          simple_obj_ref_317_gather_scatter_req_0 <= split_req_1876_symbol; -- link to DP
          split_ack_1877_symbol <= simple_obj_ref_317_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/split_ack
          word_access_1878: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access 
            signal word_access_1878_start: Boolean;
            signal Xentry_1879_symbol: Boolean;
            signal Xexit_1880_symbol: Boolean;
            signal word_access_0_1881_symbol : Boolean;
            -- 
          begin -- 
            word_access_1878_start <= split_ack_1877_symbol; -- control passed to block
            Xentry_1879_symbol  <= word_access_1878_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/$entry
            word_access_0_1881: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0 
              signal word_access_0_1881_start: Boolean;
              signal Xentry_1882_symbol: Boolean;
              signal Xexit_1883_symbol: Boolean;
              signal rr_1884_symbol : Boolean;
              signal ra_1885_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1881_start <= Xentry_1879_symbol; -- control passed to block
              Xentry_1882_symbol  <= word_access_0_1881_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/$entry
              rr_1884_symbol <= Xentry_1882_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/rr
              simple_obj_ref_317_store_0_req_0 <= rr_1884_symbol; -- link to DP
              ra_1885_symbol <= simple_obj_ref_317_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/ra
              Xexit_1883_symbol <= ra_1885_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/$exit
              word_access_0_1881_symbol <= Xexit_1883_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0
            Xexit_1880_symbol <= word_access_0_1881_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/$exit
            word_access_1878_symbol <= Xexit_1880_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access
          Xexit_1875_symbol <= word_access_1878_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/$exit
          simple_obj_ref_317_request_1873_symbol <= Xexit_1875_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request
        simple_obj_ref_317_complete_1886: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete 
          signal simple_obj_ref_317_complete_1886_start: Boolean;
          signal Xentry_1887_symbol: Boolean;
          signal Xexit_1888_symbol: Boolean;
          signal word_access_1889_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_317_complete_1886_start <= simple_obj_ref_317_active_x_x1870_symbol; -- control passed to block
          Xentry_1887_symbol  <= simple_obj_ref_317_complete_1886_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/$entry
          word_access_1889: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access 
            signal word_access_1889_start: Boolean;
            signal Xentry_1890_symbol: Boolean;
            signal Xexit_1891_symbol: Boolean;
            signal word_access_0_1892_symbol : Boolean;
            -- 
          begin -- 
            word_access_1889_start <= Xentry_1887_symbol; -- control passed to block
            Xentry_1890_symbol  <= word_access_1889_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/$entry
            word_access_0_1892: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0 
              signal word_access_0_1892_start: Boolean;
              signal Xentry_1893_symbol: Boolean;
              signal Xexit_1894_symbol: Boolean;
              signal cr_1895_symbol : Boolean;
              signal ca_1896_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1892_start <= Xentry_1890_symbol; -- control passed to block
              Xentry_1893_symbol  <= word_access_0_1892_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/$entry
              cr_1895_symbol <= Xentry_1893_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/cr
              simple_obj_ref_317_store_0_req_1 <= cr_1895_symbol; -- link to DP
              ca_1896_symbol <= simple_obj_ref_317_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/ca
              Xexit_1894_symbol <= ca_1896_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/$exit
              word_access_0_1892_symbol <= Xexit_1894_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0
            Xexit_1891_symbol <= word_access_0_1892_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/$exit
            word_access_1889_symbol <= Xexit_1891_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access
          Xexit_1888_symbol <= word_access_1889_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/$exit
          simple_obj_ref_317_complete_1886_symbol <= Xexit_1888_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete
        Xexit_1709_symbol <= assign_stmt_319_completed_x_x1867_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/$exit
        assign_stmt_307_to_assign_stmt_319_1707_symbol <= Xexit_1709_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319
      assign_stmt_325_to_assign_stmt_334_1897: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334 
        signal assign_stmt_325_to_assign_stmt_334_1897_start: Boolean;
        signal Xentry_1898_symbol: Boolean;
        signal Xexit_1899_symbol: Boolean;
        signal assign_stmt_325_active_x_x1900_symbol : Boolean;
        signal assign_stmt_325_completed_x_x1901_symbol : Boolean;
        signal ptr_deref_324_trigger_x_x1902_symbol : Boolean;
        signal ptr_deref_324_active_x_x1903_symbol : Boolean;
        signal ptr_deref_324_base_address_calculated_1904_symbol : Boolean;
        signal ptr_deref_324_root_address_calculated_1905_symbol : Boolean;
        signal ptr_deref_324_word_address_calculated_1906_symbol : Boolean;
        signal ptr_deref_324_request_1907_symbol : Boolean;
        signal ptr_deref_324_complete_1933_symbol : Boolean;
        signal assign_stmt_329_active_x_x1961_symbol : Boolean;
        signal assign_stmt_329_completed_x_x1962_symbol : Boolean;
        signal type_cast_328_active_x_x1963_symbol : Boolean;
        signal type_cast_328_trigger_x_x1964_symbol : Boolean;
        signal simple_obj_ref_327_complete_1965_symbol : Boolean;
        signal type_cast_328_complete_1966_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_325_to_assign_stmt_334_1897_start <= assign_stmt_325_to_assign_stmt_334_x_xentry_x_xx_x660_symbol; -- control passed to block
        Xentry_1898_symbol  <= assign_stmt_325_to_assign_stmt_334_1897_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/$entry
        assign_stmt_325_active_x_x1900_symbol <= ptr_deref_324_complete_1933_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_325_active_
        assign_stmt_325_completed_x_x1901_symbol <= assign_stmt_325_active_x_x1900_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_325_completed_
        ptr_deref_324_trigger_x_x1902_symbol <= ptr_deref_324_word_address_calculated_1906_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_trigger_
        ptr_deref_324_active_x_x1903_symbol <= ptr_deref_324_request_1907_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_active_
        ptr_deref_324_base_address_calculated_1904_symbol <= Xentry_1898_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_base_address_calculated
        ptr_deref_324_root_address_calculated_1905_symbol <= Xentry_1898_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_root_address_calculated
        ptr_deref_324_word_address_calculated_1906_symbol <= ptr_deref_324_root_address_calculated_1905_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_word_address_calculated
        ptr_deref_324_request_1907: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request 
          signal ptr_deref_324_request_1907_start: Boolean;
          signal Xentry_1908_symbol: Boolean;
          signal Xexit_1909_symbol: Boolean;
          signal word_access_1910_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_324_request_1907_start <= ptr_deref_324_trigger_x_x1902_symbol; -- control passed to block
          Xentry_1908_symbol  <= ptr_deref_324_request_1907_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/$entry
          word_access_1910: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access 
            signal word_access_1910_start: Boolean;
            signal Xentry_1911_symbol: Boolean;
            signal Xexit_1912_symbol: Boolean;
            signal word_access_0_1913_symbol : Boolean;
            signal word_access_1_1918_symbol : Boolean;
            signal word_access_2_1923_symbol : Boolean;
            signal word_access_3_1928_symbol : Boolean;
            -- 
          begin -- 
            word_access_1910_start <= Xentry_1908_symbol; -- control passed to block
            Xentry_1911_symbol  <= word_access_1910_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/$entry
            word_access_0_1913: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0 
              signal word_access_0_1913_start: Boolean;
              signal Xentry_1914_symbol: Boolean;
              signal Xexit_1915_symbol: Boolean;
              signal rr_1916_symbol : Boolean;
              signal ra_1917_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1913_start <= Xentry_1911_symbol; -- control passed to block
              Xentry_1914_symbol  <= word_access_0_1913_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/$entry
              rr_1916_symbol <= Xentry_1914_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/rr
              ptr_deref_324_load_0_req_0 <= rr_1916_symbol; -- link to DP
              ra_1917_symbol <= ptr_deref_324_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/ra
              Xexit_1915_symbol <= ra_1917_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/$exit
              word_access_0_1913_symbol <= Xexit_1915_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0
            word_access_1_1918: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_1 
              signal word_access_1_1918_start: Boolean;
              signal Xentry_1919_symbol: Boolean;
              signal Xexit_1920_symbol: Boolean;
              signal rr_1921_symbol : Boolean;
              signal ra_1922_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1918_start <= Xentry_1911_symbol; -- control passed to block
              Xentry_1919_symbol  <= word_access_1_1918_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_1/$entry
              rr_1921_symbol <= Xentry_1919_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_1/rr
              ptr_deref_324_load_1_req_0 <= rr_1921_symbol; -- link to DP
              ra_1922_symbol <= ptr_deref_324_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_1/ra
              Xexit_1920_symbol <= ra_1922_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_1/$exit
              word_access_1_1918_symbol <= Xexit_1920_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_1
            word_access_2_1923: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_2 
              signal word_access_2_1923_start: Boolean;
              signal Xentry_1924_symbol: Boolean;
              signal Xexit_1925_symbol: Boolean;
              signal rr_1926_symbol : Boolean;
              signal ra_1927_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1923_start <= Xentry_1911_symbol; -- control passed to block
              Xentry_1924_symbol  <= word_access_2_1923_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_2/$entry
              rr_1926_symbol <= Xentry_1924_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_2/rr
              ptr_deref_324_load_2_req_0 <= rr_1926_symbol; -- link to DP
              ra_1927_symbol <= ptr_deref_324_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_2/ra
              Xexit_1925_symbol <= ra_1927_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_2/$exit
              word_access_2_1923_symbol <= Xexit_1925_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_2
            word_access_3_1928: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_3 
              signal word_access_3_1928_start: Boolean;
              signal Xentry_1929_symbol: Boolean;
              signal Xexit_1930_symbol: Boolean;
              signal rr_1931_symbol : Boolean;
              signal ra_1932_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1928_start <= Xentry_1911_symbol; -- control passed to block
              Xentry_1929_symbol  <= word_access_3_1928_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_3/$entry
              rr_1931_symbol <= Xentry_1929_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_3/rr
              ptr_deref_324_load_3_req_0 <= rr_1931_symbol; -- link to DP
              ra_1932_symbol <= ptr_deref_324_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_3/ra
              Xexit_1930_symbol <= ra_1932_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_3/$exit
              word_access_3_1928_symbol <= Xexit_1930_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_3
            Xexit_1912_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/$exit 
              signal Xexit_1912_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1912_predecessors(0) <= word_access_0_1913_symbol;
              Xexit_1912_predecessors(1) <= word_access_1_1918_symbol;
              Xexit_1912_predecessors(2) <= word_access_2_1923_symbol;
              Xexit_1912_predecessors(3) <= word_access_3_1928_symbol;
              Xexit_1912_join: join -- 
                port map( -- 
                  preds => Xexit_1912_predecessors,
                  symbol_out => Xexit_1912_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/$exit
            word_access_1910_symbol <= Xexit_1912_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access
          Xexit_1909_symbol <= word_access_1910_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/$exit
          ptr_deref_324_request_1907_symbol <= Xexit_1909_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request
        ptr_deref_324_complete_1933: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete 
          signal ptr_deref_324_complete_1933_start: Boolean;
          signal Xentry_1934_symbol: Boolean;
          signal Xexit_1935_symbol: Boolean;
          signal word_access_1936_symbol : Boolean;
          signal merge_req_1959_symbol : Boolean;
          signal merge_ack_1960_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_324_complete_1933_start <= ptr_deref_324_active_x_x1903_symbol; -- control passed to block
          Xentry_1934_symbol  <= ptr_deref_324_complete_1933_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/$entry
          word_access_1936: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access 
            signal word_access_1936_start: Boolean;
            signal Xentry_1937_symbol: Boolean;
            signal Xexit_1938_symbol: Boolean;
            signal word_access_0_1939_symbol : Boolean;
            signal word_access_1_1944_symbol : Boolean;
            signal word_access_2_1949_symbol : Boolean;
            signal word_access_3_1954_symbol : Boolean;
            -- 
          begin -- 
            word_access_1936_start <= Xentry_1934_symbol; -- control passed to block
            Xentry_1937_symbol  <= word_access_1936_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/$entry
            word_access_0_1939: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0 
              signal word_access_0_1939_start: Boolean;
              signal Xentry_1940_symbol: Boolean;
              signal Xexit_1941_symbol: Boolean;
              signal cr_1942_symbol : Boolean;
              signal ca_1943_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1939_start <= Xentry_1937_symbol; -- control passed to block
              Xentry_1940_symbol  <= word_access_0_1939_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/$entry
              cr_1942_symbol <= Xentry_1940_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/cr
              ptr_deref_324_load_0_req_1 <= cr_1942_symbol; -- link to DP
              ca_1943_symbol <= ptr_deref_324_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/ca
              Xexit_1941_symbol <= ca_1943_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/$exit
              word_access_0_1939_symbol <= Xexit_1941_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0
            word_access_1_1944: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_1 
              signal word_access_1_1944_start: Boolean;
              signal Xentry_1945_symbol: Boolean;
              signal Xexit_1946_symbol: Boolean;
              signal cr_1947_symbol : Boolean;
              signal ca_1948_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_1944_start <= Xentry_1937_symbol; -- control passed to block
              Xentry_1945_symbol  <= word_access_1_1944_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_1/$entry
              cr_1947_symbol <= Xentry_1945_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_1/cr
              ptr_deref_324_load_1_req_1 <= cr_1947_symbol; -- link to DP
              ca_1948_symbol <= ptr_deref_324_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_1/ca
              Xexit_1946_symbol <= ca_1948_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_1/$exit
              word_access_1_1944_symbol <= Xexit_1946_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_1
            word_access_2_1949: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_2 
              signal word_access_2_1949_start: Boolean;
              signal Xentry_1950_symbol: Boolean;
              signal Xexit_1951_symbol: Boolean;
              signal cr_1952_symbol : Boolean;
              signal ca_1953_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_1949_start <= Xentry_1937_symbol; -- control passed to block
              Xentry_1950_symbol  <= word_access_2_1949_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_2/$entry
              cr_1952_symbol <= Xentry_1950_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_2/cr
              ptr_deref_324_load_2_req_1 <= cr_1952_symbol; -- link to DP
              ca_1953_symbol <= ptr_deref_324_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_2/ca
              Xexit_1951_symbol <= ca_1953_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_2/$exit
              word_access_2_1949_symbol <= Xexit_1951_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_2
            word_access_3_1954: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_3 
              signal word_access_3_1954_start: Boolean;
              signal Xentry_1955_symbol: Boolean;
              signal Xexit_1956_symbol: Boolean;
              signal cr_1957_symbol : Boolean;
              signal ca_1958_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_1954_start <= Xentry_1937_symbol; -- control passed to block
              Xentry_1955_symbol  <= word_access_3_1954_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_3/$entry
              cr_1957_symbol <= Xentry_1955_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_3/cr
              ptr_deref_324_load_3_req_1 <= cr_1957_symbol; -- link to DP
              ca_1958_symbol <= ptr_deref_324_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_3/ca
              Xexit_1956_symbol <= ca_1958_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_3/$exit
              word_access_3_1954_symbol <= Xexit_1956_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_3
            Xexit_1938_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/$exit 
              signal Xexit_1938_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_1938_predecessors(0) <= word_access_0_1939_symbol;
              Xexit_1938_predecessors(1) <= word_access_1_1944_symbol;
              Xexit_1938_predecessors(2) <= word_access_2_1949_symbol;
              Xexit_1938_predecessors(3) <= word_access_3_1954_symbol;
              Xexit_1938_join: join -- 
                port map( -- 
                  preds => Xexit_1938_predecessors,
                  symbol_out => Xexit_1938_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/$exit
            word_access_1936_symbol <= Xexit_1938_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access
          merge_req_1959_symbol <= word_access_1936_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/merge_req
          ptr_deref_324_gather_scatter_req_0 <= merge_req_1959_symbol; -- link to DP
          merge_ack_1960_symbol <= ptr_deref_324_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/merge_ack
          Xexit_1935_symbol <= merge_ack_1960_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/$exit
          ptr_deref_324_complete_1933_symbol <= Xexit_1935_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete
        assign_stmt_329_active_x_x1961_symbol <= type_cast_328_complete_1966_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_329_active_
        assign_stmt_329_completed_x_x1962_symbol <= assign_stmt_329_active_x_x1961_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_329_completed_
        type_cast_328_active_x_x1963_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_active_ 
          signal type_cast_328_active_x_x1963_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_328_active_x_x1963_predecessors(0) <= type_cast_328_trigger_x_x1964_symbol;
          type_cast_328_active_x_x1963_predecessors(1) <= simple_obj_ref_327_complete_1965_symbol;
          type_cast_328_active_x_x1963_join: join -- 
            port map( -- 
              preds => type_cast_328_active_x_x1963_predecessors,
              symbol_out => type_cast_328_active_x_x1963_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_active_
        type_cast_328_trigger_x_x1964_symbol <= Xentry_1898_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_trigger_
        simple_obj_ref_327_complete_1965_symbol <= assign_stmt_325_completed_x_x1901_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/simple_obj_ref_327_complete
        type_cast_328_complete_1966: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete 
          signal type_cast_328_complete_1966_start: Boolean;
          signal Xentry_1967_symbol: Boolean;
          signal Xexit_1968_symbol: Boolean;
          signal req_1969_symbol : Boolean;
          signal ack_1970_symbol : Boolean;
          -- 
        begin -- 
          type_cast_328_complete_1966_start <= type_cast_328_active_x_x1963_symbol; -- control passed to block
          Xentry_1967_symbol  <= type_cast_328_complete_1966_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/$entry
          req_1969_symbol <= Xentry_1967_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/req
          type_cast_328_inst_req_0 <= req_1969_symbol; -- link to DP
          ack_1970_symbol <= type_cast_328_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/ack
          Xexit_1968_symbol <= ack_1970_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/$exit
          type_cast_328_complete_1966_symbol <= Xexit_1968_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete
        Xexit_1899_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/$exit 
          signal Xexit_1899_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_1899_predecessors(0) <= ptr_deref_324_base_address_calculated_1904_symbol;
          Xexit_1899_predecessors(1) <= assign_stmt_329_completed_x_x1962_symbol;
          Xexit_1899_join: join -- 
            port map( -- 
              preds => Xexit_1899_predecessors,
              symbol_out => Xexit_1899_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/$exit
        assign_stmt_325_to_assign_stmt_334_1897_symbol <= Xexit_1899_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334
      assign_stmt_338_1971: Block -- branch_block_stmt_134/assign_stmt_338 
        signal assign_stmt_338_1971_start: Boolean;
        signal Xentry_1972_symbol: Boolean;
        signal Xexit_1973_symbol: Boolean;
        signal assign_stmt_338_active_x_x1974_symbol : Boolean;
        signal assign_stmt_338_completed_x_x1975_symbol : Boolean;
        signal type_cast_337_active_x_x1976_symbol : Boolean;
        signal type_cast_337_trigger_x_x1977_symbol : Boolean;
        signal simple_obj_ref_336_complete_1978_symbol : Boolean;
        signal type_cast_337_complete_1979_symbol : Boolean;
        signal simple_obj_ref_335_trigger_x_x1984_symbol : Boolean;
        signal simple_obj_ref_335_complete_1985_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_338_1971_start <= assign_stmt_338_x_xentry_x_xx_x662_symbol; -- control passed to block
        Xentry_1972_symbol  <= assign_stmt_338_1971_start; -- transition branch_block_stmt_134/assign_stmt_338/$entry
        assign_stmt_338_active_x_x1974_symbol <= type_cast_337_complete_1979_symbol; -- transition branch_block_stmt_134/assign_stmt_338/assign_stmt_338_active_
        assign_stmt_338_completed_x_x1975_symbol <= simple_obj_ref_335_complete_1985_symbol; -- transition branch_block_stmt_134/assign_stmt_338/assign_stmt_338_completed_
        type_cast_337_active_x_x1976_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_338/type_cast_337_active_ 
          signal type_cast_337_active_x_x1976_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_337_active_x_x1976_predecessors(0) <= type_cast_337_trigger_x_x1977_symbol;
          type_cast_337_active_x_x1976_predecessors(1) <= simple_obj_ref_336_complete_1978_symbol;
          type_cast_337_active_x_x1976_join: join -- 
            port map( -- 
              preds => type_cast_337_active_x_x1976_predecessors,
              symbol_out => type_cast_337_active_x_x1976_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_338/type_cast_337_active_
        type_cast_337_trigger_x_x1977_symbol <= Xentry_1972_symbol; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_trigger_
        simple_obj_ref_336_complete_1978_symbol <= Xentry_1972_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_336_complete
        type_cast_337_complete_1979: Block -- branch_block_stmt_134/assign_stmt_338/type_cast_337_complete 
          signal type_cast_337_complete_1979_start: Boolean;
          signal Xentry_1980_symbol: Boolean;
          signal Xexit_1981_symbol: Boolean;
          signal req_1982_symbol : Boolean;
          signal ack_1983_symbol : Boolean;
          -- 
        begin -- 
          type_cast_337_complete_1979_start <= type_cast_337_active_x_x1976_symbol; -- control passed to block
          Xentry_1980_symbol  <= type_cast_337_complete_1979_start; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/$entry
          req_1982_symbol <= Xentry_1980_symbol; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/req
          type_cast_337_inst_req_0 <= req_1982_symbol; -- link to DP
          ack_1983_symbol <= type_cast_337_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/ack
          Xexit_1981_symbol <= ack_1983_symbol; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/$exit
          type_cast_337_complete_1979_symbol <= Xexit_1981_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_338/type_cast_337_complete
        simple_obj_ref_335_trigger_x_x1984_symbol <= assign_stmt_338_active_x_x1974_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_trigger_
        simple_obj_ref_335_complete_1985: Block -- branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete 
          signal simple_obj_ref_335_complete_1985_start: Boolean;
          signal Xentry_1986_symbol: Boolean;
          signal Xexit_1987_symbol: Boolean;
          signal pipe_wreq_1988_symbol : Boolean;
          signal pipe_wack_1989_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_335_complete_1985_start <= simple_obj_ref_335_trigger_x_x1984_symbol; -- control passed to block
          Xentry_1986_symbol  <= simple_obj_ref_335_complete_1985_start; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/$entry
          pipe_wreq_1988_symbol <= Xentry_1986_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/pipe_wreq
          simple_obj_ref_335_inst_req_0 <= pipe_wreq_1988_symbol; -- link to DP
          pipe_wack_1989_symbol <= simple_obj_ref_335_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/pipe_wack
          Xexit_1987_symbol <= pipe_wack_1989_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/$exit
          simple_obj_ref_335_complete_1985_symbol <= Xexit_1987_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete
        Xexit_1973_symbol <= assign_stmt_338_completed_x_x1975_symbol; -- transition branch_block_stmt_134/assign_stmt_338/$exit
        assign_stmt_338_1971_symbol <= Xexit_1973_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_338
      assign_stmt_344_to_assign_stmt_353_1990: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353 
        signal assign_stmt_344_to_assign_stmt_353_1990_start: Boolean;
        signal Xentry_1991_symbol: Boolean;
        signal Xexit_1992_symbol: Boolean;
        signal assign_stmt_344_active_x_x1993_symbol : Boolean;
        signal assign_stmt_344_completed_x_x1994_symbol : Boolean;
        signal ptr_deref_343_trigger_x_x1995_symbol : Boolean;
        signal ptr_deref_343_active_x_x1996_symbol : Boolean;
        signal ptr_deref_343_base_address_calculated_1997_symbol : Boolean;
        signal ptr_deref_343_root_address_calculated_1998_symbol : Boolean;
        signal ptr_deref_343_word_address_calculated_1999_symbol : Boolean;
        signal ptr_deref_343_request_2000_symbol : Boolean;
        signal ptr_deref_343_complete_2011_symbol : Boolean;
        signal assign_stmt_348_active_x_x2024_symbol : Boolean;
        signal assign_stmt_348_completed_x_x2025_symbol : Boolean;
        signal type_cast_347_active_x_x2026_symbol : Boolean;
        signal type_cast_347_trigger_x_x2027_symbol : Boolean;
        signal simple_obj_ref_346_complete_2028_symbol : Boolean;
        signal type_cast_347_complete_2029_symbol : Boolean;
        signal assign_stmt_353_active_x_x2034_symbol : Boolean;
        signal assign_stmt_353_completed_x_x2035_symbol : Boolean;
        signal binary_352_active_x_x2036_symbol : Boolean;
        signal binary_352_trigger_x_x2037_symbol : Boolean;
        signal simple_obj_ref_350_complete_2038_symbol : Boolean;
        signal binary_352_complete_2039_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_344_to_assign_stmt_353_1990_start <= assign_stmt_344_to_assign_stmt_353_x_xentry_x_xx_x666_symbol; -- control passed to block
        Xentry_1991_symbol  <= assign_stmt_344_to_assign_stmt_353_1990_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/$entry
        assign_stmt_344_active_x_x1993_symbol <= ptr_deref_343_complete_2011_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_344_active_
        assign_stmt_344_completed_x_x1994_symbol <= assign_stmt_344_active_x_x1993_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_344_completed_
        ptr_deref_343_trigger_x_x1995_symbol <= ptr_deref_343_word_address_calculated_1999_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_trigger_
        ptr_deref_343_active_x_x1996_symbol <= ptr_deref_343_request_2000_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_active_
        ptr_deref_343_base_address_calculated_1997_symbol <= Xentry_1991_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_base_address_calculated
        ptr_deref_343_root_address_calculated_1998_symbol <= Xentry_1991_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_root_address_calculated
        ptr_deref_343_word_address_calculated_1999_symbol <= ptr_deref_343_root_address_calculated_1998_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_word_address_calculated
        ptr_deref_343_request_2000: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request 
          signal ptr_deref_343_request_2000_start: Boolean;
          signal Xentry_2001_symbol: Boolean;
          signal Xexit_2002_symbol: Boolean;
          signal word_access_2003_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_343_request_2000_start <= ptr_deref_343_trigger_x_x1995_symbol; -- control passed to block
          Xentry_2001_symbol  <= ptr_deref_343_request_2000_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/$entry
          word_access_2003: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access 
            signal word_access_2003_start: Boolean;
            signal Xentry_2004_symbol: Boolean;
            signal Xexit_2005_symbol: Boolean;
            signal word_access_0_2006_symbol : Boolean;
            -- 
          begin -- 
            word_access_2003_start <= Xentry_2001_symbol; -- control passed to block
            Xentry_2004_symbol  <= word_access_2003_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/$entry
            word_access_0_2006: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0 
              signal word_access_0_2006_start: Boolean;
              signal Xentry_2007_symbol: Boolean;
              signal Xexit_2008_symbol: Boolean;
              signal rr_2009_symbol : Boolean;
              signal ra_2010_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2006_start <= Xentry_2004_symbol; -- control passed to block
              Xentry_2007_symbol  <= word_access_0_2006_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/$entry
              rr_2009_symbol <= Xentry_2007_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/rr
              ptr_deref_343_load_0_req_0 <= rr_2009_symbol; -- link to DP
              ra_2010_symbol <= ptr_deref_343_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/ra
              Xexit_2008_symbol <= ra_2010_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/$exit
              word_access_0_2006_symbol <= Xexit_2008_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0
            Xexit_2005_symbol <= word_access_0_2006_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/$exit
            word_access_2003_symbol <= Xexit_2005_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access
          Xexit_2002_symbol <= word_access_2003_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/$exit
          ptr_deref_343_request_2000_symbol <= Xexit_2002_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request
        ptr_deref_343_complete_2011: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete 
          signal ptr_deref_343_complete_2011_start: Boolean;
          signal Xentry_2012_symbol: Boolean;
          signal Xexit_2013_symbol: Boolean;
          signal word_access_2014_symbol : Boolean;
          signal merge_req_2022_symbol : Boolean;
          signal merge_ack_2023_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_343_complete_2011_start <= ptr_deref_343_active_x_x1996_symbol; -- control passed to block
          Xentry_2012_symbol  <= ptr_deref_343_complete_2011_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/$entry
          word_access_2014: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access 
            signal word_access_2014_start: Boolean;
            signal Xentry_2015_symbol: Boolean;
            signal Xexit_2016_symbol: Boolean;
            signal word_access_0_2017_symbol : Boolean;
            -- 
          begin -- 
            word_access_2014_start <= Xentry_2012_symbol; -- control passed to block
            Xentry_2015_symbol  <= word_access_2014_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/$entry
            word_access_0_2017: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0 
              signal word_access_0_2017_start: Boolean;
              signal Xentry_2018_symbol: Boolean;
              signal Xexit_2019_symbol: Boolean;
              signal cr_2020_symbol : Boolean;
              signal ca_2021_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2017_start <= Xentry_2015_symbol; -- control passed to block
              Xentry_2018_symbol  <= word_access_0_2017_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/$entry
              cr_2020_symbol <= Xentry_2018_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/cr
              ptr_deref_343_load_0_req_1 <= cr_2020_symbol; -- link to DP
              ca_2021_symbol <= ptr_deref_343_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/ca
              Xexit_2019_symbol <= ca_2021_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/$exit
              word_access_0_2017_symbol <= Xexit_2019_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0
            Xexit_2016_symbol <= word_access_0_2017_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/$exit
            word_access_2014_symbol <= Xexit_2016_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access
          merge_req_2022_symbol <= word_access_2014_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/merge_req
          ptr_deref_343_gather_scatter_req_0 <= merge_req_2022_symbol; -- link to DP
          merge_ack_2023_symbol <= ptr_deref_343_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/merge_ack
          Xexit_2013_symbol <= merge_ack_2023_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/$exit
          ptr_deref_343_complete_2011_symbol <= Xexit_2013_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete
        assign_stmt_348_active_x_x2024_symbol <= type_cast_347_complete_2029_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_348_active_
        assign_stmt_348_completed_x_x2025_symbol <= assign_stmt_348_active_x_x2024_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_348_completed_
        type_cast_347_active_x_x2026_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_active_ 
          signal type_cast_347_active_x_x2026_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_347_active_x_x2026_predecessors(0) <= type_cast_347_trigger_x_x2027_symbol;
          type_cast_347_active_x_x2026_predecessors(1) <= simple_obj_ref_346_complete_2028_symbol;
          type_cast_347_active_x_x2026_join: join -- 
            port map( -- 
              preds => type_cast_347_active_x_x2026_predecessors,
              symbol_out => type_cast_347_active_x_x2026_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_active_
        type_cast_347_trigger_x_x2027_symbol <= Xentry_1991_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_trigger_
        simple_obj_ref_346_complete_2028_symbol <= assign_stmt_344_completed_x_x1994_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/simple_obj_ref_346_complete
        type_cast_347_complete_2029: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete 
          signal type_cast_347_complete_2029_start: Boolean;
          signal Xentry_2030_symbol: Boolean;
          signal Xexit_2031_symbol: Boolean;
          signal req_2032_symbol : Boolean;
          signal ack_2033_symbol : Boolean;
          -- 
        begin -- 
          type_cast_347_complete_2029_start <= type_cast_347_active_x_x2026_symbol; -- control passed to block
          Xentry_2030_symbol  <= type_cast_347_complete_2029_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/$entry
          req_2032_symbol <= Xentry_2030_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/req
          type_cast_347_inst_req_0 <= req_2032_symbol; -- link to DP
          ack_2033_symbol <= type_cast_347_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/ack
          Xexit_2031_symbol <= ack_2033_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/$exit
          type_cast_347_complete_2029_symbol <= Xexit_2031_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete
        assign_stmt_353_active_x_x2034_symbol <= binary_352_complete_2039_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_353_active_
        assign_stmt_353_completed_x_x2035_symbol <= assign_stmt_353_active_x_x2034_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_353_completed_
        binary_352_active_x_x2036_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_active_ 
          signal binary_352_active_x_x2036_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_352_active_x_x2036_predecessors(0) <= binary_352_trigger_x_x2037_symbol;
          binary_352_active_x_x2036_predecessors(1) <= simple_obj_ref_350_complete_2038_symbol;
          binary_352_active_x_x2036_join: join -- 
            port map( -- 
              preds => binary_352_active_x_x2036_predecessors,
              symbol_out => binary_352_active_x_x2036_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_active_
        binary_352_trigger_x_x2037_symbol <= Xentry_1991_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_trigger_
        simple_obj_ref_350_complete_2038_symbol <= assign_stmt_348_completed_x_x2025_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/simple_obj_ref_350_complete
        binary_352_complete_2039: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete 
          signal binary_352_complete_2039_start: Boolean;
          signal Xentry_2040_symbol: Boolean;
          signal Xexit_2041_symbol: Boolean;
          signal rr_2042_symbol : Boolean;
          signal ra_2043_symbol : Boolean;
          signal cr_2044_symbol : Boolean;
          signal ca_2045_symbol : Boolean;
          -- 
        begin -- 
          binary_352_complete_2039_start <= binary_352_active_x_x2036_symbol; -- control passed to block
          Xentry_2040_symbol  <= binary_352_complete_2039_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/$entry
          rr_2042_symbol <= Xentry_2040_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/rr
          binary_352_inst_req_0 <= rr_2042_symbol; -- link to DP
          ra_2043_symbol <= binary_352_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/ra
          cr_2044_symbol <= ra_2043_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/cr
          binary_352_inst_req_1 <= cr_2044_symbol; -- link to DP
          ca_2045_symbol <= binary_352_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/ca
          Xexit_2041_symbol <= ca_2045_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/$exit
          binary_352_complete_2039_symbol <= Xexit_2041_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete
        Xexit_1992_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/$exit 
          signal Xexit_1992_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_1992_predecessors(0) <= ptr_deref_343_base_address_calculated_1997_symbol;
          Xexit_1992_predecessors(1) <= assign_stmt_353_completed_x_x2035_symbol;
          Xexit_1992_join: join -- 
            port map( -- 
              preds => Xexit_1992_predecessors,
              symbol_out => Xexit_1992_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/$exit
        assign_stmt_344_to_assign_stmt_353_1990_symbol <= Xexit_1992_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353
      if_stmt_354_dead_link_2046: Block -- branch_block_stmt_134/if_stmt_354_dead_link 
        signal if_stmt_354_dead_link_2046_start: Boolean;
        signal Xentry_2047_symbol: Boolean;
        signal Xexit_2048_symbol: Boolean;
        signal dead_transition_2049_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_dead_link_2046_start <= if_stmt_354_x_xentry_x_xx_x668_symbol; -- control passed to block
        Xentry_2047_symbol  <= if_stmt_354_dead_link_2046_start; -- transition branch_block_stmt_134/if_stmt_354_dead_link/$entry
        dead_transition_2049_symbol <= false;
        Xexit_2048_symbol <= dead_transition_2049_symbol; -- transition branch_block_stmt_134/if_stmt_354_dead_link/$exit
        if_stmt_354_dead_link_2046_symbol <= Xexit_2048_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_dead_link
      if_stmt_354_eval_test_2050: Block -- branch_block_stmt_134/if_stmt_354_eval_test 
        signal if_stmt_354_eval_test_2050_start: Boolean;
        signal Xentry_2051_symbol: Boolean;
        signal Xexit_2052_symbol: Boolean;
        signal branch_req_2053_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_eval_test_2050_start <= if_stmt_354_x_xentry_x_xx_x668_symbol; -- control passed to block
        Xentry_2051_symbol  <= if_stmt_354_eval_test_2050_start; -- transition branch_block_stmt_134/if_stmt_354_eval_test/$entry
        branch_req_2053_symbol <= Xentry_2051_symbol; -- transition branch_block_stmt_134/if_stmt_354_eval_test/branch_req
        if_stmt_354_branch_req_0 <= branch_req_2053_symbol; -- link to DP
        Xexit_2052_symbol <= branch_req_2053_symbol; -- transition branch_block_stmt_134/if_stmt_354_eval_test/$exit
        if_stmt_354_eval_test_2050_symbol <= Xexit_2052_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_eval_test
      simple_obj_ref_355_place_2054_symbol  <=  if_stmt_354_eval_test_2050_symbol; -- place branch_block_stmt_134/simple_obj_ref_355_place (optimized away) 
      if_stmt_354_if_link_2055: Block -- branch_block_stmt_134/if_stmt_354_if_link 
        signal if_stmt_354_if_link_2055_start: Boolean;
        signal Xentry_2056_symbol: Boolean;
        signal Xexit_2057_symbol: Boolean;
        signal if_choice_transition_2058_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_if_link_2055_start <= simple_obj_ref_355_place_2054_symbol; -- control passed to block
        Xentry_2056_symbol  <= if_stmt_354_if_link_2055_start; -- transition branch_block_stmt_134/if_stmt_354_if_link/$entry
        if_choice_transition_2058_symbol <= if_stmt_354_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_354_if_link/if_choice_transition
        Xexit_2057_symbol <= if_choice_transition_2058_symbol; -- transition branch_block_stmt_134/if_stmt_354_if_link/$exit
        if_stmt_354_if_link_2055_symbol <= Xexit_2057_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_if_link
      if_stmt_354_else_link_2059: Block -- branch_block_stmt_134/if_stmt_354_else_link 
        signal if_stmt_354_else_link_2059_start: Boolean;
        signal Xentry_2060_symbol: Boolean;
        signal Xexit_2061_symbol: Boolean;
        signal else_choice_transition_2062_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_else_link_2059_start <= simple_obj_ref_355_place_2054_symbol; -- control passed to block
        Xentry_2060_symbol  <= if_stmt_354_else_link_2059_start; -- transition branch_block_stmt_134/if_stmt_354_else_link/$entry
        else_choice_transition_2062_symbol <= if_stmt_354_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_354_else_link/else_choice_transition
        Xexit_2061_symbol <= else_choice_transition_2062_symbol; -- transition branch_block_stmt_134/if_stmt_354_else_link/$exit
        if_stmt_354_else_link_2059_symbol <= Xexit_2061_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_else_link
      bb_8_bb_9_2063_symbol  <=  if_stmt_354_if_link_2055_symbol; -- place branch_block_stmt_134/bb_8_bb_9 (optimized away) 
      bb_8_bb_4_2064_symbol  <=  if_stmt_354_else_link_2059_symbol; -- place branch_block_stmt_134/bb_8_bb_4 (optimized away) 
      assign_stmt_365_2065: Block -- branch_block_stmt_134/assign_stmt_365 
        signal assign_stmt_365_2065_start: Boolean;
        signal Xentry_2066_symbol: Boolean;
        signal Xexit_2067_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_365_2065_start <= assign_stmt_365_x_xentry_x_xx_x672_symbol; -- control passed to block
        Xentry_2066_symbol  <= assign_stmt_365_2065_start; -- transition branch_block_stmt_134/assign_stmt_365/$entry
        Xexit_2067_symbol <= Xentry_2066_symbol; -- transition branch_block_stmt_134/assign_stmt_365/$exit
        assign_stmt_365_2065_symbol <= Xexit_2067_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_365
      assign_stmt_369_2068: Block -- branch_block_stmt_134/assign_stmt_369 
        signal assign_stmt_369_2068_start: Boolean;
        signal Xentry_2069_symbol: Boolean;
        signal Xexit_2070_symbol: Boolean;
        signal assign_stmt_369_active_x_x2071_symbol : Boolean;
        signal assign_stmt_369_completed_x_x2072_symbol : Boolean;
        signal type_cast_368_active_x_x2073_symbol : Boolean;
        signal type_cast_368_trigger_x_x2074_symbol : Boolean;
        signal simple_obj_ref_367_trigger_x_x2075_symbol : Boolean;
        signal simple_obj_ref_367_complete_2076_symbol : Boolean;
        signal type_cast_368_complete_2081_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_369_2068_start <= assign_stmt_369_x_xentry_x_xx_x674_symbol; -- control passed to block
        Xentry_2069_symbol  <= assign_stmt_369_2068_start; -- transition branch_block_stmt_134/assign_stmt_369/$entry
        assign_stmt_369_active_x_x2071_symbol <= type_cast_368_complete_2081_symbol; -- transition branch_block_stmt_134/assign_stmt_369/assign_stmt_369_active_
        assign_stmt_369_completed_x_x2072_symbol <= assign_stmt_369_active_x_x2071_symbol; -- transition branch_block_stmt_134/assign_stmt_369/assign_stmt_369_completed_
        type_cast_368_active_x_x2073_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_369/type_cast_368_active_ 
          signal type_cast_368_active_x_x2073_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_368_active_x_x2073_predecessors(0) <= type_cast_368_trigger_x_x2074_symbol;
          type_cast_368_active_x_x2073_predecessors(1) <= simple_obj_ref_367_complete_2076_symbol;
          type_cast_368_active_x_x2073_join: join -- 
            port map( -- 
              preds => type_cast_368_active_x_x2073_predecessors,
              symbol_out => type_cast_368_active_x_x2073_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_369/type_cast_368_active_
        type_cast_368_trigger_x_x2074_symbol <= Xentry_2069_symbol; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_trigger_
        simple_obj_ref_367_trigger_x_x2075_symbol <= Xentry_2069_symbol; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_trigger_
        simple_obj_ref_367_complete_2076: Block -- branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete 
          signal simple_obj_ref_367_complete_2076_start: Boolean;
          signal Xentry_2077_symbol: Boolean;
          signal Xexit_2078_symbol: Boolean;
          signal req_2079_symbol : Boolean;
          signal ack_2080_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_367_complete_2076_start <= simple_obj_ref_367_trigger_x_x2075_symbol; -- control passed to block
          Xentry_2077_symbol  <= simple_obj_ref_367_complete_2076_start; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/$entry
          req_2079_symbol <= Xentry_2077_symbol; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/req
          simple_obj_ref_367_inst_req_0 <= req_2079_symbol; -- link to DP
          ack_2080_symbol <= simple_obj_ref_367_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/ack
          Xexit_2078_symbol <= ack_2080_symbol; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/$exit
          simple_obj_ref_367_complete_2076_symbol <= Xexit_2078_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete
        type_cast_368_complete_2081: Block -- branch_block_stmt_134/assign_stmt_369/type_cast_368_complete 
          signal type_cast_368_complete_2081_start: Boolean;
          signal Xentry_2082_symbol: Boolean;
          signal Xexit_2083_symbol: Boolean;
          signal req_2084_symbol : Boolean;
          signal ack_2085_symbol : Boolean;
          -- 
        begin -- 
          type_cast_368_complete_2081_start <= type_cast_368_active_x_x2073_symbol; -- control passed to block
          Xentry_2082_symbol  <= type_cast_368_complete_2081_start; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/$entry
          req_2084_symbol <= Xentry_2082_symbol; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/req
          type_cast_368_inst_req_0 <= req_2084_symbol; -- link to DP
          ack_2085_symbol <= type_cast_368_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/ack
          Xexit_2083_symbol <= ack_2085_symbol; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/$exit
          type_cast_368_complete_2081_symbol <= Xexit_2083_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_369/type_cast_368_complete
        Xexit_2070_symbol <= assign_stmt_369_completed_x_x2072_symbol; -- transition branch_block_stmt_134/assign_stmt_369/$exit
        assign_stmt_369_2068_symbol <= Xexit_2070_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_369
      assign_stmt_373_to_assign_stmt_400_2086: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400 
        signal assign_stmt_373_to_assign_stmt_400_2086_start: Boolean;
        signal Xentry_2087_symbol: Boolean;
        signal Xexit_2088_symbol: Boolean;
        signal assign_stmt_373_active_x_x2089_symbol : Boolean;
        signal assign_stmt_373_completed_x_x2090_symbol : Boolean;
        signal type_cast_372_active_x_x2091_symbol : Boolean;
        signal type_cast_372_trigger_x_x2092_symbol : Boolean;
        signal simple_obj_ref_371_complete_2093_symbol : Boolean;
        signal type_cast_372_complete_2094_symbol : Boolean;
        signal assign_stmt_377_active_x_x2099_symbol : Boolean;
        signal assign_stmt_377_completed_x_x2100_symbol : Boolean;
        signal simple_obj_ref_376_complete_2101_symbol : Boolean;
        signal ptr_deref_375_trigger_x_x2102_symbol : Boolean;
        signal ptr_deref_375_active_x_x2103_symbol : Boolean;
        signal ptr_deref_375_base_address_calculated_2104_symbol : Boolean;
        signal ptr_deref_375_root_address_calculated_2105_symbol : Boolean;
        signal ptr_deref_375_word_address_calculated_2106_symbol : Boolean;
        signal ptr_deref_375_request_2107_symbol : Boolean;
        signal ptr_deref_375_complete_2135_symbol : Boolean;
        signal assign_stmt_380_active_x_x2161_symbol : Boolean;
        signal assign_stmt_380_completed_x_x2162_symbol : Boolean;
        signal simple_obj_ref_379_trigger_x_x2163_symbol : Boolean;
        signal simple_obj_ref_379_active_x_x2164_symbol : Boolean;
        signal simple_obj_ref_379_root_address_calculated_2165_symbol : Boolean;
        signal simple_obj_ref_379_word_address_calculated_2166_symbol : Boolean;
        signal simple_obj_ref_379_request_2167_symbol : Boolean;
        signal simple_obj_ref_379_complete_2178_symbol : Boolean;
        signal assign_stmt_384_active_x_x2191_symbol : Boolean;
        signal assign_stmt_384_completed_x_x2192_symbol : Boolean;
        signal ptr_deref_383_trigger_x_x2193_symbol : Boolean;
        signal ptr_deref_383_active_x_x2194_symbol : Boolean;
        signal ptr_deref_383_base_address_calculated_2195_symbol : Boolean;
        signal ptr_deref_383_root_address_calculated_2196_symbol : Boolean;
        signal ptr_deref_383_word_address_calculated_2197_symbol : Boolean;
        signal ptr_deref_383_request_2198_symbol : Boolean;
        signal ptr_deref_383_complete_2224_symbol : Boolean;
        signal assign_stmt_389_active_x_x2252_symbol : Boolean;
        signal assign_stmt_389_completed_x_x2253_symbol : Boolean;
        signal array_obj_ref_388_trigger_x_x2254_symbol : Boolean;
        signal array_obj_ref_388_active_x_x2255_symbol : Boolean;
        signal array_obj_ref_388_base_address_calculated_2256_symbol : Boolean;
        signal array_obj_ref_388_root_address_calculated_2257_symbol : Boolean;
        signal array_obj_ref_388_base_address_resized_2258_symbol : Boolean;
        signal array_obj_ref_388_base_addr_resize_2259_symbol : Boolean;
        signal array_obj_ref_388_base_plus_offset_2264_symbol : Boolean;
        signal array_obj_ref_388_complete_2269_symbol : Boolean;
        signal assign_stmt_393_active_x_x2274_symbol : Boolean;
        signal assign_stmt_393_completed_x_x2275_symbol : Boolean;
        signal simple_obj_ref_392_complete_2276_symbol : Boolean;
        signal ptr_deref_391_trigger_x_x2277_symbol : Boolean;
        signal ptr_deref_391_active_x_x2278_symbol : Boolean;
        signal ptr_deref_391_base_address_calculated_2279_symbol : Boolean;
        signal simple_obj_ref_390_complete_2280_symbol : Boolean;
        signal ptr_deref_391_root_address_calculated_2281_symbol : Boolean;
        signal ptr_deref_391_word_address_calculated_2282_symbol : Boolean;
        signal ptr_deref_391_base_address_resized_2283_symbol : Boolean;
        signal ptr_deref_391_base_addr_resize_2284_symbol : Boolean;
        signal ptr_deref_391_base_plus_offset_2289_symbol : Boolean;
        signal ptr_deref_391_word_addrgen_2294_symbol : Boolean;
        signal ptr_deref_391_request_2325_symbol : Boolean;
        signal ptr_deref_391_complete_2353_symbol : Boolean;
        signal assign_stmt_397_active_x_x2379_symbol : Boolean;
        signal assign_stmt_397_completed_x_x2380_symbol : Boolean;
        signal ptr_deref_396_trigger_x_x2381_symbol : Boolean;
        signal ptr_deref_396_active_x_x2382_symbol : Boolean;
        signal ptr_deref_396_base_address_calculated_2383_symbol : Boolean;
        signal ptr_deref_396_root_address_calculated_2384_symbol : Boolean;
        signal ptr_deref_396_word_address_calculated_2385_symbol : Boolean;
        signal ptr_deref_396_request_2386_symbol : Boolean;
        signal ptr_deref_396_complete_2412_symbol : Boolean;
        signal assign_stmt_400_active_x_x2440_symbol : Boolean;
        signal assign_stmt_400_completed_x_x2441_symbol : Boolean;
        signal simple_obj_ref_399_complete_2442_symbol : Boolean;
        signal simple_obj_ref_398_trigger_x_x2443_symbol : Boolean;
        signal simple_obj_ref_398_active_x_x2444_symbol : Boolean;
        signal simple_obj_ref_398_root_address_calculated_2445_symbol : Boolean;
        signal simple_obj_ref_398_word_address_calculated_2446_symbol : Boolean;
        signal simple_obj_ref_398_request_2447_symbol : Boolean;
        signal simple_obj_ref_398_complete_2460_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_373_to_assign_stmt_400_2086_start <= assign_stmt_373_to_assign_stmt_400_x_xentry_x_xx_x676_symbol; -- control passed to block
        Xentry_2087_symbol  <= assign_stmt_373_to_assign_stmt_400_2086_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/$entry
        assign_stmt_373_active_x_x2089_symbol <= type_cast_372_complete_2094_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_373_active_
        assign_stmt_373_completed_x_x2090_symbol <= assign_stmt_373_active_x_x2089_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_373_completed_
        type_cast_372_active_x_x2091_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_active_ 
          signal type_cast_372_active_x_x2091_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_372_active_x_x2091_predecessors(0) <= type_cast_372_trigger_x_x2092_symbol;
          type_cast_372_active_x_x2091_predecessors(1) <= simple_obj_ref_371_complete_2093_symbol;
          type_cast_372_active_x_x2091_join: join -- 
            port map( -- 
              preds => type_cast_372_active_x_x2091_predecessors,
              symbol_out => type_cast_372_active_x_x2091_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_active_
        type_cast_372_trigger_x_x2092_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_trigger_
        simple_obj_ref_371_complete_2093_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_371_complete
        type_cast_372_complete_2094: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete 
          signal type_cast_372_complete_2094_start: Boolean;
          signal Xentry_2095_symbol: Boolean;
          signal Xexit_2096_symbol: Boolean;
          signal req_2097_symbol : Boolean;
          signal ack_2098_symbol : Boolean;
          -- 
        begin -- 
          type_cast_372_complete_2094_start <= type_cast_372_active_x_x2091_symbol; -- control passed to block
          Xentry_2095_symbol  <= type_cast_372_complete_2094_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/$entry
          req_2097_symbol <= Xentry_2095_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/req
          type_cast_372_inst_req_0 <= req_2097_symbol; -- link to DP
          ack_2098_symbol <= type_cast_372_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/ack
          Xexit_2096_symbol <= ack_2098_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/$exit
          type_cast_372_complete_2094_symbol <= Xexit_2096_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete
        assign_stmt_377_active_x_x2099_symbol <= simple_obj_ref_376_complete_2101_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_377_active_
        assign_stmt_377_completed_x_x2100_symbol <= ptr_deref_375_complete_2135_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_377_completed_
        simple_obj_ref_376_complete_2101_symbol <= assign_stmt_373_completed_x_x2090_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_376_complete
        ptr_deref_375_trigger_x_x2102_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_trigger_ 
          signal ptr_deref_375_trigger_x_x2102_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_375_trigger_x_x2102_predecessors(0) <= ptr_deref_375_word_address_calculated_2106_symbol;
          ptr_deref_375_trigger_x_x2102_predecessors(1) <= assign_stmt_377_active_x_x2099_symbol;
          ptr_deref_375_trigger_x_x2102_join: join -- 
            port map( -- 
              preds => ptr_deref_375_trigger_x_x2102_predecessors,
              symbol_out => ptr_deref_375_trigger_x_x2102_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_trigger_
        ptr_deref_375_active_x_x2103_symbol <= ptr_deref_375_request_2107_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_active_
        ptr_deref_375_base_address_calculated_2104_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_base_address_calculated
        ptr_deref_375_root_address_calculated_2105_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_root_address_calculated
        ptr_deref_375_word_address_calculated_2106_symbol <= ptr_deref_375_root_address_calculated_2105_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_word_address_calculated
        ptr_deref_375_request_2107: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request 
          signal ptr_deref_375_request_2107_start: Boolean;
          signal Xentry_2108_symbol: Boolean;
          signal Xexit_2109_symbol: Boolean;
          signal split_req_2110_symbol : Boolean;
          signal split_ack_2111_symbol : Boolean;
          signal word_access_2112_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_375_request_2107_start <= ptr_deref_375_trigger_x_x2102_symbol; -- control passed to block
          Xentry_2108_symbol  <= ptr_deref_375_request_2107_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/$entry
          split_req_2110_symbol <= Xentry_2108_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/split_req
          ptr_deref_375_gather_scatter_req_0 <= split_req_2110_symbol; -- link to DP
          split_ack_2111_symbol <= ptr_deref_375_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/split_ack
          word_access_2112: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access 
            signal word_access_2112_start: Boolean;
            signal Xentry_2113_symbol: Boolean;
            signal Xexit_2114_symbol: Boolean;
            signal word_access_0_2115_symbol : Boolean;
            signal word_access_1_2120_symbol : Boolean;
            signal word_access_2_2125_symbol : Boolean;
            signal word_access_3_2130_symbol : Boolean;
            -- 
          begin -- 
            word_access_2112_start <= split_ack_2111_symbol; -- control passed to block
            Xentry_2113_symbol  <= word_access_2112_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/$entry
            word_access_0_2115: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0 
              signal word_access_0_2115_start: Boolean;
              signal Xentry_2116_symbol: Boolean;
              signal Xexit_2117_symbol: Boolean;
              signal rr_2118_symbol : Boolean;
              signal ra_2119_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2115_start <= Xentry_2113_symbol; -- control passed to block
              Xentry_2116_symbol  <= word_access_0_2115_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/$entry
              rr_2118_symbol <= Xentry_2116_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/rr
              ptr_deref_375_store_0_req_0 <= rr_2118_symbol; -- link to DP
              ra_2119_symbol <= ptr_deref_375_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/ra
              Xexit_2117_symbol <= ra_2119_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/$exit
              word_access_0_2115_symbol <= Xexit_2117_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0
            word_access_1_2120: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_1 
              signal word_access_1_2120_start: Boolean;
              signal Xentry_2121_symbol: Boolean;
              signal Xexit_2122_symbol: Boolean;
              signal rr_2123_symbol : Boolean;
              signal ra_2124_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2120_start <= Xentry_2113_symbol; -- control passed to block
              Xentry_2121_symbol  <= word_access_1_2120_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_1/$entry
              rr_2123_symbol <= Xentry_2121_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_1/rr
              ptr_deref_375_store_1_req_0 <= rr_2123_symbol; -- link to DP
              ra_2124_symbol <= ptr_deref_375_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_1/ra
              Xexit_2122_symbol <= ra_2124_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_1/$exit
              word_access_1_2120_symbol <= Xexit_2122_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_1
            word_access_2_2125: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_2 
              signal word_access_2_2125_start: Boolean;
              signal Xentry_2126_symbol: Boolean;
              signal Xexit_2127_symbol: Boolean;
              signal rr_2128_symbol : Boolean;
              signal ra_2129_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2125_start <= Xentry_2113_symbol; -- control passed to block
              Xentry_2126_symbol  <= word_access_2_2125_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_2/$entry
              rr_2128_symbol <= Xentry_2126_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_2/rr
              ptr_deref_375_store_2_req_0 <= rr_2128_symbol; -- link to DP
              ra_2129_symbol <= ptr_deref_375_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_2/ra
              Xexit_2127_symbol <= ra_2129_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_2/$exit
              word_access_2_2125_symbol <= Xexit_2127_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_2
            word_access_3_2130: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_3 
              signal word_access_3_2130_start: Boolean;
              signal Xentry_2131_symbol: Boolean;
              signal Xexit_2132_symbol: Boolean;
              signal rr_2133_symbol : Boolean;
              signal ra_2134_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2130_start <= Xentry_2113_symbol; -- control passed to block
              Xentry_2131_symbol  <= word_access_3_2130_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_3/$entry
              rr_2133_symbol <= Xentry_2131_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_3/rr
              ptr_deref_375_store_3_req_0 <= rr_2133_symbol; -- link to DP
              ra_2134_symbol <= ptr_deref_375_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_3/ra
              Xexit_2132_symbol <= ra_2134_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_3/$exit
              word_access_3_2130_symbol <= Xexit_2132_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_3
            Xexit_2114_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/$exit 
              signal Xexit_2114_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2114_predecessors(0) <= word_access_0_2115_symbol;
              Xexit_2114_predecessors(1) <= word_access_1_2120_symbol;
              Xexit_2114_predecessors(2) <= word_access_2_2125_symbol;
              Xexit_2114_predecessors(3) <= word_access_3_2130_symbol;
              Xexit_2114_join: join -- 
                port map( -- 
                  preds => Xexit_2114_predecessors,
                  symbol_out => Xexit_2114_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/$exit
            word_access_2112_symbol <= Xexit_2114_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access
          Xexit_2109_symbol <= word_access_2112_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/$exit
          ptr_deref_375_request_2107_symbol <= Xexit_2109_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request
        ptr_deref_375_complete_2135: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete 
          signal ptr_deref_375_complete_2135_start: Boolean;
          signal Xentry_2136_symbol: Boolean;
          signal Xexit_2137_symbol: Boolean;
          signal word_access_2138_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_375_complete_2135_start <= ptr_deref_375_active_x_x2103_symbol; -- control passed to block
          Xentry_2136_symbol  <= ptr_deref_375_complete_2135_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/$entry
          word_access_2138: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access 
            signal word_access_2138_start: Boolean;
            signal Xentry_2139_symbol: Boolean;
            signal Xexit_2140_symbol: Boolean;
            signal word_access_0_2141_symbol : Boolean;
            signal word_access_1_2146_symbol : Boolean;
            signal word_access_2_2151_symbol : Boolean;
            signal word_access_3_2156_symbol : Boolean;
            -- 
          begin -- 
            word_access_2138_start <= Xentry_2136_symbol; -- control passed to block
            Xentry_2139_symbol  <= word_access_2138_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/$entry
            word_access_0_2141: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0 
              signal word_access_0_2141_start: Boolean;
              signal Xentry_2142_symbol: Boolean;
              signal Xexit_2143_symbol: Boolean;
              signal cr_2144_symbol : Boolean;
              signal ca_2145_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2141_start <= Xentry_2139_symbol; -- control passed to block
              Xentry_2142_symbol  <= word_access_0_2141_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/$entry
              cr_2144_symbol <= Xentry_2142_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/cr
              ptr_deref_375_store_0_req_1 <= cr_2144_symbol; -- link to DP
              ca_2145_symbol <= ptr_deref_375_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/ca
              Xexit_2143_symbol <= ca_2145_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/$exit
              word_access_0_2141_symbol <= Xexit_2143_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0
            word_access_1_2146: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_1 
              signal word_access_1_2146_start: Boolean;
              signal Xentry_2147_symbol: Boolean;
              signal Xexit_2148_symbol: Boolean;
              signal cr_2149_symbol : Boolean;
              signal ca_2150_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2146_start <= Xentry_2139_symbol; -- control passed to block
              Xentry_2147_symbol  <= word_access_1_2146_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_1/$entry
              cr_2149_symbol <= Xentry_2147_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_1/cr
              ptr_deref_375_store_1_req_1 <= cr_2149_symbol; -- link to DP
              ca_2150_symbol <= ptr_deref_375_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_1/ca
              Xexit_2148_symbol <= ca_2150_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_1/$exit
              word_access_1_2146_symbol <= Xexit_2148_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_1
            word_access_2_2151: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_2 
              signal word_access_2_2151_start: Boolean;
              signal Xentry_2152_symbol: Boolean;
              signal Xexit_2153_symbol: Boolean;
              signal cr_2154_symbol : Boolean;
              signal ca_2155_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2151_start <= Xentry_2139_symbol; -- control passed to block
              Xentry_2152_symbol  <= word_access_2_2151_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_2/$entry
              cr_2154_symbol <= Xentry_2152_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_2/cr
              ptr_deref_375_store_2_req_1 <= cr_2154_symbol; -- link to DP
              ca_2155_symbol <= ptr_deref_375_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_2/ca
              Xexit_2153_symbol <= ca_2155_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_2/$exit
              word_access_2_2151_symbol <= Xexit_2153_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_2
            word_access_3_2156: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_3 
              signal word_access_3_2156_start: Boolean;
              signal Xentry_2157_symbol: Boolean;
              signal Xexit_2158_symbol: Boolean;
              signal cr_2159_symbol : Boolean;
              signal ca_2160_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2156_start <= Xentry_2139_symbol; -- control passed to block
              Xentry_2157_symbol  <= word_access_3_2156_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_3/$entry
              cr_2159_symbol <= Xentry_2157_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_3/cr
              ptr_deref_375_store_3_req_1 <= cr_2159_symbol; -- link to DP
              ca_2160_symbol <= ptr_deref_375_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_3/ca
              Xexit_2158_symbol <= ca_2160_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_3/$exit
              word_access_3_2156_symbol <= Xexit_2158_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_3
            Xexit_2140_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/$exit 
              signal Xexit_2140_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2140_predecessors(0) <= word_access_0_2141_symbol;
              Xexit_2140_predecessors(1) <= word_access_1_2146_symbol;
              Xexit_2140_predecessors(2) <= word_access_2_2151_symbol;
              Xexit_2140_predecessors(3) <= word_access_3_2156_symbol;
              Xexit_2140_join: join -- 
                port map( -- 
                  preds => Xexit_2140_predecessors,
                  symbol_out => Xexit_2140_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/$exit
            word_access_2138_symbol <= Xexit_2140_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access
          Xexit_2137_symbol <= word_access_2138_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/$exit
          ptr_deref_375_complete_2135_symbol <= Xexit_2137_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete
        assign_stmt_380_active_x_x2161_symbol <= simple_obj_ref_379_complete_2178_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_380_active_
        assign_stmt_380_completed_x_x2162_symbol <= assign_stmt_380_active_x_x2161_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_380_completed_
        simple_obj_ref_379_trigger_x_x2163_symbol <= simple_obj_ref_379_word_address_calculated_2166_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_trigger_
        simple_obj_ref_379_active_x_x2164_symbol <= simple_obj_ref_379_request_2167_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_active_
        simple_obj_ref_379_root_address_calculated_2165_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_root_address_calculated
        simple_obj_ref_379_word_address_calculated_2166_symbol <= simple_obj_ref_379_root_address_calculated_2165_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_word_address_calculated
        simple_obj_ref_379_request_2167: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request 
          signal simple_obj_ref_379_request_2167_start: Boolean;
          signal Xentry_2168_symbol: Boolean;
          signal Xexit_2169_symbol: Boolean;
          signal word_access_2170_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_379_request_2167_start <= simple_obj_ref_379_trigger_x_x2163_symbol; -- control passed to block
          Xentry_2168_symbol  <= simple_obj_ref_379_request_2167_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/$entry
          word_access_2170: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access 
            signal word_access_2170_start: Boolean;
            signal Xentry_2171_symbol: Boolean;
            signal Xexit_2172_symbol: Boolean;
            signal word_access_0_2173_symbol : Boolean;
            -- 
          begin -- 
            word_access_2170_start <= Xentry_2168_symbol; -- control passed to block
            Xentry_2171_symbol  <= word_access_2170_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/$entry
            word_access_0_2173: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0 
              signal word_access_0_2173_start: Boolean;
              signal Xentry_2174_symbol: Boolean;
              signal Xexit_2175_symbol: Boolean;
              signal rr_2176_symbol : Boolean;
              signal ra_2177_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2173_start <= Xentry_2171_symbol; -- control passed to block
              Xentry_2174_symbol  <= word_access_0_2173_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/$entry
              rr_2176_symbol <= Xentry_2174_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/rr
              simple_obj_ref_379_load_0_req_0 <= rr_2176_symbol; -- link to DP
              ra_2177_symbol <= simple_obj_ref_379_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/ra
              Xexit_2175_symbol <= ra_2177_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/$exit
              word_access_0_2173_symbol <= Xexit_2175_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0
            Xexit_2172_symbol <= word_access_0_2173_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/$exit
            word_access_2170_symbol <= Xexit_2172_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access
          Xexit_2169_symbol <= word_access_2170_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/$exit
          simple_obj_ref_379_request_2167_symbol <= Xexit_2169_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request
        simple_obj_ref_379_complete_2178: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete 
          signal simple_obj_ref_379_complete_2178_start: Boolean;
          signal Xentry_2179_symbol: Boolean;
          signal Xexit_2180_symbol: Boolean;
          signal word_access_2181_symbol : Boolean;
          signal merge_req_2189_symbol : Boolean;
          signal merge_ack_2190_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_379_complete_2178_start <= simple_obj_ref_379_active_x_x2164_symbol; -- control passed to block
          Xentry_2179_symbol  <= simple_obj_ref_379_complete_2178_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/$entry
          word_access_2181: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access 
            signal word_access_2181_start: Boolean;
            signal Xentry_2182_symbol: Boolean;
            signal Xexit_2183_symbol: Boolean;
            signal word_access_0_2184_symbol : Boolean;
            -- 
          begin -- 
            word_access_2181_start <= Xentry_2179_symbol; -- control passed to block
            Xentry_2182_symbol  <= word_access_2181_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/$entry
            word_access_0_2184: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0 
              signal word_access_0_2184_start: Boolean;
              signal Xentry_2185_symbol: Boolean;
              signal Xexit_2186_symbol: Boolean;
              signal cr_2187_symbol : Boolean;
              signal ca_2188_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2184_start <= Xentry_2182_symbol; -- control passed to block
              Xentry_2185_symbol  <= word_access_0_2184_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/$entry
              cr_2187_symbol <= Xentry_2185_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/cr
              simple_obj_ref_379_load_0_req_1 <= cr_2187_symbol; -- link to DP
              ca_2188_symbol <= simple_obj_ref_379_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/ca
              Xexit_2186_symbol <= ca_2188_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/$exit
              word_access_0_2184_symbol <= Xexit_2186_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0
            Xexit_2183_symbol <= word_access_0_2184_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/$exit
            word_access_2181_symbol <= Xexit_2183_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access
          merge_req_2189_symbol <= word_access_2181_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/merge_req
          simple_obj_ref_379_gather_scatter_req_0 <= merge_req_2189_symbol; -- link to DP
          merge_ack_2190_symbol <= simple_obj_ref_379_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/merge_ack
          Xexit_2180_symbol <= merge_ack_2190_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/$exit
          simple_obj_ref_379_complete_2178_symbol <= Xexit_2180_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete
        assign_stmt_384_active_x_x2191_symbol <= ptr_deref_383_complete_2224_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_384_active_
        assign_stmt_384_completed_x_x2192_symbol <= assign_stmt_384_active_x_x2191_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_384_completed_
        ptr_deref_383_trigger_x_x2193_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_trigger_ 
          signal ptr_deref_383_trigger_x_x2193_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_383_trigger_x_x2193_predecessors(0) <= ptr_deref_383_word_address_calculated_2197_symbol;
          ptr_deref_383_trigger_x_x2193_predecessors(1) <= ptr_deref_375_active_x_x2103_symbol;
          ptr_deref_383_trigger_x_x2193_join: join -- 
            port map( -- 
              preds => ptr_deref_383_trigger_x_x2193_predecessors,
              symbol_out => ptr_deref_383_trigger_x_x2193_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_trigger_
        ptr_deref_383_active_x_x2194_symbol <= ptr_deref_383_request_2198_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_active_
        ptr_deref_383_base_address_calculated_2195_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_base_address_calculated
        ptr_deref_383_root_address_calculated_2196_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_root_address_calculated
        ptr_deref_383_word_address_calculated_2197_symbol <= ptr_deref_383_root_address_calculated_2196_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_word_address_calculated
        ptr_deref_383_request_2198: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request 
          signal ptr_deref_383_request_2198_start: Boolean;
          signal Xentry_2199_symbol: Boolean;
          signal Xexit_2200_symbol: Boolean;
          signal word_access_2201_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_383_request_2198_start <= ptr_deref_383_trigger_x_x2193_symbol; -- control passed to block
          Xentry_2199_symbol  <= ptr_deref_383_request_2198_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/$entry
          word_access_2201: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access 
            signal word_access_2201_start: Boolean;
            signal Xentry_2202_symbol: Boolean;
            signal Xexit_2203_symbol: Boolean;
            signal word_access_0_2204_symbol : Boolean;
            signal word_access_1_2209_symbol : Boolean;
            signal word_access_2_2214_symbol : Boolean;
            signal word_access_3_2219_symbol : Boolean;
            -- 
          begin -- 
            word_access_2201_start <= Xentry_2199_symbol; -- control passed to block
            Xentry_2202_symbol  <= word_access_2201_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/$entry
            word_access_0_2204: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0 
              signal word_access_0_2204_start: Boolean;
              signal Xentry_2205_symbol: Boolean;
              signal Xexit_2206_symbol: Boolean;
              signal rr_2207_symbol : Boolean;
              signal ra_2208_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2204_start <= Xentry_2202_symbol; -- control passed to block
              Xentry_2205_symbol  <= word_access_0_2204_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/$entry
              rr_2207_symbol <= Xentry_2205_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/rr
              ptr_deref_383_load_0_req_0 <= rr_2207_symbol; -- link to DP
              ra_2208_symbol <= ptr_deref_383_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/ra
              Xexit_2206_symbol <= ra_2208_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/$exit
              word_access_0_2204_symbol <= Xexit_2206_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0
            word_access_1_2209: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_1 
              signal word_access_1_2209_start: Boolean;
              signal Xentry_2210_symbol: Boolean;
              signal Xexit_2211_symbol: Boolean;
              signal rr_2212_symbol : Boolean;
              signal ra_2213_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2209_start <= Xentry_2202_symbol; -- control passed to block
              Xentry_2210_symbol  <= word_access_1_2209_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_1/$entry
              rr_2212_symbol <= Xentry_2210_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_1/rr
              ptr_deref_383_load_1_req_0 <= rr_2212_symbol; -- link to DP
              ra_2213_symbol <= ptr_deref_383_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_1/ra
              Xexit_2211_symbol <= ra_2213_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_1/$exit
              word_access_1_2209_symbol <= Xexit_2211_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_1
            word_access_2_2214: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_2 
              signal word_access_2_2214_start: Boolean;
              signal Xentry_2215_symbol: Boolean;
              signal Xexit_2216_symbol: Boolean;
              signal rr_2217_symbol : Boolean;
              signal ra_2218_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2214_start <= Xentry_2202_symbol; -- control passed to block
              Xentry_2215_symbol  <= word_access_2_2214_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_2/$entry
              rr_2217_symbol <= Xentry_2215_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_2/rr
              ptr_deref_383_load_2_req_0 <= rr_2217_symbol; -- link to DP
              ra_2218_symbol <= ptr_deref_383_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_2/ra
              Xexit_2216_symbol <= ra_2218_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_2/$exit
              word_access_2_2214_symbol <= Xexit_2216_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_2
            word_access_3_2219: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_3 
              signal word_access_3_2219_start: Boolean;
              signal Xentry_2220_symbol: Boolean;
              signal Xexit_2221_symbol: Boolean;
              signal rr_2222_symbol : Boolean;
              signal ra_2223_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2219_start <= Xentry_2202_symbol; -- control passed to block
              Xentry_2220_symbol  <= word_access_3_2219_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_3/$entry
              rr_2222_symbol <= Xentry_2220_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_3/rr
              ptr_deref_383_load_3_req_0 <= rr_2222_symbol; -- link to DP
              ra_2223_symbol <= ptr_deref_383_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_3/ra
              Xexit_2221_symbol <= ra_2223_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_3/$exit
              word_access_3_2219_symbol <= Xexit_2221_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_3
            Xexit_2203_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/$exit 
              signal Xexit_2203_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2203_predecessors(0) <= word_access_0_2204_symbol;
              Xexit_2203_predecessors(1) <= word_access_1_2209_symbol;
              Xexit_2203_predecessors(2) <= word_access_2_2214_symbol;
              Xexit_2203_predecessors(3) <= word_access_3_2219_symbol;
              Xexit_2203_join: join -- 
                port map( -- 
                  preds => Xexit_2203_predecessors,
                  symbol_out => Xexit_2203_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/$exit
            word_access_2201_symbol <= Xexit_2203_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access
          Xexit_2200_symbol <= word_access_2201_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/$exit
          ptr_deref_383_request_2198_symbol <= Xexit_2200_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request
        ptr_deref_383_complete_2224: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete 
          signal ptr_deref_383_complete_2224_start: Boolean;
          signal Xentry_2225_symbol: Boolean;
          signal Xexit_2226_symbol: Boolean;
          signal word_access_2227_symbol : Boolean;
          signal merge_req_2250_symbol : Boolean;
          signal merge_ack_2251_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_383_complete_2224_start <= ptr_deref_383_active_x_x2194_symbol; -- control passed to block
          Xentry_2225_symbol  <= ptr_deref_383_complete_2224_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/$entry
          word_access_2227: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access 
            signal word_access_2227_start: Boolean;
            signal Xentry_2228_symbol: Boolean;
            signal Xexit_2229_symbol: Boolean;
            signal word_access_0_2230_symbol : Boolean;
            signal word_access_1_2235_symbol : Boolean;
            signal word_access_2_2240_symbol : Boolean;
            signal word_access_3_2245_symbol : Boolean;
            -- 
          begin -- 
            word_access_2227_start <= Xentry_2225_symbol; -- control passed to block
            Xentry_2228_symbol  <= word_access_2227_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/$entry
            word_access_0_2230: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0 
              signal word_access_0_2230_start: Boolean;
              signal Xentry_2231_symbol: Boolean;
              signal Xexit_2232_symbol: Boolean;
              signal cr_2233_symbol : Boolean;
              signal ca_2234_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2230_start <= Xentry_2228_symbol; -- control passed to block
              Xentry_2231_symbol  <= word_access_0_2230_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/$entry
              cr_2233_symbol <= Xentry_2231_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/cr
              ptr_deref_383_load_0_req_1 <= cr_2233_symbol; -- link to DP
              ca_2234_symbol <= ptr_deref_383_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/ca
              Xexit_2232_symbol <= ca_2234_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/$exit
              word_access_0_2230_symbol <= Xexit_2232_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0
            word_access_1_2235: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_1 
              signal word_access_1_2235_start: Boolean;
              signal Xentry_2236_symbol: Boolean;
              signal Xexit_2237_symbol: Boolean;
              signal cr_2238_symbol : Boolean;
              signal ca_2239_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2235_start <= Xentry_2228_symbol; -- control passed to block
              Xentry_2236_symbol  <= word_access_1_2235_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_1/$entry
              cr_2238_symbol <= Xentry_2236_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_1/cr
              ptr_deref_383_load_1_req_1 <= cr_2238_symbol; -- link to DP
              ca_2239_symbol <= ptr_deref_383_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_1/ca
              Xexit_2237_symbol <= ca_2239_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_1/$exit
              word_access_1_2235_symbol <= Xexit_2237_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_1
            word_access_2_2240: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_2 
              signal word_access_2_2240_start: Boolean;
              signal Xentry_2241_symbol: Boolean;
              signal Xexit_2242_symbol: Boolean;
              signal cr_2243_symbol : Boolean;
              signal ca_2244_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2240_start <= Xentry_2228_symbol; -- control passed to block
              Xentry_2241_symbol  <= word_access_2_2240_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_2/$entry
              cr_2243_symbol <= Xentry_2241_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_2/cr
              ptr_deref_383_load_2_req_1 <= cr_2243_symbol; -- link to DP
              ca_2244_symbol <= ptr_deref_383_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_2/ca
              Xexit_2242_symbol <= ca_2244_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_2/$exit
              word_access_2_2240_symbol <= Xexit_2242_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_2
            word_access_3_2245: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_3 
              signal word_access_3_2245_start: Boolean;
              signal Xentry_2246_symbol: Boolean;
              signal Xexit_2247_symbol: Boolean;
              signal cr_2248_symbol : Boolean;
              signal ca_2249_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2245_start <= Xentry_2228_symbol; -- control passed to block
              Xentry_2246_symbol  <= word_access_3_2245_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_3/$entry
              cr_2248_symbol <= Xentry_2246_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_3/cr
              ptr_deref_383_load_3_req_1 <= cr_2248_symbol; -- link to DP
              ca_2249_symbol <= ptr_deref_383_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_3/ca
              Xexit_2247_symbol <= ca_2249_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_3/$exit
              word_access_3_2245_symbol <= Xexit_2247_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_3
            Xexit_2229_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/$exit 
              signal Xexit_2229_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2229_predecessors(0) <= word_access_0_2230_symbol;
              Xexit_2229_predecessors(1) <= word_access_1_2235_symbol;
              Xexit_2229_predecessors(2) <= word_access_2_2240_symbol;
              Xexit_2229_predecessors(3) <= word_access_3_2245_symbol;
              Xexit_2229_join: join -- 
                port map( -- 
                  preds => Xexit_2229_predecessors,
                  symbol_out => Xexit_2229_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/$exit
            word_access_2227_symbol <= Xexit_2229_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access
          merge_req_2250_symbol <= word_access_2227_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/merge_req
          ptr_deref_383_gather_scatter_req_0 <= merge_req_2250_symbol; -- link to DP
          merge_ack_2251_symbol <= ptr_deref_383_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/merge_ack
          Xexit_2226_symbol <= merge_ack_2251_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/$exit
          ptr_deref_383_complete_2224_symbol <= Xexit_2226_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete
        assign_stmt_389_active_x_x2252_symbol <= array_obj_ref_388_complete_2269_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_389_active_
        assign_stmt_389_completed_x_x2253_symbol <= assign_stmt_389_active_x_x2252_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_389_completed_
        array_obj_ref_388_trigger_x_x2254_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_trigger_
        array_obj_ref_388_active_x_x2255_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_active_ 
          signal array_obj_ref_388_active_x_x2255_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_388_active_x_x2255_predecessors(0) <= array_obj_ref_388_trigger_x_x2254_symbol;
          array_obj_ref_388_active_x_x2255_predecessors(1) <= array_obj_ref_388_root_address_calculated_2257_symbol;
          array_obj_ref_388_active_x_x2255_join: join -- 
            port map( -- 
              preds => array_obj_ref_388_active_x_x2255_predecessors,
              symbol_out => array_obj_ref_388_active_x_x2255_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_active_
        array_obj_ref_388_base_address_calculated_2256_symbol <= assign_stmt_384_completed_x_x2192_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_address_calculated
        array_obj_ref_388_root_address_calculated_2257_symbol <= array_obj_ref_388_base_plus_offset_2264_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_root_address_calculated
        array_obj_ref_388_base_address_resized_2258_symbol <= array_obj_ref_388_base_addr_resize_2259_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_address_resized
        array_obj_ref_388_base_addr_resize_2259: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize 
          signal array_obj_ref_388_base_addr_resize_2259_start: Boolean;
          signal Xentry_2260_symbol: Boolean;
          signal Xexit_2261_symbol: Boolean;
          signal base_resize_req_2262_symbol : Boolean;
          signal base_resize_ack_2263_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_388_base_addr_resize_2259_start <= array_obj_ref_388_base_address_calculated_2256_symbol; -- control passed to block
          Xentry_2260_symbol  <= array_obj_ref_388_base_addr_resize_2259_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/$entry
          base_resize_req_2262_symbol <= Xentry_2260_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/base_resize_req
          array_obj_ref_388_base_resize_req_0 <= base_resize_req_2262_symbol; -- link to DP
          base_resize_ack_2263_symbol <= array_obj_ref_388_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/base_resize_ack
          Xexit_2261_symbol <= base_resize_ack_2263_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/$exit
          array_obj_ref_388_base_addr_resize_2259_symbol <= Xexit_2261_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize
        array_obj_ref_388_base_plus_offset_2264: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset 
          signal array_obj_ref_388_base_plus_offset_2264_start: Boolean;
          signal Xentry_2265_symbol: Boolean;
          signal Xexit_2266_symbol: Boolean;
          signal sum_rename_req_2267_symbol : Boolean;
          signal sum_rename_ack_2268_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_388_base_plus_offset_2264_start <= array_obj_ref_388_base_address_resized_2258_symbol; -- control passed to block
          Xentry_2265_symbol  <= array_obj_ref_388_base_plus_offset_2264_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/$entry
          sum_rename_req_2267_symbol <= Xentry_2265_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/sum_rename_req
          array_obj_ref_388_root_address_inst_req_0 <= sum_rename_req_2267_symbol; -- link to DP
          sum_rename_ack_2268_symbol <= array_obj_ref_388_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/sum_rename_ack
          Xexit_2266_symbol <= sum_rename_ack_2268_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/$exit
          array_obj_ref_388_base_plus_offset_2264_symbol <= Xexit_2266_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset
        array_obj_ref_388_complete_2269: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete 
          signal array_obj_ref_388_complete_2269_start: Boolean;
          signal Xentry_2270_symbol: Boolean;
          signal Xexit_2271_symbol: Boolean;
          signal final_reg_req_2272_symbol : Boolean;
          signal final_reg_ack_2273_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_388_complete_2269_start <= array_obj_ref_388_active_x_x2255_symbol; -- control passed to block
          Xentry_2270_symbol  <= array_obj_ref_388_complete_2269_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/$entry
          final_reg_req_2272_symbol <= Xentry_2270_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/final_reg_req
          array_obj_ref_388_final_reg_req_0 <= final_reg_req_2272_symbol; -- link to DP
          final_reg_ack_2273_symbol <= array_obj_ref_388_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/final_reg_ack
          Xexit_2271_symbol <= final_reg_ack_2273_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/$exit
          array_obj_ref_388_complete_2269_symbol <= Xexit_2271_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete
        assign_stmt_393_active_x_x2274_symbol <= simple_obj_ref_392_complete_2276_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_393_active_
        assign_stmt_393_completed_x_x2275_symbol <= ptr_deref_391_complete_2353_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_393_completed_
        simple_obj_ref_392_complete_2276_symbol <= assign_stmt_380_completed_x_x2162_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_392_complete
        ptr_deref_391_trigger_x_x2277_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_trigger_ 
          signal ptr_deref_391_trigger_x_x2277_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          ptr_deref_391_trigger_x_x2277_predecessors(0) <= ptr_deref_391_word_address_calculated_2282_symbol;
          ptr_deref_391_trigger_x_x2277_predecessors(1) <= ptr_deref_391_base_address_calculated_2279_symbol;
          ptr_deref_391_trigger_x_x2277_predecessors(2) <= assign_stmt_393_active_x_x2274_symbol;
          ptr_deref_391_trigger_x_x2277_predecessors(3) <= ptr_deref_383_active_x_x2194_symbol;
          ptr_deref_391_trigger_x_x2277_join: join -- 
            port map( -- 
              preds => ptr_deref_391_trigger_x_x2277_predecessors,
              symbol_out => ptr_deref_391_trigger_x_x2277_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_trigger_
        ptr_deref_391_active_x_x2278_symbol <= ptr_deref_391_request_2325_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_active_
        ptr_deref_391_base_address_calculated_2279_symbol <= simple_obj_ref_390_complete_2280_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_address_calculated
        simple_obj_ref_390_complete_2280_symbol <= assign_stmt_389_completed_x_x2253_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_390_complete
        ptr_deref_391_root_address_calculated_2281_symbol <= ptr_deref_391_base_plus_offset_2289_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_root_address_calculated
        ptr_deref_391_word_address_calculated_2282_symbol <= ptr_deref_391_word_addrgen_2294_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_address_calculated
        ptr_deref_391_base_address_resized_2283_symbol <= ptr_deref_391_base_addr_resize_2284_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_address_resized
        ptr_deref_391_base_addr_resize_2284: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize 
          signal ptr_deref_391_base_addr_resize_2284_start: Boolean;
          signal Xentry_2285_symbol: Boolean;
          signal Xexit_2286_symbol: Boolean;
          signal base_resize_req_2287_symbol : Boolean;
          signal base_resize_ack_2288_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_base_addr_resize_2284_start <= ptr_deref_391_base_address_calculated_2279_symbol; -- control passed to block
          Xentry_2285_symbol  <= ptr_deref_391_base_addr_resize_2284_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/$entry
          base_resize_req_2287_symbol <= Xentry_2285_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/base_resize_req
          ptr_deref_391_base_resize_req_0 <= base_resize_req_2287_symbol; -- link to DP
          base_resize_ack_2288_symbol <= ptr_deref_391_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/base_resize_ack
          Xexit_2286_symbol <= base_resize_ack_2288_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/$exit
          ptr_deref_391_base_addr_resize_2284_symbol <= Xexit_2286_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize
        ptr_deref_391_base_plus_offset_2289: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset 
          signal ptr_deref_391_base_plus_offset_2289_start: Boolean;
          signal Xentry_2290_symbol: Boolean;
          signal Xexit_2291_symbol: Boolean;
          signal sum_rename_req_2292_symbol : Boolean;
          signal sum_rename_ack_2293_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_base_plus_offset_2289_start <= ptr_deref_391_base_address_resized_2283_symbol; -- control passed to block
          Xentry_2290_symbol  <= ptr_deref_391_base_plus_offset_2289_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/$entry
          sum_rename_req_2292_symbol <= Xentry_2290_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/sum_rename_req
          ptr_deref_391_root_address_inst_req_0 <= sum_rename_req_2292_symbol; -- link to DP
          sum_rename_ack_2293_symbol <= ptr_deref_391_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/sum_rename_ack
          Xexit_2291_symbol <= sum_rename_ack_2293_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/$exit
          ptr_deref_391_base_plus_offset_2289_symbol <= Xexit_2291_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset
        ptr_deref_391_word_addrgen_2294: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen 
          signal ptr_deref_391_word_addrgen_2294_start: Boolean;
          signal Xentry_2295_symbol: Boolean;
          signal Xexit_2296_symbol: Boolean;
          signal word_0_2297_symbol : Boolean;
          signal word_1_2304_symbol : Boolean;
          signal word_2_2311_symbol : Boolean;
          signal word_3_2318_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_word_addrgen_2294_start <= ptr_deref_391_root_address_calculated_2281_symbol; -- control passed to block
          Xentry_2295_symbol  <= ptr_deref_391_word_addrgen_2294_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/$entry
          word_0_2297: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0 
            signal word_0_2297_start: Boolean;
            signal Xentry_2298_symbol: Boolean;
            signal Xexit_2299_symbol: Boolean;
            signal rr_2300_symbol : Boolean;
            signal ra_2301_symbol : Boolean;
            signal cr_2302_symbol : Boolean;
            signal ca_2303_symbol : Boolean;
            -- 
          begin -- 
            word_0_2297_start <= Xentry_2295_symbol; -- control passed to block
            Xentry_2298_symbol  <= word_0_2297_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0/$entry
            rr_2300_symbol <= Xentry_2298_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0/rr
            ptr_deref_391_addr_0_req_0 <= rr_2300_symbol; -- link to DP
            ra_2301_symbol <= ptr_deref_391_addr_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0/ra
            cr_2302_symbol <= ra_2301_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0/cr
            ptr_deref_391_addr_0_req_1 <= cr_2302_symbol; -- link to DP
            ca_2303_symbol <= ptr_deref_391_addr_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0/ca
            Xexit_2299_symbol <= ca_2303_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0/$exit
            word_0_2297_symbol <= Xexit_2299_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_0
          word_1_2304: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1 
            signal word_1_2304_start: Boolean;
            signal Xentry_2305_symbol: Boolean;
            signal Xexit_2306_symbol: Boolean;
            signal rr_2307_symbol : Boolean;
            signal ra_2308_symbol : Boolean;
            signal cr_2309_symbol : Boolean;
            signal ca_2310_symbol : Boolean;
            -- 
          begin -- 
            word_1_2304_start <= Xentry_2295_symbol; -- control passed to block
            Xentry_2305_symbol  <= word_1_2304_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1/$entry
            rr_2307_symbol <= Xentry_2305_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1/rr
            ptr_deref_391_addr_1_req_0 <= rr_2307_symbol; -- link to DP
            ra_2308_symbol <= ptr_deref_391_addr_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1/ra
            cr_2309_symbol <= ra_2308_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1/cr
            ptr_deref_391_addr_1_req_1 <= cr_2309_symbol; -- link to DP
            ca_2310_symbol <= ptr_deref_391_addr_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1/ca
            Xexit_2306_symbol <= ca_2310_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1/$exit
            word_1_2304_symbol <= Xexit_2306_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_1
          word_2_2311: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2 
            signal word_2_2311_start: Boolean;
            signal Xentry_2312_symbol: Boolean;
            signal Xexit_2313_symbol: Boolean;
            signal rr_2314_symbol : Boolean;
            signal ra_2315_symbol : Boolean;
            signal cr_2316_symbol : Boolean;
            signal ca_2317_symbol : Boolean;
            -- 
          begin -- 
            word_2_2311_start <= Xentry_2295_symbol; -- control passed to block
            Xentry_2312_symbol  <= word_2_2311_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2/$entry
            rr_2314_symbol <= Xentry_2312_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2/rr
            ptr_deref_391_addr_2_req_0 <= rr_2314_symbol; -- link to DP
            ra_2315_symbol <= ptr_deref_391_addr_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2/ra
            cr_2316_symbol <= ra_2315_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2/cr
            ptr_deref_391_addr_2_req_1 <= cr_2316_symbol; -- link to DP
            ca_2317_symbol <= ptr_deref_391_addr_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2/ca
            Xexit_2313_symbol <= ca_2317_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2/$exit
            word_2_2311_symbol <= Xexit_2313_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_2
          word_3_2318: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3 
            signal word_3_2318_start: Boolean;
            signal Xentry_2319_symbol: Boolean;
            signal Xexit_2320_symbol: Boolean;
            signal rr_2321_symbol : Boolean;
            signal ra_2322_symbol : Boolean;
            signal cr_2323_symbol : Boolean;
            signal ca_2324_symbol : Boolean;
            -- 
          begin -- 
            word_3_2318_start <= Xentry_2295_symbol; -- control passed to block
            Xentry_2319_symbol  <= word_3_2318_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3/$entry
            rr_2321_symbol <= Xentry_2319_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3/rr
            ptr_deref_391_addr_3_req_0 <= rr_2321_symbol; -- link to DP
            ra_2322_symbol <= ptr_deref_391_addr_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3/ra
            cr_2323_symbol <= ra_2322_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3/cr
            ptr_deref_391_addr_3_req_1 <= cr_2323_symbol; -- link to DP
            ca_2324_symbol <= ptr_deref_391_addr_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3/ca
            Xexit_2320_symbol <= ca_2324_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3/$exit
            word_3_2318_symbol <= Xexit_2320_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/word_3
          Xexit_2296_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/$exit 
            signal Xexit_2296_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_2296_predecessors(0) <= word_0_2297_symbol;
            Xexit_2296_predecessors(1) <= word_1_2304_symbol;
            Xexit_2296_predecessors(2) <= word_2_2311_symbol;
            Xexit_2296_predecessors(3) <= word_3_2318_symbol;
            Xexit_2296_join: join -- 
              port map( -- 
                preds => Xexit_2296_predecessors,
                symbol_out => Xexit_2296_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/$exit
          ptr_deref_391_word_addrgen_2294_symbol <= Xexit_2296_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen
        ptr_deref_391_request_2325: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request 
          signal ptr_deref_391_request_2325_start: Boolean;
          signal Xentry_2326_symbol: Boolean;
          signal Xexit_2327_symbol: Boolean;
          signal split_req_2328_symbol : Boolean;
          signal split_ack_2329_symbol : Boolean;
          signal word_access_2330_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_request_2325_start <= ptr_deref_391_trigger_x_x2277_symbol; -- control passed to block
          Xentry_2326_symbol  <= ptr_deref_391_request_2325_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/$entry
          split_req_2328_symbol <= Xentry_2326_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/split_req
          ptr_deref_391_gather_scatter_req_0 <= split_req_2328_symbol; -- link to DP
          split_ack_2329_symbol <= ptr_deref_391_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/split_ack
          word_access_2330: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access 
            signal word_access_2330_start: Boolean;
            signal Xentry_2331_symbol: Boolean;
            signal Xexit_2332_symbol: Boolean;
            signal word_access_0_2333_symbol : Boolean;
            signal word_access_1_2338_symbol : Boolean;
            signal word_access_2_2343_symbol : Boolean;
            signal word_access_3_2348_symbol : Boolean;
            -- 
          begin -- 
            word_access_2330_start <= split_ack_2329_symbol; -- control passed to block
            Xentry_2331_symbol  <= word_access_2330_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/$entry
            word_access_0_2333: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0 
              signal word_access_0_2333_start: Boolean;
              signal Xentry_2334_symbol: Boolean;
              signal Xexit_2335_symbol: Boolean;
              signal rr_2336_symbol : Boolean;
              signal ra_2337_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2333_start <= Xentry_2331_symbol; -- control passed to block
              Xentry_2334_symbol  <= word_access_0_2333_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/$entry
              rr_2336_symbol <= Xentry_2334_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/rr
              ptr_deref_391_store_0_req_0 <= rr_2336_symbol; -- link to DP
              ra_2337_symbol <= ptr_deref_391_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/ra
              Xexit_2335_symbol <= ra_2337_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/$exit
              word_access_0_2333_symbol <= Xexit_2335_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0
            word_access_1_2338: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_1 
              signal word_access_1_2338_start: Boolean;
              signal Xentry_2339_symbol: Boolean;
              signal Xexit_2340_symbol: Boolean;
              signal rr_2341_symbol : Boolean;
              signal ra_2342_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2338_start <= Xentry_2331_symbol; -- control passed to block
              Xentry_2339_symbol  <= word_access_1_2338_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_1/$entry
              rr_2341_symbol <= Xentry_2339_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_1/rr
              ptr_deref_391_store_1_req_0 <= rr_2341_symbol; -- link to DP
              ra_2342_symbol <= ptr_deref_391_store_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_1/ra
              Xexit_2340_symbol <= ra_2342_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_1/$exit
              word_access_1_2338_symbol <= Xexit_2340_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_1
            word_access_2_2343: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_2 
              signal word_access_2_2343_start: Boolean;
              signal Xentry_2344_symbol: Boolean;
              signal Xexit_2345_symbol: Boolean;
              signal rr_2346_symbol : Boolean;
              signal ra_2347_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2343_start <= Xentry_2331_symbol; -- control passed to block
              Xentry_2344_symbol  <= word_access_2_2343_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_2/$entry
              rr_2346_symbol <= Xentry_2344_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_2/rr
              ptr_deref_391_store_2_req_0 <= rr_2346_symbol; -- link to DP
              ra_2347_symbol <= ptr_deref_391_store_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_2/ra
              Xexit_2345_symbol <= ra_2347_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_2/$exit
              word_access_2_2343_symbol <= Xexit_2345_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_2
            word_access_3_2348: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_3 
              signal word_access_3_2348_start: Boolean;
              signal Xentry_2349_symbol: Boolean;
              signal Xexit_2350_symbol: Boolean;
              signal rr_2351_symbol : Boolean;
              signal ra_2352_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2348_start <= Xentry_2331_symbol; -- control passed to block
              Xentry_2349_symbol  <= word_access_3_2348_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_3/$entry
              rr_2351_symbol <= Xentry_2349_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_3/rr
              ptr_deref_391_store_3_req_0 <= rr_2351_symbol; -- link to DP
              ra_2352_symbol <= ptr_deref_391_store_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_3/ra
              Xexit_2350_symbol <= ra_2352_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_3/$exit
              word_access_3_2348_symbol <= Xexit_2350_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_3
            Xexit_2332_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/$exit 
              signal Xexit_2332_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2332_predecessors(0) <= word_access_0_2333_symbol;
              Xexit_2332_predecessors(1) <= word_access_1_2338_symbol;
              Xexit_2332_predecessors(2) <= word_access_2_2343_symbol;
              Xexit_2332_predecessors(3) <= word_access_3_2348_symbol;
              Xexit_2332_join: join -- 
                port map( -- 
                  preds => Xexit_2332_predecessors,
                  symbol_out => Xexit_2332_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/$exit
            word_access_2330_symbol <= Xexit_2332_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access
          Xexit_2327_symbol <= word_access_2330_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/$exit
          ptr_deref_391_request_2325_symbol <= Xexit_2327_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request
        ptr_deref_391_complete_2353: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete 
          signal ptr_deref_391_complete_2353_start: Boolean;
          signal Xentry_2354_symbol: Boolean;
          signal Xexit_2355_symbol: Boolean;
          signal word_access_2356_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_complete_2353_start <= ptr_deref_391_active_x_x2278_symbol; -- control passed to block
          Xentry_2354_symbol  <= ptr_deref_391_complete_2353_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/$entry
          word_access_2356: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access 
            signal word_access_2356_start: Boolean;
            signal Xentry_2357_symbol: Boolean;
            signal Xexit_2358_symbol: Boolean;
            signal word_access_0_2359_symbol : Boolean;
            signal word_access_1_2364_symbol : Boolean;
            signal word_access_2_2369_symbol : Boolean;
            signal word_access_3_2374_symbol : Boolean;
            -- 
          begin -- 
            word_access_2356_start <= Xentry_2354_symbol; -- control passed to block
            Xentry_2357_symbol  <= word_access_2356_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/$entry
            word_access_0_2359: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0 
              signal word_access_0_2359_start: Boolean;
              signal Xentry_2360_symbol: Boolean;
              signal Xexit_2361_symbol: Boolean;
              signal cr_2362_symbol : Boolean;
              signal ca_2363_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2359_start <= Xentry_2357_symbol; -- control passed to block
              Xentry_2360_symbol  <= word_access_0_2359_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/$entry
              cr_2362_symbol <= Xentry_2360_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/cr
              ptr_deref_391_store_0_req_1 <= cr_2362_symbol; -- link to DP
              ca_2363_symbol <= ptr_deref_391_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/ca
              Xexit_2361_symbol <= ca_2363_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/$exit
              word_access_0_2359_symbol <= Xexit_2361_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0
            word_access_1_2364: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_1 
              signal word_access_1_2364_start: Boolean;
              signal Xentry_2365_symbol: Boolean;
              signal Xexit_2366_symbol: Boolean;
              signal cr_2367_symbol : Boolean;
              signal ca_2368_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2364_start <= Xentry_2357_symbol; -- control passed to block
              Xentry_2365_symbol  <= word_access_1_2364_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_1/$entry
              cr_2367_symbol <= Xentry_2365_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_1/cr
              ptr_deref_391_store_1_req_1 <= cr_2367_symbol; -- link to DP
              ca_2368_symbol <= ptr_deref_391_store_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_1/ca
              Xexit_2366_symbol <= ca_2368_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_1/$exit
              word_access_1_2364_symbol <= Xexit_2366_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_1
            word_access_2_2369: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_2 
              signal word_access_2_2369_start: Boolean;
              signal Xentry_2370_symbol: Boolean;
              signal Xexit_2371_symbol: Boolean;
              signal cr_2372_symbol : Boolean;
              signal ca_2373_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2369_start <= Xentry_2357_symbol; -- control passed to block
              Xentry_2370_symbol  <= word_access_2_2369_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_2/$entry
              cr_2372_symbol <= Xentry_2370_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_2/cr
              ptr_deref_391_store_2_req_1 <= cr_2372_symbol; -- link to DP
              ca_2373_symbol <= ptr_deref_391_store_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_2/ca
              Xexit_2371_symbol <= ca_2373_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_2/$exit
              word_access_2_2369_symbol <= Xexit_2371_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_2
            word_access_3_2374: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_3 
              signal word_access_3_2374_start: Boolean;
              signal Xentry_2375_symbol: Boolean;
              signal Xexit_2376_symbol: Boolean;
              signal cr_2377_symbol : Boolean;
              signal ca_2378_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2374_start <= Xentry_2357_symbol; -- control passed to block
              Xentry_2375_symbol  <= word_access_3_2374_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_3/$entry
              cr_2377_symbol <= Xentry_2375_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_3/cr
              ptr_deref_391_store_3_req_1 <= cr_2377_symbol; -- link to DP
              ca_2378_symbol <= ptr_deref_391_store_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_3/ca
              Xexit_2376_symbol <= ca_2378_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_3/$exit
              word_access_3_2374_symbol <= Xexit_2376_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_3
            Xexit_2358_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/$exit 
              signal Xexit_2358_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2358_predecessors(0) <= word_access_0_2359_symbol;
              Xexit_2358_predecessors(1) <= word_access_1_2364_symbol;
              Xexit_2358_predecessors(2) <= word_access_2_2369_symbol;
              Xexit_2358_predecessors(3) <= word_access_3_2374_symbol;
              Xexit_2358_join: join -- 
                port map( -- 
                  preds => Xexit_2358_predecessors,
                  symbol_out => Xexit_2358_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/$exit
            word_access_2356_symbol <= Xexit_2358_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access
          Xexit_2355_symbol <= word_access_2356_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/$exit
          ptr_deref_391_complete_2353_symbol <= Xexit_2355_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete
        assign_stmt_397_active_x_x2379_symbol <= ptr_deref_396_complete_2412_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_397_active_
        assign_stmt_397_completed_x_x2380_symbol <= assign_stmt_397_active_x_x2379_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_397_completed_
        ptr_deref_396_trigger_x_x2381_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_trigger_ 
          signal ptr_deref_396_trigger_x_x2381_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_396_trigger_x_x2381_predecessors(0) <= ptr_deref_396_word_address_calculated_2385_symbol;
          ptr_deref_396_trigger_x_x2381_predecessors(1) <= ptr_deref_391_active_x_x2278_symbol;
          ptr_deref_396_trigger_x_x2381_join: join -- 
            port map( -- 
              preds => ptr_deref_396_trigger_x_x2381_predecessors,
              symbol_out => ptr_deref_396_trigger_x_x2381_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_trigger_
        ptr_deref_396_active_x_x2382_symbol <= ptr_deref_396_request_2386_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_active_
        ptr_deref_396_base_address_calculated_2383_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_base_address_calculated
        ptr_deref_396_root_address_calculated_2384_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_root_address_calculated
        ptr_deref_396_word_address_calculated_2385_symbol <= ptr_deref_396_root_address_calculated_2384_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_word_address_calculated
        ptr_deref_396_request_2386: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request 
          signal ptr_deref_396_request_2386_start: Boolean;
          signal Xentry_2387_symbol: Boolean;
          signal Xexit_2388_symbol: Boolean;
          signal word_access_2389_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_396_request_2386_start <= ptr_deref_396_trigger_x_x2381_symbol; -- control passed to block
          Xentry_2387_symbol  <= ptr_deref_396_request_2386_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/$entry
          word_access_2389: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access 
            signal word_access_2389_start: Boolean;
            signal Xentry_2390_symbol: Boolean;
            signal Xexit_2391_symbol: Boolean;
            signal word_access_0_2392_symbol : Boolean;
            signal word_access_1_2397_symbol : Boolean;
            signal word_access_2_2402_symbol : Boolean;
            signal word_access_3_2407_symbol : Boolean;
            -- 
          begin -- 
            word_access_2389_start <= Xentry_2387_symbol; -- control passed to block
            Xentry_2390_symbol  <= word_access_2389_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/$entry
            word_access_0_2392: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0 
              signal word_access_0_2392_start: Boolean;
              signal Xentry_2393_symbol: Boolean;
              signal Xexit_2394_symbol: Boolean;
              signal rr_2395_symbol : Boolean;
              signal ra_2396_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2392_start <= Xentry_2390_symbol; -- control passed to block
              Xentry_2393_symbol  <= word_access_0_2392_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/$entry
              rr_2395_symbol <= Xentry_2393_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/rr
              ptr_deref_396_load_0_req_0 <= rr_2395_symbol; -- link to DP
              ra_2396_symbol <= ptr_deref_396_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/ra
              Xexit_2394_symbol <= ra_2396_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/$exit
              word_access_0_2392_symbol <= Xexit_2394_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0
            word_access_1_2397: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_1 
              signal word_access_1_2397_start: Boolean;
              signal Xentry_2398_symbol: Boolean;
              signal Xexit_2399_symbol: Boolean;
              signal rr_2400_symbol : Boolean;
              signal ra_2401_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2397_start <= Xentry_2390_symbol; -- control passed to block
              Xentry_2398_symbol  <= word_access_1_2397_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_1/$entry
              rr_2400_symbol <= Xentry_2398_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_1/rr
              ptr_deref_396_load_1_req_0 <= rr_2400_symbol; -- link to DP
              ra_2401_symbol <= ptr_deref_396_load_1_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_1/ra
              Xexit_2399_symbol <= ra_2401_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_1/$exit
              word_access_1_2397_symbol <= Xexit_2399_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_1
            word_access_2_2402: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_2 
              signal word_access_2_2402_start: Boolean;
              signal Xentry_2403_symbol: Boolean;
              signal Xexit_2404_symbol: Boolean;
              signal rr_2405_symbol : Boolean;
              signal ra_2406_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2402_start <= Xentry_2390_symbol; -- control passed to block
              Xentry_2403_symbol  <= word_access_2_2402_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_2/$entry
              rr_2405_symbol <= Xentry_2403_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_2/rr
              ptr_deref_396_load_2_req_0 <= rr_2405_symbol; -- link to DP
              ra_2406_symbol <= ptr_deref_396_load_2_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_2/ra
              Xexit_2404_symbol <= ra_2406_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_2/$exit
              word_access_2_2402_symbol <= Xexit_2404_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_2
            word_access_3_2407: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_3 
              signal word_access_3_2407_start: Boolean;
              signal Xentry_2408_symbol: Boolean;
              signal Xexit_2409_symbol: Boolean;
              signal rr_2410_symbol : Boolean;
              signal ra_2411_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2407_start <= Xentry_2390_symbol; -- control passed to block
              Xentry_2408_symbol  <= word_access_3_2407_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_3/$entry
              rr_2410_symbol <= Xentry_2408_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_3/rr
              ptr_deref_396_load_3_req_0 <= rr_2410_symbol; -- link to DP
              ra_2411_symbol <= ptr_deref_396_load_3_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_3/ra
              Xexit_2409_symbol <= ra_2411_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_3/$exit
              word_access_3_2407_symbol <= Xexit_2409_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_3
            Xexit_2391_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/$exit 
              signal Xexit_2391_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2391_predecessors(0) <= word_access_0_2392_symbol;
              Xexit_2391_predecessors(1) <= word_access_1_2397_symbol;
              Xexit_2391_predecessors(2) <= word_access_2_2402_symbol;
              Xexit_2391_predecessors(3) <= word_access_3_2407_symbol;
              Xexit_2391_join: join -- 
                port map( -- 
                  preds => Xexit_2391_predecessors,
                  symbol_out => Xexit_2391_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/$exit
            word_access_2389_symbol <= Xexit_2391_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access
          Xexit_2388_symbol <= word_access_2389_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/$exit
          ptr_deref_396_request_2386_symbol <= Xexit_2388_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request
        ptr_deref_396_complete_2412: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete 
          signal ptr_deref_396_complete_2412_start: Boolean;
          signal Xentry_2413_symbol: Boolean;
          signal Xexit_2414_symbol: Boolean;
          signal word_access_2415_symbol : Boolean;
          signal merge_req_2438_symbol : Boolean;
          signal merge_ack_2439_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_396_complete_2412_start <= ptr_deref_396_active_x_x2382_symbol; -- control passed to block
          Xentry_2413_symbol  <= ptr_deref_396_complete_2412_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/$entry
          word_access_2415: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access 
            signal word_access_2415_start: Boolean;
            signal Xentry_2416_symbol: Boolean;
            signal Xexit_2417_symbol: Boolean;
            signal word_access_0_2418_symbol : Boolean;
            signal word_access_1_2423_symbol : Boolean;
            signal word_access_2_2428_symbol : Boolean;
            signal word_access_3_2433_symbol : Boolean;
            -- 
          begin -- 
            word_access_2415_start <= Xentry_2413_symbol; -- control passed to block
            Xentry_2416_symbol  <= word_access_2415_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/$entry
            word_access_0_2418: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0 
              signal word_access_0_2418_start: Boolean;
              signal Xentry_2419_symbol: Boolean;
              signal Xexit_2420_symbol: Boolean;
              signal cr_2421_symbol : Boolean;
              signal ca_2422_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2418_start <= Xentry_2416_symbol; -- control passed to block
              Xentry_2419_symbol  <= word_access_0_2418_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/$entry
              cr_2421_symbol <= Xentry_2419_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/cr
              ptr_deref_396_load_0_req_1 <= cr_2421_symbol; -- link to DP
              ca_2422_symbol <= ptr_deref_396_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/ca
              Xexit_2420_symbol <= ca_2422_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/$exit
              word_access_0_2418_symbol <= Xexit_2420_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0
            word_access_1_2423: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_1 
              signal word_access_1_2423_start: Boolean;
              signal Xentry_2424_symbol: Boolean;
              signal Xexit_2425_symbol: Boolean;
              signal cr_2426_symbol : Boolean;
              signal ca_2427_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2423_start <= Xentry_2416_symbol; -- control passed to block
              Xentry_2424_symbol  <= word_access_1_2423_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_1/$entry
              cr_2426_symbol <= Xentry_2424_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_1/cr
              ptr_deref_396_load_1_req_1 <= cr_2426_symbol; -- link to DP
              ca_2427_symbol <= ptr_deref_396_load_1_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_1/ca
              Xexit_2425_symbol <= ca_2427_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_1/$exit
              word_access_1_2423_symbol <= Xexit_2425_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_1
            word_access_2_2428: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_2 
              signal word_access_2_2428_start: Boolean;
              signal Xentry_2429_symbol: Boolean;
              signal Xexit_2430_symbol: Boolean;
              signal cr_2431_symbol : Boolean;
              signal ca_2432_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2428_start <= Xentry_2416_symbol; -- control passed to block
              Xentry_2429_symbol  <= word_access_2_2428_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_2/$entry
              cr_2431_symbol <= Xentry_2429_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_2/cr
              ptr_deref_396_load_2_req_1 <= cr_2431_symbol; -- link to DP
              ca_2432_symbol <= ptr_deref_396_load_2_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_2/ca
              Xexit_2430_symbol <= ca_2432_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_2/$exit
              word_access_2_2428_symbol <= Xexit_2430_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_2
            word_access_3_2433: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_3 
              signal word_access_3_2433_start: Boolean;
              signal Xentry_2434_symbol: Boolean;
              signal Xexit_2435_symbol: Boolean;
              signal cr_2436_symbol : Boolean;
              signal ca_2437_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2433_start <= Xentry_2416_symbol; -- control passed to block
              Xentry_2434_symbol  <= word_access_3_2433_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_3/$entry
              cr_2436_symbol <= Xentry_2434_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_3/cr
              ptr_deref_396_load_3_req_1 <= cr_2436_symbol; -- link to DP
              ca_2437_symbol <= ptr_deref_396_load_3_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_3/ca
              Xexit_2435_symbol <= ca_2437_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_3/$exit
              word_access_3_2433_symbol <= Xexit_2435_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_3
            Xexit_2417_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/$exit 
              signal Xexit_2417_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2417_predecessors(0) <= word_access_0_2418_symbol;
              Xexit_2417_predecessors(1) <= word_access_1_2423_symbol;
              Xexit_2417_predecessors(2) <= word_access_2_2428_symbol;
              Xexit_2417_predecessors(3) <= word_access_3_2433_symbol;
              Xexit_2417_join: join -- 
                port map( -- 
                  preds => Xexit_2417_predecessors,
                  symbol_out => Xexit_2417_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/$exit
            word_access_2415_symbol <= Xexit_2417_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access
          merge_req_2438_symbol <= word_access_2415_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/merge_req
          ptr_deref_396_gather_scatter_req_0 <= merge_req_2438_symbol; -- link to DP
          merge_ack_2439_symbol <= ptr_deref_396_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/merge_ack
          Xexit_2414_symbol <= merge_ack_2439_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/$exit
          ptr_deref_396_complete_2412_symbol <= Xexit_2414_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete
        assign_stmt_400_active_x_x2440_symbol <= simple_obj_ref_399_complete_2442_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_400_active_
        assign_stmt_400_completed_x_x2441_symbol <= simple_obj_ref_398_complete_2460_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_400_completed_
        simple_obj_ref_399_complete_2442_symbol <= assign_stmt_397_completed_x_x2380_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_399_complete
        simple_obj_ref_398_trigger_x_x2443_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_trigger_ 
          signal simple_obj_ref_398_trigger_x_x2443_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          simple_obj_ref_398_trigger_x_x2443_predecessors(0) <= simple_obj_ref_398_word_address_calculated_2446_symbol;
          simple_obj_ref_398_trigger_x_x2443_predecessors(1) <= assign_stmt_400_active_x_x2440_symbol;
          simple_obj_ref_398_trigger_x_x2443_predecessors(2) <= simple_obj_ref_379_active_x_x2164_symbol;
          simple_obj_ref_398_trigger_x_x2443_join: join -- 
            port map( -- 
              preds => simple_obj_ref_398_trigger_x_x2443_predecessors,
              symbol_out => simple_obj_ref_398_trigger_x_x2443_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_trigger_
        simple_obj_ref_398_active_x_x2444_symbol <= simple_obj_ref_398_request_2447_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_active_
        simple_obj_ref_398_root_address_calculated_2445_symbol <= Xentry_2087_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_root_address_calculated
        simple_obj_ref_398_word_address_calculated_2446_symbol <= simple_obj_ref_398_root_address_calculated_2445_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_word_address_calculated
        simple_obj_ref_398_request_2447: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request 
          signal simple_obj_ref_398_request_2447_start: Boolean;
          signal Xentry_2448_symbol: Boolean;
          signal Xexit_2449_symbol: Boolean;
          signal split_req_2450_symbol : Boolean;
          signal split_ack_2451_symbol : Boolean;
          signal word_access_2452_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_398_request_2447_start <= simple_obj_ref_398_trigger_x_x2443_symbol; -- control passed to block
          Xentry_2448_symbol  <= simple_obj_ref_398_request_2447_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/$entry
          split_req_2450_symbol <= Xentry_2448_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/split_req
          simple_obj_ref_398_gather_scatter_req_0 <= split_req_2450_symbol; -- link to DP
          split_ack_2451_symbol <= simple_obj_ref_398_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/split_ack
          word_access_2452: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access 
            signal word_access_2452_start: Boolean;
            signal Xentry_2453_symbol: Boolean;
            signal Xexit_2454_symbol: Boolean;
            signal word_access_0_2455_symbol : Boolean;
            -- 
          begin -- 
            word_access_2452_start <= split_ack_2451_symbol; -- control passed to block
            Xentry_2453_symbol  <= word_access_2452_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/$entry
            word_access_0_2455: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0 
              signal word_access_0_2455_start: Boolean;
              signal Xentry_2456_symbol: Boolean;
              signal Xexit_2457_symbol: Boolean;
              signal rr_2458_symbol : Boolean;
              signal ra_2459_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2455_start <= Xentry_2453_symbol; -- control passed to block
              Xentry_2456_symbol  <= word_access_0_2455_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/$entry
              rr_2458_symbol <= Xentry_2456_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/rr
              simple_obj_ref_398_store_0_req_0 <= rr_2458_symbol; -- link to DP
              ra_2459_symbol <= simple_obj_ref_398_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/ra
              Xexit_2457_symbol <= ra_2459_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/$exit
              word_access_0_2455_symbol <= Xexit_2457_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0
            Xexit_2454_symbol <= word_access_0_2455_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/$exit
            word_access_2452_symbol <= Xexit_2454_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access
          Xexit_2449_symbol <= word_access_2452_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/$exit
          simple_obj_ref_398_request_2447_symbol <= Xexit_2449_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request
        simple_obj_ref_398_complete_2460: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete 
          signal simple_obj_ref_398_complete_2460_start: Boolean;
          signal Xentry_2461_symbol: Boolean;
          signal Xexit_2462_symbol: Boolean;
          signal word_access_2463_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_398_complete_2460_start <= simple_obj_ref_398_active_x_x2444_symbol; -- control passed to block
          Xentry_2461_symbol  <= simple_obj_ref_398_complete_2460_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/$entry
          word_access_2463: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access 
            signal word_access_2463_start: Boolean;
            signal Xentry_2464_symbol: Boolean;
            signal Xexit_2465_symbol: Boolean;
            signal word_access_0_2466_symbol : Boolean;
            -- 
          begin -- 
            word_access_2463_start <= Xentry_2461_symbol; -- control passed to block
            Xentry_2464_symbol  <= word_access_2463_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/$entry
            word_access_0_2466: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0 
              signal word_access_0_2466_start: Boolean;
              signal Xentry_2467_symbol: Boolean;
              signal Xexit_2468_symbol: Boolean;
              signal cr_2469_symbol : Boolean;
              signal ca_2470_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2466_start <= Xentry_2464_symbol; -- control passed to block
              Xentry_2467_symbol  <= word_access_0_2466_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/$entry
              cr_2469_symbol <= Xentry_2467_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/cr
              simple_obj_ref_398_store_0_req_1 <= cr_2469_symbol; -- link to DP
              ca_2470_symbol <= simple_obj_ref_398_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/ca
              Xexit_2468_symbol <= ca_2470_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/$exit
              word_access_0_2466_symbol <= Xexit_2468_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0
            Xexit_2465_symbol <= word_access_0_2466_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/$exit
            word_access_2463_symbol <= Xexit_2465_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access
          Xexit_2462_symbol <= word_access_2463_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/$exit
          simple_obj_ref_398_complete_2460_symbol <= Xexit_2462_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete
        Xexit_2088_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/$exit 
          signal Xexit_2088_predecessors: BooleanArray(5 downto 0);
          -- 
        begin -- 
          Xexit_2088_predecessors(0) <= assign_stmt_377_completed_x_x2100_symbol;
          Xexit_2088_predecessors(1) <= ptr_deref_375_base_address_calculated_2104_symbol;
          Xexit_2088_predecessors(2) <= ptr_deref_383_base_address_calculated_2195_symbol;
          Xexit_2088_predecessors(3) <= assign_stmt_393_completed_x_x2275_symbol;
          Xexit_2088_predecessors(4) <= ptr_deref_396_base_address_calculated_2383_symbol;
          Xexit_2088_predecessors(5) <= assign_stmt_400_completed_x_x2441_symbol;
          Xexit_2088_join: join -- 
            port map( -- 
              preds => Xexit_2088_predecessors,
              symbol_out => Xexit_2088_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/$exit
        assign_stmt_373_to_assign_stmt_400_2086_symbol <= Xexit_2088_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400
      bb_0_bb_1_PhiReq_2471: Block -- branch_block_stmt_134/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_2471_start: Boolean;
        signal Xentry_2472_symbol: Boolean;
        signal Xexit_2473_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_2471_start <= bb_0_bb_1_624_symbol; -- control passed to block
        Xentry_2472_symbol  <= bb_0_bb_1_PhiReq_2471_start; -- transition branch_block_stmt_134/bb_0_bb_1_PhiReq/$entry
        Xexit_2473_symbol <= Xentry_2472_symbol; -- transition branch_block_stmt_134/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_2471_symbol <= Xexit_2473_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_0_bb_1_PhiReq
      bb_2_bb_1_PhiReq_2474: Block -- branch_block_stmt_134/bb_2_bb_1_PhiReq 
        signal bb_2_bb_1_PhiReq_2474_start: Boolean;
        signal Xentry_2475_symbol: Boolean;
        signal Xexit_2476_symbol: Boolean;
        -- 
      begin -- 
        bb_2_bb_1_PhiReq_2474_start <= bb_2_bb_1_634_symbol; -- control passed to block
        Xentry_2475_symbol  <= bb_2_bb_1_PhiReq_2474_start; -- transition branch_block_stmt_134/bb_2_bb_1_PhiReq/$entry
        Xexit_2476_symbol <= Xentry_2475_symbol; -- transition branch_block_stmt_134/bb_2_bb_1_PhiReq/$exit
        bb_2_bb_1_PhiReq_2474_symbol <= Xexit_2476_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_2_bb_1_PhiReq
      merge_stmt_160_PhiReqMerge_2477_symbol  <=  bb_0_bb_1_PhiReq_2471_symbol or bb_2_bb_1_PhiReq_2474_symbol; -- place branch_block_stmt_134/merge_stmt_160_PhiReqMerge (optimized away) 
      merge_stmt_160_PhiAck_2478: Block -- branch_block_stmt_134/merge_stmt_160_PhiAck 
        signal merge_stmt_160_PhiAck_2478_start: Boolean;
        signal Xentry_2479_symbol: Boolean;
        signal Xexit_2480_symbol: Boolean;
        signal dummy_2481_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_160_PhiAck_2478_start <= merge_stmt_160_PhiReqMerge_2477_symbol; -- control passed to block
        Xentry_2479_symbol  <= merge_stmt_160_PhiAck_2478_start; -- transition branch_block_stmt_134/merge_stmt_160_PhiAck/$entry
        dummy_2481_symbol <= Xentry_2479_symbol; -- transition branch_block_stmt_134/merge_stmt_160_PhiAck/dummy
        Xexit_2480_symbol <= dummy_2481_symbol; -- transition branch_block_stmt_134/merge_stmt_160_PhiAck/$exit
        merge_stmt_160_PhiAck_2478_symbol <= Xexit_2480_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_160_PhiAck
      merge_stmt_180_dead_link_2482: Block -- branch_block_stmt_134/merge_stmt_180_dead_link 
        signal merge_stmt_180_dead_link_2482_start: Boolean;
        signal Xentry_2483_symbol: Boolean;
        signal Xexit_2484_symbol: Boolean;
        signal dead_transition_2485_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_180_dead_link_2482_start <= merge_stmt_180_x_xentry_x_xx_x630_symbol; -- control passed to block
        Xentry_2483_symbol  <= merge_stmt_180_dead_link_2482_start; -- transition branch_block_stmt_134/merge_stmt_180_dead_link/$entry
        dead_transition_2485_symbol <= false;
        Xexit_2484_symbol <= dead_transition_2485_symbol; -- transition branch_block_stmt_134/merge_stmt_180_dead_link/$exit
        merge_stmt_180_dead_link_2482_symbol <= Xexit_2484_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_180_dead_link
      bb_1_bb_2_PhiReq_2486: Block -- branch_block_stmt_134/bb_1_bb_2_PhiReq 
        signal bb_1_bb_2_PhiReq_2486_start: Boolean;
        signal Xentry_2487_symbol: Boolean;
        signal Xexit_2488_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_2_PhiReq_2486_start <= bb_1_bb_2_845_symbol; -- control passed to block
        Xentry_2487_symbol  <= bb_1_bb_2_PhiReq_2486_start; -- transition branch_block_stmt_134/bb_1_bb_2_PhiReq/$entry
        Xexit_2488_symbol <= Xentry_2487_symbol; -- transition branch_block_stmt_134/bb_1_bb_2_PhiReq/$exit
        bb_1_bb_2_PhiReq_2486_symbol <= Xexit_2488_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_1_bb_2_PhiReq
      merge_stmt_180_PhiReqMerge_2489_symbol  <=  bb_1_bb_2_PhiReq_2486_symbol; -- place branch_block_stmt_134/merge_stmt_180_PhiReqMerge (optimized away) 
      merge_stmt_180_PhiAck_2490: Block -- branch_block_stmt_134/merge_stmt_180_PhiAck 
        signal merge_stmt_180_PhiAck_2490_start: Boolean;
        signal Xentry_2491_symbol: Boolean;
        signal Xexit_2492_symbol: Boolean;
        signal dummy_2493_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_180_PhiAck_2490_start <= merge_stmt_180_PhiReqMerge_2489_symbol; -- control passed to block
        Xentry_2491_symbol  <= merge_stmt_180_PhiAck_2490_start; -- transition branch_block_stmt_134/merge_stmt_180_PhiAck/$entry
        dummy_2493_symbol <= Xentry_2491_symbol; -- transition branch_block_stmt_134/merge_stmt_180_PhiAck/dummy
        Xexit_2492_symbol <= dummy_2493_symbol; -- transition branch_block_stmt_134/merge_stmt_180_PhiAck/$exit
        merge_stmt_180_PhiAck_2490_symbol <= Xexit_2492_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_180_PhiAck
      bb_1_bb_3_PhiReq_2494: Block -- branch_block_stmt_134/bb_1_bb_3_PhiReq 
        signal bb_1_bb_3_PhiReq_2494_start: Boolean;
        signal Xentry_2495_symbol: Boolean;
        signal Xexit_2496_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_3_PhiReq_2494_start <= bb_1_bb_3_846_symbol; -- control passed to block
        Xentry_2495_symbol  <= bb_1_bb_3_PhiReq_2494_start; -- transition branch_block_stmt_134/bb_1_bb_3_PhiReq/$entry
        Xexit_2496_symbol <= Xentry_2495_symbol; -- transition branch_block_stmt_134/bb_1_bb_3_PhiReq/$exit
        bb_1_bb_3_PhiReq_2494_symbol <= Xexit_2496_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_1_bb_3_PhiReq
      merge_stmt_227_PhiReqMerge_2497_symbol  <=  bb_1_bb_3_PhiReq_2494_symbol; -- place branch_block_stmt_134/merge_stmt_227_PhiReqMerge (optimized away) 
      merge_stmt_227_PhiAck_2498: Block -- branch_block_stmt_134/merge_stmt_227_PhiAck 
        signal merge_stmt_227_PhiAck_2498_start: Boolean;
        signal Xentry_2499_symbol: Boolean;
        signal Xexit_2500_symbol: Boolean;
        signal dummy_2501_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_227_PhiAck_2498_start <= merge_stmt_227_PhiReqMerge_2497_symbol; -- control passed to block
        Xentry_2499_symbol  <= merge_stmt_227_PhiAck_2498_start; -- transition branch_block_stmt_134/merge_stmt_227_PhiAck/$entry
        dummy_2501_symbol <= Xentry_2499_symbol; -- transition branch_block_stmt_134/merge_stmt_227_PhiAck/dummy
        Xexit_2500_symbol <= dummy_2501_symbol; -- transition branch_block_stmt_134/merge_stmt_227_PhiAck/$exit
        merge_stmt_227_PhiAck_2498_symbol <= Xexit_2500_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_227_PhiAck
      bb_3_bb_4_PhiReq_2502: Block -- branch_block_stmt_134/bb_3_bb_4_PhiReq 
        signal bb_3_bb_4_PhiReq_2502_start: Boolean;
        signal Xentry_2503_symbol: Boolean;
        signal Xexit_2504_symbol: Boolean;
        -- 
      begin -- 
        bb_3_bb_4_PhiReq_2502_start <= bb_3_bb_4_638_symbol; -- control passed to block
        Xentry_2503_symbol  <= bb_3_bb_4_PhiReq_2502_start; -- transition branch_block_stmt_134/bb_3_bb_4_PhiReq/$entry
        Xexit_2504_symbol <= Xentry_2503_symbol; -- transition branch_block_stmt_134/bb_3_bb_4_PhiReq/$exit
        bb_3_bb_4_PhiReq_2502_symbol <= Xexit_2504_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_3_bb_4_PhiReq
      bb_7_bb_4_PhiReq_2505: Block -- branch_block_stmt_134/bb_7_bb_4_PhiReq 
        signal bb_7_bb_4_PhiReq_2505_start: Boolean;
        signal Xentry_2506_symbol: Boolean;
        signal Xexit_2507_symbol: Boolean;
        -- 
      begin -- 
        bb_7_bb_4_PhiReq_2505_start <= bb_7_bb_4_664_symbol; -- control passed to block
        Xentry_2506_symbol  <= bb_7_bb_4_PhiReq_2505_start; -- transition branch_block_stmt_134/bb_7_bb_4_PhiReq/$entry
        Xexit_2507_symbol <= Xentry_2506_symbol; -- transition branch_block_stmt_134/bb_7_bb_4_PhiReq/$exit
        bb_7_bb_4_PhiReq_2505_symbol <= Xexit_2507_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_7_bb_4_PhiReq
      bb_8_bb_4_PhiReq_2508: Block -- branch_block_stmt_134/bb_8_bb_4_PhiReq 
        signal bb_8_bb_4_PhiReq_2508_start: Boolean;
        signal Xentry_2509_symbol: Boolean;
        signal Xexit_2510_symbol: Boolean;
        -- 
      begin -- 
        bb_8_bb_4_PhiReq_2508_start <= bb_8_bb_4_2064_symbol; -- control passed to block
        Xentry_2509_symbol  <= bb_8_bb_4_PhiReq_2508_start; -- transition branch_block_stmt_134/bb_8_bb_4_PhiReq/$entry
        Xexit_2510_symbol <= Xentry_2509_symbol; -- transition branch_block_stmt_134/bb_8_bb_4_PhiReq/$exit
        bb_8_bb_4_PhiReq_2508_symbol <= Xexit_2510_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_8_bb_4_PhiReq
      bb_9_bb_4_PhiReq_2511: Block -- branch_block_stmt_134/bb_9_bb_4_PhiReq 
        signal bb_9_bb_4_PhiReq_2511_start: Boolean;
        signal Xentry_2512_symbol: Boolean;
        signal Xexit_2513_symbol: Boolean;
        -- 
      begin -- 
        bb_9_bb_4_PhiReq_2511_start <= bb_9_bb_4_678_symbol; -- control passed to block
        Xentry_2512_symbol  <= bb_9_bb_4_PhiReq_2511_start; -- transition branch_block_stmt_134/bb_9_bb_4_PhiReq/$entry
        Xexit_2513_symbol <= Xentry_2512_symbol; -- transition branch_block_stmt_134/bb_9_bb_4_PhiReq/$exit
        bb_9_bb_4_PhiReq_2511_symbol <= Xexit_2513_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_9_bb_4_PhiReq
      merge_stmt_247_PhiReqMerge_2514_symbol  <=  bb_3_bb_4_PhiReq_2502_symbol or bb_7_bb_4_PhiReq_2505_symbol or bb_8_bb_4_PhiReq_2508_symbol or bb_9_bb_4_PhiReq_2511_symbol; -- place branch_block_stmt_134/merge_stmt_247_PhiReqMerge (optimized away) 
      merge_stmt_247_PhiAck_2515: Block -- branch_block_stmt_134/merge_stmt_247_PhiAck 
        signal merge_stmt_247_PhiAck_2515_start: Boolean;
        signal Xentry_2516_symbol: Boolean;
        signal Xexit_2517_symbol: Boolean;
        signal dummy_2518_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_247_PhiAck_2515_start <= merge_stmt_247_PhiReqMerge_2514_symbol; -- control passed to block
        Xentry_2516_symbol  <= merge_stmt_247_PhiAck_2515_start; -- transition branch_block_stmt_134/merge_stmt_247_PhiAck/$entry
        dummy_2518_symbol <= Xentry_2516_symbol; -- transition branch_block_stmt_134/merge_stmt_247_PhiAck/dummy
        Xexit_2517_symbol <= dummy_2518_symbol; -- transition branch_block_stmt_134/merge_stmt_247_PhiAck/$exit
        merge_stmt_247_PhiAck_2515_symbol <= Xexit_2517_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_247_PhiAck
      merge_stmt_280_dead_link_2519: Block -- branch_block_stmt_134/merge_stmt_280_dead_link 
        signal merge_stmt_280_dead_link_2519_start: Boolean;
        signal Xentry_2520_symbol: Boolean;
        signal Xexit_2521_symbol: Boolean;
        signal dead_transition_2522_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_280_dead_link_2519_start <= merge_stmt_280_x_xentry_x_xx_x648_symbol; -- control passed to block
        Xentry_2520_symbol  <= merge_stmt_280_dead_link_2519_start; -- transition branch_block_stmt_134/merge_stmt_280_dead_link/$entry
        dead_transition_2522_symbol <= false;
        Xexit_2521_symbol <= dead_transition_2522_symbol; -- transition branch_block_stmt_134/merge_stmt_280_dead_link/$exit
        merge_stmt_280_dead_link_2519_symbol <= Xexit_2521_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_280_dead_link
      bb_4_bb_5_PhiReq_2523: Block -- branch_block_stmt_134/bb_4_bb_5_PhiReq 
        signal bb_4_bb_5_PhiReq_2523_start: Boolean;
        signal Xentry_2524_symbol: Boolean;
        signal Xexit_2525_symbol: Boolean;
        -- 
      begin -- 
        bb_4_bb_5_PhiReq_2523_start <= bb_4_bb_5_1540_symbol; -- control passed to block
        Xentry_2524_symbol  <= bb_4_bb_5_PhiReq_2523_start; -- transition branch_block_stmt_134/bb_4_bb_5_PhiReq/$entry
        Xexit_2525_symbol <= Xentry_2524_symbol; -- transition branch_block_stmt_134/bb_4_bb_5_PhiReq/$exit
        bb_4_bb_5_PhiReq_2523_symbol <= Xexit_2525_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_4_bb_5_PhiReq
      merge_stmt_280_PhiReqMerge_2526_symbol  <=  bb_4_bb_5_PhiReq_2523_symbol; -- place branch_block_stmt_134/merge_stmt_280_PhiReqMerge (optimized away) 
      merge_stmt_280_PhiAck_2527: Block -- branch_block_stmt_134/merge_stmt_280_PhiAck 
        signal merge_stmt_280_PhiAck_2527_start: Boolean;
        signal Xentry_2528_symbol: Boolean;
        signal Xexit_2529_symbol: Boolean;
        signal dummy_2530_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_280_PhiAck_2527_start <= merge_stmt_280_PhiReqMerge_2526_symbol; -- control passed to block
        Xentry_2528_symbol  <= merge_stmt_280_PhiAck_2527_start; -- transition branch_block_stmt_134/merge_stmt_280_PhiAck/$entry
        dummy_2530_symbol <= Xentry_2528_symbol; -- transition branch_block_stmt_134/merge_stmt_280_PhiAck/dummy
        Xexit_2529_symbol <= dummy_2530_symbol; -- transition branch_block_stmt_134/merge_stmt_280_PhiAck/$exit
        merge_stmt_280_PhiAck_2527_symbol <= Xexit_2529_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_280_PhiAck
      merge_stmt_304_dead_link_2531: Block -- branch_block_stmt_134/merge_stmt_304_dead_link 
        signal merge_stmt_304_dead_link_2531_start: Boolean;
        signal Xentry_2532_symbol: Boolean;
        signal Xexit_2533_symbol: Boolean;
        signal dead_transition_2534_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_304_dead_link_2531_start <= merge_stmt_304_x_xentry_x_xx_x654_symbol; -- control passed to block
        Xentry_2532_symbol  <= merge_stmt_304_dead_link_2531_start; -- transition branch_block_stmt_134/merge_stmt_304_dead_link/$entry
        dead_transition_2534_symbol <= false;
        Xexit_2533_symbol <= dead_transition_2534_symbol; -- transition branch_block_stmt_134/merge_stmt_304_dead_link/$exit
        merge_stmt_304_dead_link_2531_symbol <= Xexit_2533_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_304_dead_link
      bb_5_bb_6_PhiReq_2535: Block -- branch_block_stmt_134/bb_5_bb_6_PhiReq 
        signal bb_5_bb_6_PhiReq_2535_start: Boolean;
        signal Xentry_2536_symbol: Boolean;
        signal Xexit_2537_symbol: Boolean;
        -- 
      begin -- 
        bb_5_bb_6_PhiReq_2535_start <= bb_5_bb_6_1705_symbol; -- control passed to block
        Xentry_2536_symbol  <= bb_5_bb_6_PhiReq_2535_start; -- transition branch_block_stmt_134/bb_5_bb_6_PhiReq/$entry
        Xexit_2537_symbol <= Xentry_2536_symbol; -- transition branch_block_stmt_134/bb_5_bb_6_PhiReq/$exit
        bb_5_bb_6_PhiReq_2535_symbol <= Xexit_2537_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_5_bb_6_PhiReq
      merge_stmt_304_PhiReqMerge_2538_symbol  <=  bb_5_bb_6_PhiReq_2535_symbol; -- place branch_block_stmt_134/merge_stmt_304_PhiReqMerge (optimized away) 
      merge_stmt_304_PhiAck_2539: Block -- branch_block_stmt_134/merge_stmt_304_PhiAck 
        signal merge_stmt_304_PhiAck_2539_start: Boolean;
        signal Xentry_2540_symbol: Boolean;
        signal Xexit_2541_symbol: Boolean;
        signal dummy_2542_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_304_PhiAck_2539_start <= merge_stmt_304_PhiReqMerge_2538_symbol; -- control passed to block
        Xentry_2540_symbol  <= merge_stmt_304_PhiAck_2539_start; -- transition branch_block_stmt_134/merge_stmt_304_PhiAck/$entry
        dummy_2542_symbol <= Xentry_2540_symbol; -- transition branch_block_stmt_134/merge_stmt_304_PhiAck/dummy
        Xexit_2541_symbol <= dummy_2542_symbol; -- transition branch_block_stmt_134/merge_stmt_304_PhiAck/$exit
        merge_stmt_304_PhiAck_2539_symbol <= Xexit_2541_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_304_PhiAck
      bb_5_bb_7_PhiReq_2543: Block -- branch_block_stmt_134/bb_5_bb_7_PhiReq 
        signal bb_5_bb_7_PhiReq_2543_start: Boolean;
        signal Xentry_2544_symbol: Boolean;
        signal Xexit_2545_symbol: Boolean;
        -- 
      begin -- 
        bb_5_bb_7_PhiReq_2543_start <= bb_5_bb_7_1706_symbol; -- control passed to block
        Xentry_2544_symbol  <= bb_5_bb_7_PhiReq_2543_start; -- transition branch_block_stmt_134/bb_5_bb_7_PhiReq/$entry
        Xexit_2545_symbol <= Xentry_2544_symbol; -- transition branch_block_stmt_134/bb_5_bb_7_PhiReq/$exit
        bb_5_bb_7_PhiReq_2543_symbol <= Xexit_2545_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_5_bb_7_PhiReq
      bb_6_bb_7_PhiReq_2546: Block -- branch_block_stmt_134/bb_6_bb_7_PhiReq 
        signal bb_6_bb_7_PhiReq_2546_start: Boolean;
        signal Xentry_2547_symbol: Boolean;
        signal Xexit_2548_symbol: Boolean;
        -- 
      begin -- 
        bb_6_bb_7_PhiReq_2546_start <= bb_6_bb_7_658_symbol; -- control passed to block
        Xentry_2547_symbol  <= bb_6_bb_7_PhiReq_2546_start; -- transition branch_block_stmt_134/bb_6_bb_7_PhiReq/$entry
        Xexit_2548_symbol <= Xentry_2547_symbol; -- transition branch_block_stmt_134/bb_6_bb_7_PhiReq/$exit
        bb_6_bb_7_PhiReq_2546_symbol <= Xexit_2548_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_6_bb_7_PhiReq
      merge_stmt_321_PhiReqMerge_2549_symbol  <=  bb_5_bb_7_PhiReq_2543_symbol or bb_6_bb_7_PhiReq_2546_symbol; -- place branch_block_stmt_134/merge_stmt_321_PhiReqMerge (optimized away) 
      merge_stmt_321_PhiAck_2550: Block -- branch_block_stmt_134/merge_stmt_321_PhiAck 
        signal merge_stmt_321_PhiAck_2550_start: Boolean;
        signal Xentry_2551_symbol: Boolean;
        signal Xexit_2552_symbol: Boolean;
        signal dummy_2553_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_321_PhiAck_2550_start <= merge_stmt_321_PhiReqMerge_2549_symbol; -- control passed to block
        Xentry_2551_symbol  <= merge_stmt_321_PhiAck_2550_start; -- transition branch_block_stmt_134/merge_stmt_321_PhiAck/$entry
        dummy_2553_symbol <= Xentry_2551_symbol; -- transition branch_block_stmt_134/merge_stmt_321_PhiAck/dummy
        Xexit_2552_symbol <= dummy_2553_symbol; -- transition branch_block_stmt_134/merge_stmt_321_PhiAck/$exit
        merge_stmt_321_PhiAck_2550_symbol <= Xexit_2552_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_321_PhiAck
      bb_4_bb_8_PhiReq_2554: Block -- branch_block_stmt_134/bb_4_bb_8_PhiReq 
        signal bb_4_bb_8_PhiReq_2554_start: Boolean;
        signal Xentry_2555_symbol: Boolean;
        signal Xexit_2556_symbol: Boolean;
        -- 
      begin -- 
        bb_4_bb_8_PhiReq_2554_start <= bb_4_bb_8_1541_symbol; -- control passed to block
        Xentry_2555_symbol  <= bb_4_bb_8_PhiReq_2554_start; -- transition branch_block_stmt_134/bb_4_bb_8_PhiReq/$entry
        Xexit_2556_symbol <= Xentry_2555_symbol; -- transition branch_block_stmt_134/bb_4_bb_8_PhiReq/$exit
        bb_4_bb_8_PhiReq_2554_symbol <= Xexit_2556_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_4_bb_8_PhiReq
      merge_stmt_340_PhiReqMerge_2557_symbol  <=  bb_4_bb_8_PhiReq_2554_symbol; -- place branch_block_stmt_134/merge_stmt_340_PhiReqMerge (optimized away) 
      merge_stmt_340_PhiAck_2558: Block -- branch_block_stmt_134/merge_stmt_340_PhiAck 
        signal merge_stmt_340_PhiAck_2558_start: Boolean;
        signal Xentry_2559_symbol: Boolean;
        signal Xexit_2560_symbol: Boolean;
        signal dummy_2561_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_340_PhiAck_2558_start <= merge_stmt_340_PhiReqMerge_2557_symbol; -- control passed to block
        Xentry_2559_symbol  <= merge_stmt_340_PhiAck_2558_start; -- transition branch_block_stmt_134/merge_stmt_340_PhiAck/$entry
        dummy_2561_symbol <= Xentry_2559_symbol; -- transition branch_block_stmt_134/merge_stmt_340_PhiAck/dummy
        Xexit_2560_symbol <= dummy_2561_symbol; -- transition branch_block_stmt_134/merge_stmt_340_PhiAck/$exit
        merge_stmt_340_PhiAck_2558_symbol <= Xexit_2560_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_340_PhiAck
      merge_stmt_360_dead_link_2562: Block -- branch_block_stmt_134/merge_stmt_360_dead_link 
        signal merge_stmt_360_dead_link_2562_start: Boolean;
        signal Xentry_2563_symbol: Boolean;
        signal Xexit_2564_symbol: Boolean;
        signal dead_transition_2565_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_360_dead_link_2562_start <= merge_stmt_360_x_xentry_x_xx_x670_symbol; -- control passed to block
        Xentry_2563_symbol  <= merge_stmt_360_dead_link_2562_start; -- transition branch_block_stmt_134/merge_stmt_360_dead_link/$entry
        dead_transition_2565_symbol <= false;
        Xexit_2564_symbol <= dead_transition_2565_symbol; -- transition branch_block_stmt_134/merge_stmt_360_dead_link/$exit
        merge_stmt_360_dead_link_2562_symbol <= Xexit_2564_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_360_dead_link
      bb_8_bb_9_PhiReq_2566: Block -- branch_block_stmt_134/bb_8_bb_9_PhiReq 
        signal bb_8_bb_9_PhiReq_2566_start: Boolean;
        signal Xentry_2567_symbol: Boolean;
        signal Xexit_2568_symbol: Boolean;
        -- 
      begin -- 
        bb_8_bb_9_PhiReq_2566_start <= bb_8_bb_9_2063_symbol; -- control passed to block
        Xentry_2567_symbol  <= bb_8_bb_9_PhiReq_2566_start; -- transition branch_block_stmt_134/bb_8_bb_9_PhiReq/$entry
        Xexit_2568_symbol <= Xentry_2567_symbol; -- transition branch_block_stmt_134/bb_8_bb_9_PhiReq/$exit
        bb_8_bb_9_PhiReq_2566_symbol <= Xexit_2568_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_8_bb_9_PhiReq
      merge_stmt_360_PhiReqMerge_2569_symbol  <=  bb_8_bb_9_PhiReq_2566_symbol; -- place branch_block_stmt_134/merge_stmt_360_PhiReqMerge (optimized away) 
      merge_stmt_360_PhiAck_2570: Block -- branch_block_stmt_134/merge_stmt_360_PhiAck 
        signal merge_stmt_360_PhiAck_2570_start: Boolean;
        signal Xentry_2571_symbol: Boolean;
        signal Xexit_2572_symbol: Boolean;
        signal dummy_2573_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_360_PhiAck_2570_start <= merge_stmt_360_PhiReqMerge_2569_symbol; -- control passed to block
        Xentry_2571_symbol  <= merge_stmt_360_PhiAck_2570_start; -- transition branch_block_stmt_134/merge_stmt_360_PhiAck/$entry
        dummy_2573_symbol <= Xentry_2571_symbol; -- transition branch_block_stmt_134/merge_stmt_360_PhiAck/dummy
        Xexit_2572_symbol <= dummy_2573_symbol; -- transition branch_block_stmt_134/merge_stmt_360_PhiAck/$exit
        merge_stmt_360_PhiAck_2570_symbol <= Xexit_2572_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_360_PhiAck
      Xexit_619_symbol <= branch_block_stmt_134_x_xexit_x_xx_x621_symbol; -- transition branch_block_stmt_134/$exit
      branch_block_stmt_134_617_symbol <= Xexit_619_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_134
    Xexit_616_symbol <= branch_block_stmt_134_617_symbol; -- transition $exit
    fin  <=  '1' when Xexit_616_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_192_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_192_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_192_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_192_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_201_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_201_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_201_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_201_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_207_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_207_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_311_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_311_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_388_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_388_root_address : std_logic_vector(5 downto 0);
    signal command_146 : std_logic_vector(31 downto 0);
    signal expr_157_wire_constant : std_logic_vector(31 downto 0);
    signal expr_187_wire_constant : std_logic_vector(31 downto 0);
    signal expr_219_wire_constant : std_logic_vector(31 downto 0);
    signal expr_236_wire_constant : std_logic_vector(31 downto 0);
    signal expr_271_wire_constant : std_logic_vector(31 downto 0);
    signal expr_351_wire_constant : std_logic_vector(31 downto 0);
    signal iNsTr_10_208 : std_logic_vector(31 downto 0);
    signal iNsTr_12_216 : std_logic_vector(31 downto 0);
    signal iNsTr_13_221 : std_logic_vector(31 downto 0);
    signal iNsTr_16_233 : std_logic_vector(31 downto 0);
    signal iNsTr_18_242 : std_logic_vector(31 downto 0);
    signal iNsTr_21_252 : std_logic_vector(31 downto 0);
    signal iNsTr_22_256 : std_logic_vector(7 downto 0);
    signal iNsTr_24_264 : std_logic_vector(7 downto 0);
    signal iNsTr_25_268 : std_logic_vector(31 downto 0);
    signal iNsTr_26_273 : std_logic_vector(0 downto 0);
    signal iNsTr_28_283 : std_logic_vector(31 downto 0);
    signal iNsTr_2_164 : std_logic_vector(31 downto 0);
    signal iNsTr_30_290 : std_logic_vector(31 downto 0);
    signal iNsTr_31_297 : std_logic_vector(0 downto 0);
    signal iNsTr_33_344 : std_logic_vector(7 downto 0);
    signal iNsTr_34_348 : std_logic_vector(31 downto 0);
    signal iNsTr_35_353 : std_logic_vector(0 downto 0);
    signal iNsTr_37_307 : std_logic_vector(31 downto 0);
    signal iNsTr_38_312 : std_logic_vector(31 downto 0);
    signal iNsTr_39_316 : std_logic_vector(31 downto 0);
    signal iNsTr_3_173 : std_logic_vector(0 downto 0);
    signal iNsTr_42_325 : std_logic_vector(31 downto 0);
    signal iNsTr_43_329 : std_logic_vector(31 downto 0);
    signal iNsTr_44_334 : std_logic_vector(31 downto 0);
    signal iNsTr_47_365 : std_logic_vector(31 downto 0);
    signal iNsTr_48_369 : std_logic_vector(31 downto 0);
    signal iNsTr_49_373 : std_logic_vector(31 downto 0);
    signal iNsTr_51_380 : std_logic_vector(31 downto 0);
    signal iNsTr_52_384 : std_logic_vector(31 downto 0);
    signal iNsTr_53_389 : std_logic_vector(31 downto 0);
    signal iNsTr_55_397 : std_logic_vector(31 downto 0);
    signal iNsTr_5_184 : std_logic_vector(31 downto 0);
    signal iNsTr_6_189 : std_logic_vector(31 downto 0);
    signal iNsTr_7_194 : std_logic_vector(31 downto 0);
    signal iNsTr_8_198 : std_logic_vector(31 downto 0);
    signal iNsTr_9_203 : std_logic_vector(31 downto 0);
    signal i_142 : std_logic_vector(31 downto 0);
    signal ptr_deref_156_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_156_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_156_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_156_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_156_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_156_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_156_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_156_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_156_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_163_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_163_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_163_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_163_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_163_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_163_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_163_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_163_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_183_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_183_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_183_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_183_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_183_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_183_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_183_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_183_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_197_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_197_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_197_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_197_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_197_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_197_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_197_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_197_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_210_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_210_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_210_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_210_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_210_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_210_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_210_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_210_word_offset_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_215_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_215_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_215_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_215_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_215_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_215_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_215_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_215_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_223_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_223_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_223_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_223_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_223_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_223_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_223_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_223_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_223_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_235_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_235_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_235_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_235_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_235_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_235_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_235_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_235_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_235_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_258_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_258_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_258_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_263_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_263_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_285_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_285_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_285_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_285_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_285_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_285_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_285_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_285_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_285_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_315_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_315_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_315_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_315_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_315_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_315_word_offset_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_324_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_324_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_324_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_324_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_324_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_324_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_324_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_324_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_343_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_343_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_375_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_375_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_375_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_375_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_375_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_375_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_375_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_375_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_375_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_383_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_383_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_383_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_383_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_383_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_383_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_383_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_383_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_391_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_391_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_391_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_391_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_391_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_391_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_391_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_391_word_offset_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_396_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_396_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_396_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_396_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_396_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_396_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_396_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_396_word_address_3 : std_logic_vector(5 downto 0);
    signal put_link_154 : std_logic_vector(31 downto 0);
    signal ret_150 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_191_resized : std_logic_vector(5 downto 0);
    signal simple_obj_ref_191_scaled : std_logic_vector(5 downto 0);
    signal simple_obj_ref_200_resized : std_logic_vector(5 downto 0);
    signal simple_obj_ref_200_scaled : std_logic_vector(5 downto 0);
    signal simple_obj_ref_243_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_243_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_254_wire : std_logic_vector(7 downto 0);
    signal simple_obj_ref_282_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_282_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_289_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_289_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_306_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_306_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_317_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_317_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_367_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_379_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_379_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_398_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_398_word_address_0 : std_logic_vector(0 downto 0);
    signal type_cast_168_wire : std_logic_vector(31 downto 0);
    signal type_cast_170_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_293_wire : std_logic_vector(31 downto 0);
    signal type_cast_295_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_337_wire : std_logic_vector(31 downto 0);
    signal xxfree_queue_managerxxbodyxxcommand_alloc_base_address : std_logic_vector(5 downto 0);
    signal xxfree_queue_managerxxbodyxxi_alloc_base_address : std_logic_vector(5 downto 0);
    signal xxfree_queue_managerxxbodyxxput_link_alloc_base_address : std_logic_vector(5 downto 0);
    signal xxfree_queue_managerxxbodyxxret_alloc_base_address : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    array_obj_ref_192_offset_scale_factor_0 <= "001000";
    array_obj_ref_192_resized_base_address <= "000000";
    array_obj_ref_201_offset_scale_factor_0 <= "001000";
    array_obj_ref_201_resized_base_address <= "000000";
    command_146 <= "00000000000000000000000000100000";
    expr_157_wire_constant <= "00000000000000000000000000000001";
    expr_187_wire_constant <= "00000000000000000000000000000001";
    expr_219_wire_constant <= "00000000000000000000000000000001";
    expr_236_wire_constant <= "00000000000000000000000000000000";
    expr_271_wire_constant <= "00000000000000000000000000000010";
    expr_351_wire_constant <= "00000000000000000000000000000001";
    iNsTr_16_233 <= "00000000000000000000000000010000";
    iNsTr_18_242 <= "00000000000000000000000000001000";
    iNsTr_21_252 <= "00000000000000000000000000000000";
    iNsTr_44_334 <= "00000000000000000000000000000000";
    iNsTr_47_365 <= "00000000000000000000000000000000";
    i_142 <= "00000000000000000000000000011100";
    ptr_deref_156_word_address_0 <= "011100";
    ptr_deref_156_word_address_1 <= "011101";
    ptr_deref_156_word_address_2 <= "011110";
    ptr_deref_156_word_address_3 <= "011111";
    ptr_deref_163_word_address_0 <= "011100";
    ptr_deref_163_word_address_1 <= "011101";
    ptr_deref_163_word_address_2 <= "011110";
    ptr_deref_163_word_address_3 <= "011111";
    ptr_deref_183_word_address_0 <= "011100";
    ptr_deref_183_word_address_1 <= "011101";
    ptr_deref_183_word_address_2 <= "011110";
    ptr_deref_183_word_address_3 <= "011111";
    ptr_deref_197_word_address_0 <= "011100";
    ptr_deref_197_word_address_1 <= "011101";
    ptr_deref_197_word_address_2 <= "011110";
    ptr_deref_197_word_address_3 <= "011111";
    ptr_deref_210_word_offset_0 <= "000000";
    ptr_deref_210_word_offset_1 <= "000001";
    ptr_deref_210_word_offset_2 <= "000010";
    ptr_deref_210_word_offset_3 <= "000011";
    ptr_deref_215_word_address_0 <= "011100";
    ptr_deref_215_word_address_1 <= "011101";
    ptr_deref_215_word_address_2 <= "011110";
    ptr_deref_215_word_address_3 <= "011111";
    ptr_deref_223_word_address_0 <= "011100";
    ptr_deref_223_word_address_1 <= "011101";
    ptr_deref_223_word_address_2 <= "011110";
    ptr_deref_223_word_address_3 <= "011111";
    ptr_deref_235_word_address_0 <= "010000";
    ptr_deref_235_word_address_1 <= "010001";
    ptr_deref_235_word_address_2 <= "010010";
    ptr_deref_235_word_address_3 <= "010011";
    ptr_deref_258_word_address_0 <= "100000";
    ptr_deref_263_word_address_0 <= "100000";
    ptr_deref_285_word_address_0 <= "100001";
    ptr_deref_285_word_address_1 <= "100010";
    ptr_deref_285_word_address_2 <= "100011";
    ptr_deref_285_word_address_3 <= "100100";
    ptr_deref_315_word_offset_0 <= "000000";
    ptr_deref_315_word_offset_1 <= "000001";
    ptr_deref_315_word_offset_2 <= "000010";
    ptr_deref_315_word_offset_3 <= "000011";
    ptr_deref_324_word_address_0 <= "100001";
    ptr_deref_324_word_address_1 <= "100010";
    ptr_deref_324_word_address_2 <= "100011";
    ptr_deref_324_word_address_3 <= "100100";
    ptr_deref_343_word_address_0 <= "100000";
    ptr_deref_375_word_address_0 <= "100101";
    ptr_deref_375_word_address_1 <= "100110";
    ptr_deref_375_word_address_2 <= "100111";
    ptr_deref_375_word_address_3 <= "101000";
    ptr_deref_383_word_address_0 <= "100101";
    ptr_deref_383_word_address_1 <= "100110";
    ptr_deref_383_word_address_2 <= "100111";
    ptr_deref_383_word_address_3 <= "101000";
    ptr_deref_391_word_offset_0 <= "000000";
    ptr_deref_391_word_offset_1 <= "000001";
    ptr_deref_391_word_offset_2 <= "000010";
    ptr_deref_391_word_offset_3 <= "000011";
    ptr_deref_396_word_address_0 <= "100101";
    ptr_deref_396_word_address_1 <= "100110";
    ptr_deref_396_word_address_2 <= "100111";
    ptr_deref_396_word_address_3 <= "101000";
    put_link_154 <= "00000000000000000000000000100101";
    ret_150 <= "00000000000000000000000000100001";
    simple_obj_ref_243_word_address_0 <= "0";
    simple_obj_ref_282_word_address_0 <= "0";
    simple_obj_ref_289_word_address_0 <= "0";
    simple_obj_ref_306_word_address_0 <= "0";
    simple_obj_ref_317_word_address_0 <= "0";
    simple_obj_ref_379_word_address_0 <= "0";
    simple_obj_ref_398_word_address_0 <= "0";
    type_cast_170_wire_constant <= "00000000000000000000000000000010";
    type_cast_295_wire_constant <= "00000000000000000000000000000000";
    xxfree_queue_managerxxbodyxxcommand_alloc_base_address <= "100000";
    xxfree_queue_managerxxbodyxxi_alloc_base_address <= "011100";
    xxfree_queue_managerxxbodyxxput_link_alloc_base_address <= "100101";
    xxfree_queue_managerxxbodyxxret_alloc_base_address <= "100001";
    addr_of_193_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_192_root_address, dout => iNsTr_7_194, req => addr_of_193_final_reg_req_0, ack => addr_of_193_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_202_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_201_root_address, dout => iNsTr_9_203, req => addr_of_202_final_reg_req_0, ack => addr_of_202_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_192_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_6_189, dout => simple_obj_ref_191_resized, req => array_obj_ref_192_index_0_resize_req_0, ack => array_obj_ref_192_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_192_offset_inst: RegisterBase generic map(in_data_width => 6,out_data_width => 6) -- 
      port map( din => simple_obj_ref_191_scaled, dout => array_obj_ref_192_final_offset, req => array_obj_ref_192_offset_inst_req_0, ack => array_obj_ref_192_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_201_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_8_198, dout => simple_obj_ref_200_resized, req => array_obj_ref_201_index_0_resize_req_0, ack => array_obj_ref_201_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_201_offset_inst: RegisterBase generic map(in_data_width => 6,out_data_width => 6) -- 
      port map( din => simple_obj_ref_200_scaled, dout => array_obj_ref_201_final_offset, req => array_obj_ref_201_offset_inst_req_0, ack => array_obj_ref_201_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_207_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_9_203, dout => array_obj_ref_207_resized_base_address, req => array_obj_ref_207_base_resize_req_0, ack => array_obj_ref_207_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_207_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_207_root_address, dout => iNsTr_10_208, req => array_obj_ref_207_final_reg_req_0, ack => array_obj_ref_207_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_311_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_37_307, dout => array_obj_ref_311_resized_base_address, req => array_obj_ref_311_base_resize_req_0, ack => array_obj_ref_311_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_311_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_311_root_address, dout => iNsTr_38_312, req => array_obj_ref_311_final_reg_req_0, ack => array_obj_ref_311_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_388_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_52_384, dout => array_obj_ref_388_resized_base_address, req => array_obj_ref_388_base_resize_req_0, ack => array_obj_ref_388_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_388_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_388_root_address, dout => iNsTr_53_389, req => array_obj_ref_388_final_reg_req_0, ack => array_obj_ref_388_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_210_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_10_208, dout => ptr_deref_210_resized_base_address, req => ptr_deref_210_base_resize_req_0, ack => ptr_deref_210_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_315_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_38_312, dout => ptr_deref_315_resized_base_address, req => ptr_deref_315_base_resize_req_0, ack => ptr_deref_315_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_391_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_53_389, dout => ptr_deref_391_resized_base_address, req => ptr_deref_391_base_resize_req_0, ack => ptr_deref_391_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_255_inst: RegisterBase generic map(in_data_width => 8,out_data_width => 8) -- 
      port map( din => simple_obj_ref_254_wire, dout => iNsTr_22_256, req => type_cast_255_inst_req_0, ack => type_cast_255_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_267_inst: RegisterBase generic map(in_data_width => 8,out_data_width => 32) -- 
      port map( din => iNsTr_24_264, dout => iNsTr_25_268, req => type_cast_267_inst_req_0, ack => type_cast_267_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_328_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_42_325, dout => iNsTr_43_329, req => type_cast_328_inst_req_0, ack => type_cast_328_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_337_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_43_329, dout => type_cast_337_wire, req => type_cast_337_inst_req_0, ack => type_cast_337_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_347_inst: RegisterBase generic map(in_data_width => 8,out_data_width => 32) -- 
      port map( din => iNsTr_33_344, dout => iNsTr_34_348, req => type_cast_347_inst_req_0, ack => type_cast_347_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_368_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_367_wire, dout => iNsTr_48_369, req => type_cast_368_inst_req_0, ack => type_cast_368_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_372_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_48_369, dout => iNsTr_49_373, req => type_cast_372_inst_req_0, ack => type_cast_372_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_192_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      array_obj_ref_192_root_address_inst_ack_0 <= array_obj_ref_192_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_192_final_offset;
      array_obj_ref_192_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    array_obj_ref_201_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      array_obj_ref_201_root_address_inst_ack_0 <= array_obj_ref_201_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_201_final_offset;
      array_obj_ref_201_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    array_obj_ref_207_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      array_obj_ref_207_root_address_inst_ack_0 <= array_obj_ref_207_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_207_resized_base_address;
      array_obj_ref_207_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    array_obj_ref_311_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      array_obj_ref_311_root_address_inst_ack_0 <= array_obj_ref_311_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_311_resized_base_address;
      array_obj_ref_311_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    array_obj_ref_388_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      array_obj_ref_388_root_address_inst_ack_0 <= array_obj_ref_388_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_388_resized_base_address;
      array_obj_ref_388_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_156_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_156_gather_scatter_ack_0 <= ptr_deref_156_gather_scatter_req_0;
      aggregated_sig <= expr_157_wire_constant;
      ptr_deref_156_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_156_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_156_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_156_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_163_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_163_gather_scatter_ack_0 <= ptr_deref_163_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_163_data_0 & ptr_deref_163_data_1 & ptr_deref_163_data_2 & ptr_deref_163_data_3;
      iNsTr_2_164 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_183_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_183_gather_scatter_ack_0 <= ptr_deref_183_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_183_data_0 & ptr_deref_183_data_1 & ptr_deref_183_data_2 & ptr_deref_183_data_3;
      iNsTr_5_184 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_197_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_197_gather_scatter_ack_0 <= ptr_deref_197_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_197_data_0 & ptr_deref_197_data_1 & ptr_deref_197_data_2 & ptr_deref_197_data_3;
      iNsTr_8_198 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_210_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_210_gather_scatter_ack_0 <= ptr_deref_210_gather_scatter_req_0;
      aggregated_sig <= iNsTr_7_194;
      ptr_deref_210_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_210_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_210_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_210_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_210_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_210_root_address_inst_ack_0 <= ptr_deref_210_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_210_resized_base_address;
      ptr_deref_210_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_215_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_215_gather_scatter_ack_0 <= ptr_deref_215_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_215_data_0 & ptr_deref_215_data_1 & ptr_deref_215_data_2 & ptr_deref_215_data_3;
      iNsTr_12_216 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_223_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_223_gather_scatter_ack_0 <= ptr_deref_223_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_221;
      ptr_deref_223_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_223_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_223_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_223_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_235_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_235_gather_scatter_ack_0 <= ptr_deref_235_gather_scatter_req_0;
      aggregated_sig <= expr_236_wire_constant;
      ptr_deref_235_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_235_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_235_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_235_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_258_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_258_gather_scatter_ack_0 <= ptr_deref_258_gather_scatter_req_0;
      aggregated_sig <= iNsTr_22_256;
      ptr_deref_258_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_263_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_263_gather_scatter_ack_0 <= ptr_deref_263_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_263_data_0;
      iNsTr_24_264 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_285_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_285_gather_scatter_ack_0 <= ptr_deref_285_gather_scatter_req_0;
      aggregated_sig <= iNsTr_28_283;
      ptr_deref_285_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_285_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_285_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_285_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_315_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_315_gather_scatter_ack_0 <= ptr_deref_315_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_315_data_0 & ptr_deref_315_data_1 & ptr_deref_315_data_2 & ptr_deref_315_data_3;
      iNsTr_39_316 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_315_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_315_root_address_inst_ack_0 <= ptr_deref_315_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_315_resized_base_address;
      ptr_deref_315_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_324_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_324_gather_scatter_ack_0 <= ptr_deref_324_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_324_data_0 & ptr_deref_324_data_1 & ptr_deref_324_data_2 & ptr_deref_324_data_3;
      iNsTr_42_325 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_343_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_343_gather_scatter_ack_0 <= ptr_deref_343_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_343_data_0;
      iNsTr_33_344 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_375_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_375_gather_scatter_ack_0 <= ptr_deref_375_gather_scatter_req_0;
      aggregated_sig <= iNsTr_49_373;
      ptr_deref_375_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_375_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_375_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_375_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_383_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_383_gather_scatter_ack_0 <= ptr_deref_383_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_383_data_0 & ptr_deref_383_data_1 & ptr_deref_383_data_2 & ptr_deref_383_data_3;
      iNsTr_52_384 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_391_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_391_gather_scatter_ack_0 <= ptr_deref_391_gather_scatter_req_0;
      aggregated_sig <= iNsTr_51_380;
      ptr_deref_391_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_391_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_391_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_391_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_391_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_391_root_address_inst_ack_0 <= ptr_deref_391_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_391_resized_base_address;
      ptr_deref_391_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_396_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_396_gather_scatter_ack_0 <= ptr_deref_396_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_396_data_0 & ptr_deref_396_data_1 & ptr_deref_396_data_2 & ptr_deref_396_data_3;
      iNsTr_55_397 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_243_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_243_gather_scatter_ack_0 <= simple_obj_ref_243_gather_scatter_req_0;
      aggregated_sig <= iNsTr_18_242;
      simple_obj_ref_243_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_282_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_282_gather_scatter_ack_0 <= simple_obj_ref_282_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_282_data_0;
      iNsTr_28_283 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_289_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_289_gather_scatter_ack_0 <= simple_obj_ref_289_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_289_data_0;
      iNsTr_30_290 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_306_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_306_gather_scatter_ack_0 <= simple_obj_ref_306_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_306_data_0;
      iNsTr_37_307 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_317_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_317_gather_scatter_ack_0 <= simple_obj_ref_317_gather_scatter_req_0;
      aggregated_sig <= iNsTr_39_316;
      simple_obj_ref_317_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_379_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_379_gather_scatter_ack_0 <= simple_obj_ref_379_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_379_data_0;
      iNsTr_51_380 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_398_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_398_gather_scatter_ack_0 <= simple_obj_ref_398_gather_scatter_req_0;
      aggregated_sig <= iNsTr_55_397;
      simple_obj_ref_398_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_174_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_173;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_174_branch_req_0,
          ack0 => if_stmt_174_branch_ack_0,
          ack1 => if_stmt_174_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_274_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_26_273;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_274_branch_req_0,
          ack0 => if_stmt_274_branch_ack_0,
          ack1 => if_stmt_274_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_298_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_31_297;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_298_branch_req_0,
          ack0 => if_stmt_298_branch_ack_0,
          ack1 => if_stmt_298_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_354_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_35_353;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_354_branch_req_0,
          ack0 => if_stmt_354_branch_ack_0,
          ack1 => if_stmt_354_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_192_index_0_scale 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_191_resized;
      simple_obj_ref_191_scaled <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "001000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_192_index_0_scale_req_0,
          ackL => array_obj_ref_192_index_0_scale_ack_0,
          reqR => array_obj_ref_192_index_0_scale_req_1,
          ackR => array_obj_ref_192_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_201_index_0_scale 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_200_resized;
      simple_obj_ref_200_scaled <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "001000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_201_index_0_scale_req_0,
          ackL => array_obj_ref_201_index_0_scale_ack_0,
          reqR => array_obj_ref_201_index_0_scale_req_1,
          ackR => array_obj_ref_201_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_171_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_168_wire;
      iNsTr_3_173 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_171_inst_req_0,
          ackL => binary_171_inst_ack_0,
          reqR => binary_171_inst_req_1,
          ackR => binary_171_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_188_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_5_184;
      iNsTr_6_189 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_188_inst_req_0,
          ackL => binary_188_inst_ack_0,
          reqR => binary_188_inst_req_1,
          ackR => binary_188_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_220_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_216;
      iNsTr_13_221 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_220_inst_req_0,
          ackL => binary_220_inst_ack_0,
          reqR => binary_220_inst_req_1,
          ackR => binary_220_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_272_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_25_268;
      iNsTr_26_273 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_272_inst_req_0,
          ackL => binary_272_inst_ack_0,
          reqR => binary_272_inst_req_1,
          ackR => binary_272_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_296_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_293_wire;
      iNsTr_31_297 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_296_inst_req_0,
          ackL => binary_296_inst_ack_0,
          reqR => binary_296_inst_req_1,
          ackR => binary_296_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_352_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_34_348;
      iNsTr_35_353 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_352_inst_req_0,
          ackL => binary_352_inst_ack_0,
          reqR => binary_352_inst_req_1,
          ackR => binary_352_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : ptr_deref_210_addr_0 ptr_deref_315_addr_0 ptr_deref_391_addr_0 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(17 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_210_root_address & ptr_deref_315_root_address & ptr_deref_391_root_address;
      ptr_deref_210_word_address_0 <= data_out(17 downto 12);
      ptr_deref_315_word_address_0 <= data_out(11 downto 6);
      ptr_deref_391_word_address_0 <= data_out(5 downto 0);
      reqL(2) <= ptr_deref_210_addr_0_req_0;
      reqL(1) <= ptr_deref_315_addr_0_req_0;
      reqL(0) <= ptr_deref_391_addr_0_req_0;
      ptr_deref_210_addr_0_ack_0 <= ackL(2);
      ptr_deref_315_addr_0_ack_0 <= ackL(1);
      ptr_deref_391_addr_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_210_addr_0_req_1;
      reqR(1) <= ptr_deref_315_addr_0_req_1;
      reqR(0) <= ptr_deref_391_addr_0_req_1;
      ptr_deref_210_addr_0_ack_1 <= ackR(2);
      ptr_deref_315_addr_0_ack_1 <= ackR(1);
      ptr_deref_391_addr_0_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000000",
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true, 
          num_reqs => 3--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : ptr_deref_210_addr_1 ptr_deref_315_addr_1 ptr_deref_391_addr_1 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(17 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_210_root_address & ptr_deref_315_root_address & ptr_deref_391_root_address;
      ptr_deref_210_word_address_1 <= data_out(17 downto 12);
      ptr_deref_315_word_address_1 <= data_out(11 downto 6);
      ptr_deref_391_word_address_1 <= data_out(5 downto 0);
      reqL(2) <= ptr_deref_210_addr_1_req_0;
      reqL(1) <= ptr_deref_315_addr_1_req_0;
      reqL(0) <= ptr_deref_391_addr_1_req_0;
      ptr_deref_210_addr_1_ack_0 <= ackL(2);
      ptr_deref_315_addr_1_ack_0 <= ackL(1);
      ptr_deref_391_addr_1_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_210_addr_1_req_1;
      reqR(1) <= ptr_deref_315_addr_1_req_1;
      reqR(0) <= ptr_deref_391_addr_1_req_1;
      ptr_deref_210_addr_1_ack_1 <= ackR(2);
      ptr_deref_315_addr_1_ack_1 <= ackR(1);
      ptr_deref_391_addr_1_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000001",
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true, 
          num_reqs => 3--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : ptr_deref_391_addr_2 ptr_deref_210_addr_2 ptr_deref_315_addr_2 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(17 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_391_root_address & ptr_deref_210_root_address & ptr_deref_315_root_address;
      ptr_deref_391_word_address_2 <= data_out(17 downto 12);
      ptr_deref_210_word_address_2 <= data_out(11 downto 6);
      ptr_deref_315_word_address_2 <= data_out(5 downto 0);
      reqL(2) <= ptr_deref_391_addr_2_req_0;
      reqL(1) <= ptr_deref_210_addr_2_req_0;
      reqL(0) <= ptr_deref_315_addr_2_req_0;
      ptr_deref_391_addr_2_ack_0 <= ackL(2);
      ptr_deref_210_addr_2_ack_0 <= ackL(1);
      ptr_deref_315_addr_2_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_391_addr_2_req_1;
      reqR(1) <= ptr_deref_210_addr_2_req_1;
      reqR(0) <= ptr_deref_315_addr_2_req_1;
      ptr_deref_391_addr_2_ack_1 <= ackR(2);
      ptr_deref_210_addr_2_ack_1 <= ackR(1);
      ptr_deref_315_addr_2_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000010",
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true, 
          num_reqs => 3--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_315_addr_3 ptr_deref_210_addr_3 ptr_deref_391_addr_3 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(17 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_315_root_address & ptr_deref_210_root_address & ptr_deref_391_root_address;
      ptr_deref_315_word_address_3 <= data_out(17 downto 12);
      ptr_deref_210_word_address_3 <= data_out(11 downto 6);
      ptr_deref_391_word_address_3 <= data_out(5 downto 0);
      reqL(2) <= ptr_deref_315_addr_3_req_0;
      reqL(1) <= ptr_deref_210_addr_3_req_0;
      reqL(0) <= ptr_deref_391_addr_3_req_0;
      ptr_deref_315_addr_3_ack_0 <= ackL(2);
      ptr_deref_210_addr_3_ack_0 <= ackL(1);
      ptr_deref_391_addr_3_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_315_addr_3_req_1;
      reqR(1) <= ptr_deref_210_addr_3_req_1;
      reqR(0) <= ptr_deref_391_addr_3_req_1;
      ptr_deref_315_addr_3_ack_1 <= ackR(2);
      ptr_deref_210_addr_3_ack_1 <= ackR(1);
      ptr_deref_391_addr_3_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000011",
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true, 
          num_reqs => 3--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : type_cast_168_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_2_164;
      type_cast_168_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => type_cast_168_inst_req_0,
          ackL => type_cast_168_inst_ack_0,
          reqR => type_cast_168_inst_req_1,
          ackR => type_cast_168_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : type_cast_293_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_30_290;
      type_cast_293_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => type_cast_293_inst_req_0,
          ackL => type_cast_293_inst_ack_0,
          reqR => type_cast_293_inst_req_1,
          ackR => type_cast_293_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared load operator group (0) : ptr_deref_183_load_0 ptr_deref_263_load_0 ptr_deref_163_load_0 ptr_deref_324_load_0 ptr_deref_383_load_0 ptr_deref_315_load_0 ptr_deref_343_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(41 downto 0);
      signal data_out: std_logic_vector(55 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 6 downto 0);
      -- 
    begin -- 
      reqL(6) <= ptr_deref_183_load_0_req_0;
      reqL(5) <= ptr_deref_263_load_0_req_0;
      reqL(4) <= ptr_deref_163_load_0_req_0;
      reqL(3) <= ptr_deref_324_load_0_req_0;
      reqL(2) <= ptr_deref_383_load_0_req_0;
      reqL(1) <= ptr_deref_315_load_0_req_0;
      reqL(0) <= ptr_deref_343_load_0_req_0;
      ptr_deref_183_load_0_ack_0 <= ackL(6);
      ptr_deref_263_load_0_ack_0 <= ackL(5);
      ptr_deref_163_load_0_ack_0 <= ackL(4);
      ptr_deref_324_load_0_ack_0 <= ackL(3);
      ptr_deref_383_load_0_ack_0 <= ackL(2);
      ptr_deref_315_load_0_ack_0 <= ackL(1);
      ptr_deref_343_load_0_ack_0 <= ackL(0);
      reqR(6) <= ptr_deref_183_load_0_req_1;
      reqR(5) <= ptr_deref_263_load_0_req_1;
      reqR(4) <= ptr_deref_163_load_0_req_1;
      reqR(3) <= ptr_deref_324_load_0_req_1;
      reqR(2) <= ptr_deref_383_load_0_req_1;
      reqR(1) <= ptr_deref_315_load_0_req_1;
      reqR(0) <= ptr_deref_343_load_0_req_1;
      ptr_deref_183_load_0_ack_1 <= ackR(6);
      ptr_deref_263_load_0_ack_1 <= ackR(5);
      ptr_deref_163_load_0_ack_1 <= ackR(4);
      ptr_deref_324_load_0_ack_1 <= ackR(3);
      ptr_deref_383_load_0_ack_1 <= ackR(2);
      ptr_deref_315_load_0_ack_1 <= ackR(1);
      ptr_deref_343_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_183_word_address_0 & ptr_deref_263_word_address_0 & ptr_deref_163_word_address_0 & ptr_deref_324_word_address_0 & ptr_deref_383_word_address_0 & ptr_deref_315_word_address_0 & ptr_deref_343_word_address_0;
      ptr_deref_183_data_0 <= data_out(55 downto 48);
      ptr_deref_263_data_0 <= data_out(47 downto 40);
      ptr_deref_163_data_0 <= data_out(39 downto 32);
      ptr_deref_324_data_0 <= data_out(31 downto 24);
      ptr_deref_383_data_0 <= data_out(23 downto 16);
      ptr_deref_315_data_0 <= data_out(15 downto 8);
      ptr_deref_343_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 7,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(11),
          mack => memory_space_1_lr_ack(11),
          maddr => memory_space_1_lr_addr(71 downto 66),
          mtag => memory_space_1_lr_tag(35 downto 33),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 7,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(11),
          mack => memory_space_1_lc_ack(11),
          mdata => memory_space_1_lc_data(95 downto 88),
          mtag => memory_space_1_lc_tag(35 downto 33),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_183_load_1 ptr_deref_324_load_1 ptr_deref_315_load_1 ptr_deref_383_load_1 ptr_deref_163_load_1 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(39 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= ptr_deref_183_load_1_req_0;
      reqL(3) <= ptr_deref_324_load_1_req_0;
      reqL(2) <= ptr_deref_315_load_1_req_0;
      reqL(1) <= ptr_deref_383_load_1_req_0;
      reqL(0) <= ptr_deref_163_load_1_req_0;
      ptr_deref_183_load_1_ack_0 <= ackL(4);
      ptr_deref_324_load_1_ack_0 <= ackL(3);
      ptr_deref_315_load_1_ack_0 <= ackL(2);
      ptr_deref_383_load_1_ack_0 <= ackL(1);
      ptr_deref_163_load_1_ack_0 <= ackL(0);
      reqR(4) <= ptr_deref_183_load_1_req_1;
      reqR(3) <= ptr_deref_324_load_1_req_1;
      reqR(2) <= ptr_deref_315_load_1_req_1;
      reqR(1) <= ptr_deref_383_load_1_req_1;
      reqR(0) <= ptr_deref_163_load_1_req_1;
      ptr_deref_183_load_1_ack_1 <= ackR(4);
      ptr_deref_324_load_1_ack_1 <= ackR(3);
      ptr_deref_315_load_1_ack_1 <= ackR(2);
      ptr_deref_383_load_1_ack_1 <= ackR(1);
      ptr_deref_163_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_183_word_address_1 & ptr_deref_324_word_address_1 & ptr_deref_315_word_address_1 & ptr_deref_383_word_address_1 & ptr_deref_163_word_address_1;
      ptr_deref_183_data_1 <= data_out(39 downto 32);
      ptr_deref_324_data_1 <= data_out(31 downto 24);
      ptr_deref_315_data_1 <= data_out(23 downto 16);
      ptr_deref_383_data_1 <= data_out(15 downto 8);
      ptr_deref_163_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 5,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(10),
          mack => memory_space_1_lr_ack(10),
          maddr => memory_space_1_lr_addr(65 downto 60),
          mtag => memory_space_1_lr_tag(32 downto 30),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 5,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(10),
          mack => memory_space_1_lc_ack(10),
          mdata => memory_space_1_lc_data(87 downto 80),
          mtag => memory_space_1_lc_tag(32 downto 30),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_183_load_2 ptr_deref_315_load_2 ptr_deref_383_load_2 ptr_deref_324_load_2 ptr_deref_163_load_2 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(39 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= ptr_deref_183_load_2_req_0;
      reqL(3) <= ptr_deref_315_load_2_req_0;
      reqL(2) <= ptr_deref_383_load_2_req_0;
      reqL(1) <= ptr_deref_324_load_2_req_0;
      reqL(0) <= ptr_deref_163_load_2_req_0;
      ptr_deref_183_load_2_ack_0 <= ackL(4);
      ptr_deref_315_load_2_ack_0 <= ackL(3);
      ptr_deref_383_load_2_ack_0 <= ackL(2);
      ptr_deref_324_load_2_ack_0 <= ackL(1);
      ptr_deref_163_load_2_ack_0 <= ackL(0);
      reqR(4) <= ptr_deref_183_load_2_req_1;
      reqR(3) <= ptr_deref_315_load_2_req_1;
      reqR(2) <= ptr_deref_383_load_2_req_1;
      reqR(1) <= ptr_deref_324_load_2_req_1;
      reqR(0) <= ptr_deref_163_load_2_req_1;
      ptr_deref_183_load_2_ack_1 <= ackR(4);
      ptr_deref_315_load_2_ack_1 <= ackR(3);
      ptr_deref_383_load_2_ack_1 <= ackR(2);
      ptr_deref_324_load_2_ack_1 <= ackR(1);
      ptr_deref_163_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_183_word_address_2 & ptr_deref_315_word_address_2 & ptr_deref_383_word_address_2 & ptr_deref_324_word_address_2 & ptr_deref_163_word_address_2;
      ptr_deref_183_data_2 <= data_out(39 downto 32);
      ptr_deref_315_data_2 <= data_out(31 downto 24);
      ptr_deref_383_data_2 <= data_out(23 downto 16);
      ptr_deref_324_data_2 <= data_out(15 downto 8);
      ptr_deref_163_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 5,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(9),
          mack => memory_space_1_lr_ack(9),
          maddr => memory_space_1_lr_addr(59 downto 54),
          mtag => memory_space_1_lr_tag(29 downto 27),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 5,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(9),
          mack => memory_space_1_lc_ack(9),
          mdata => memory_space_1_lc_data(79 downto 72),
          mtag => memory_space_1_lc_tag(29 downto 27),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_183_load_3 ptr_deref_163_load_3 ptr_deref_315_load_3 ptr_deref_383_load_3 ptr_deref_324_load_3 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(39 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= ptr_deref_183_load_3_req_0;
      reqL(3) <= ptr_deref_163_load_3_req_0;
      reqL(2) <= ptr_deref_315_load_3_req_0;
      reqL(1) <= ptr_deref_383_load_3_req_0;
      reqL(0) <= ptr_deref_324_load_3_req_0;
      ptr_deref_183_load_3_ack_0 <= ackL(4);
      ptr_deref_163_load_3_ack_0 <= ackL(3);
      ptr_deref_315_load_3_ack_0 <= ackL(2);
      ptr_deref_383_load_3_ack_0 <= ackL(1);
      ptr_deref_324_load_3_ack_0 <= ackL(0);
      reqR(4) <= ptr_deref_183_load_3_req_1;
      reqR(3) <= ptr_deref_163_load_3_req_1;
      reqR(2) <= ptr_deref_315_load_3_req_1;
      reqR(1) <= ptr_deref_383_load_3_req_1;
      reqR(0) <= ptr_deref_324_load_3_req_1;
      ptr_deref_183_load_3_ack_1 <= ackR(4);
      ptr_deref_163_load_3_ack_1 <= ackR(3);
      ptr_deref_315_load_3_ack_1 <= ackR(2);
      ptr_deref_383_load_3_ack_1 <= ackR(1);
      ptr_deref_324_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_183_word_address_3 & ptr_deref_163_word_address_3 & ptr_deref_315_word_address_3 & ptr_deref_383_word_address_3 & ptr_deref_324_word_address_3;
      ptr_deref_183_data_3 <= data_out(39 downto 32);
      ptr_deref_163_data_3 <= data_out(31 downto 24);
      ptr_deref_315_data_3 <= data_out(23 downto 16);
      ptr_deref_383_data_3 <= data_out(15 downto 8);
      ptr_deref_324_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 5,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(8),
          mack => memory_space_1_lr_ack(8),
          maddr => memory_space_1_lr_addr(53 downto 48),
          mtag => memory_space_1_lr_tag(26 downto 24),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 5,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(8),
          mack => memory_space_1_lc_ack(8),
          mdata => memory_space_1_lc_data(71 downto 64),
          mtag => memory_space_1_lc_tag(26 downto 24),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_197_load_0 ptr_deref_396_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_197_load_0_req_0;
      reqL(0) <= ptr_deref_396_load_0_req_0;
      ptr_deref_197_load_0_ack_0 <= ackL(1);
      ptr_deref_396_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_197_load_0_req_1;
      reqR(0) <= ptr_deref_396_load_0_req_1;
      ptr_deref_197_load_0_ack_1 <= ackR(1);
      ptr_deref_396_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_197_word_address_0 & ptr_deref_396_word_address_0;
      ptr_deref_197_data_0 <= data_out(15 downto 8);
      ptr_deref_396_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(7),
          mack => memory_space_1_lr_ack(7),
          maddr => memory_space_1_lr_addr(47 downto 42),
          mtag => memory_space_1_lr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(7),
          mack => memory_space_1_lc_ack(7),
          mdata => memory_space_1_lc_data(63 downto 56),
          mtag => memory_space_1_lc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_197_load_1 ptr_deref_396_load_1 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_197_load_1_req_0;
      reqL(0) <= ptr_deref_396_load_1_req_0;
      ptr_deref_197_load_1_ack_0 <= ackL(1);
      ptr_deref_396_load_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_197_load_1_req_1;
      reqR(0) <= ptr_deref_396_load_1_req_1;
      ptr_deref_197_load_1_ack_1 <= ackR(1);
      ptr_deref_396_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_197_word_address_1 & ptr_deref_396_word_address_1;
      ptr_deref_197_data_1 <= data_out(15 downto 8);
      ptr_deref_396_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(6),
          mack => memory_space_1_lr_ack(6),
          maddr => memory_space_1_lr_addr(41 downto 36),
          mtag => memory_space_1_lr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(6),
          mack => memory_space_1_lc_ack(6),
          mdata => memory_space_1_lc_data(55 downto 48),
          mtag => memory_space_1_lc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_197_load_2 ptr_deref_396_load_2 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_197_load_2_req_0;
      reqL(0) <= ptr_deref_396_load_2_req_0;
      ptr_deref_197_load_2_ack_0 <= ackL(1);
      ptr_deref_396_load_2_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_197_load_2_req_1;
      reqR(0) <= ptr_deref_396_load_2_req_1;
      ptr_deref_197_load_2_ack_1 <= ackR(1);
      ptr_deref_396_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_197_word_address_2 & ptr_deref_396_word_address_2;
      ptr_deref_197_data_2 <= data_out(15 downto 8);
      ptr_deref_396_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(5),
          mack => memory_space_1_lr_ack(5),
          maddr => memory_space_1_lr_addr(35 downto 30),
          mtag => memory_space_1_lr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(5),
          mack => memory_space_1_lc_ack(5),
          mdata => memory_space_1_lc_data(47 downto 40),
          mtag => memory_space_1_lc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_197_load_3 ptr_deref_396_load_3 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_197_load_3_req_0;
      reqL(0) <= ptr_deref_396_load_3_req_0;
      ptr_deref_197_load_3_ack_0 <= ackL(1);
      ptr_deref_396_load_3_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_197_load_3_req_1;
      reqR(0) <= ptr_deref_396_load_3_req_1;
      ptr_deref_197_load_3_ack_1 <= ackR(1);
      ptr_deref_396_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_197_word_address_3 & ptr_deref_396_word_address_3;
      ptr_deref_197_data_3 <= data_out(15 downto 8);
      ptr_deref_396_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(4),
          mack => memory_space_1_lr_ack(4),
          maddr => memory_space_1_lr_addr(29 downto 24),
          mtag => memory_space_1_lr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(4),
          mack => memory_space_1_lc_ack(4),
          mdata => memory_space_1_lc_data(39 downto 32),
          mtag => memory_space_1_lc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared load operator group (8) : ptr_deref_215_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_215_load_0_req_0;
      ptr_deref_215_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_215_load_0_req_1;
      ptr_deref_215_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_215_word_address_0;
      ptr_deref_215_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(3),
          mack => memory_space_1_lr_ack(3),
          maddr => memory_space_1_lr_addr(23 downto 18),
          mtag => memory_space_1_lr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(3),
          mack => memory_space_1_lc_ack(3),
          mdata => memory_space_1_lc_data(31 downto 24),
          mtag => memory_space_1_lc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- shared load operator group (9) : ptr_deref_215_load_1 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_215_load_1_req_0;
      ptr_deref_215_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_215_load_1_req_1;
      ptr_deref_215_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_215_word_address_1;
      ptr_deref_215_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(2),
          mack => memory_space_1_lr_ack(2),
          maddr => memory_space_1_lr_addr(17 downto 12),
          mtag => memory_space_1_lr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(2),
          mack => memory_space_1_lc_ack(2),
          mdata => memory_space_1_lc_data(23 downto 16),
          mtag => memory_space_1_lc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    -- shared load operator group (10) : ptr_deref_215_load_2 
    LoadGroup10: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_215_load_2_req_0;
      ptr_deref_215_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_215_load_2_req_1;
      ptr_deref_215_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_215_word_address_2;
      ptr_deref_215_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(1),
          mack => memory_space_1_lr_ack(1),
          maddr => memory_space_1_lr_addr(11 downto 6),
          mtag => memory_space_1_lr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(1),
          mack => memory_space_1_lc_ack(1),
          mdata => memory_space_1_lc_data(15 downto 8),
          mtag => memory_space_1_lc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 10
    -- shared load operator group (11) : ptr_deref_215_load_3 
    LoadGroup11: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_215_load_3_req_0;
      ptr_deref_215_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_215_load_3_req_1;
      ptr_deref_215_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_215_word_address_3;
      ptr_deref_215_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(5 downto 0),
          mtag => memory_space_1_lr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 11
    -- shared load operator group (12) : simple_obj_ref_282_load_0 simple_obj_ref_306_load_0 simple_obj_ref_379_load_0 
    LoadGroup12: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= simple_obj_ref_282_load_0_req_0;
      reqL(1) <= simple_obj_ref_306_load_0_req_0;
      reqL(0) <= simple_obj_ref_379_load_0_req_0;
      simple_obj_ref_282_load_0_ack_0 <= ackL(2);
      simple_obj_ref_306_load_0_ack_0 <= ackL(1);
      simple_obj_ref_379_load_0_ack_0 <= ackL(0);
      reqR(2) <= simple_obj_ref_282_load_0_req_1;
      reqR(1) <= simple_obj_ref_306_load_0_req_1;
      reqR(0) <= simple_obj_ref_379_load_0_req_1;
      simple_obj_ref_282_load_0_ack_1 <= ackR(2);
      simple_obj_ref_306_load_0_ack_1 <= ackR(1);
      simple_obj_ref_379_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_282_word_address_0 & simple_obj_ref_306_word_address_0 & simple_obj_ref_379_word_address_0;
      simple_obj_ref_282_data_0 <= data_out(95 downto 64);
      simple_obj_ref_306_data_0 <= data_out(63 downto 32);
      simple_obj_ref_379_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 3,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(1),
          mack => memory_space_2_lr_ack(1),
          maddr => memory_space_2_lr_addr(1 downto 1),
          mtag => memory_space_2_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(1),
          mack => memory_space_2_lc_ack(1),
          mdata => memory_space_2_lc_data(63 downto 32),
          mtag => memory_space_2_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 12
    -- shared load operator group (13) : simple_obj_ref_289_load_0 
    LoadGroup13: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_289_load_0_req_0;
      simple_obj_ref_289_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_289_load_0_req_1;
      simple_obj_ref_289_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_289_word_address_0;
      simple_obj_ref_289_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 13
    -- shared store operator group (0) : ptr_deref_156_store_0 ptr_deref_258_store_0 ptr_deref_235_store_0 ptr_deref_210_store_0 ptr_deref_375_store_0 ptr_deref_285_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(35 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_156_store_0_req_0;
      reqL(4) <= ptr_deref_258_store_0_req_0;
      reqL(3) <= ptr_deref_235_store_0_req_0;
      reqL(2) <= ptr_deref_210_store_0_req_0;
      reqL(1) <= ptr_deref_375_store_0_req_0;
      reqL(0) <= ptr_deref_285_store_0_req_0;
      ptr_deref_156_store_0_ack_0 <= ackL(5);
      ptr_deref_258_store_0_ack_0 <= ackL(4);
      ptr_deref_235_store_0_ack_0 <= ackL(3);
      ptr_deref_210_store_0_ack_0 <= ackL(2);
      ptr_deref_375_store_0_ack_0 <= ackL(1);
      ptr_deref_285_store_0_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_156_store_0_req_1;
      reqR(4) <= ptr_deref_258_store_0_req_1;
      reqR(3) <= ptr_deref_235_store_0_req_1;
      reqR(2) <= ptr_deref_210_store_0_req_1;
      reqR(1) <= ptr_deref_375_store_0_req_1;
      reqR(0) <= ptr_deref_285_store_0_req_1;
      ptr_deref_156_store_0_ack_1 <= ackR(5);
      ptr_deref_258_store_0_ack_1 <= ackR(4);
      ptr_deref_235_store_0_ack_1 <= ackR(3);
      ptr_deref_210_store_0_ack_1 <= ackR(2);
      ptr_deref_375_store_0_ack_1 <= ackR(1);
      ptr_deref_285_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_156_word_address_0 & ptr_deref_258_word_address_0 & ptr_deref_235_word_address_0 & ptr_deref_210_word_address_0 & ptr_deref_375_word_address_0 & ptr_deref_285_word_address_0;
      data_in <= ptr_deref_156_data_0 & ptr_deref_258_data_0 & ptr_deref_235_data_0 & ptr_deref_210_data_0 & ptr_deref_375_data_0 & ptr_deref_285_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 6,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(7),
          mack => memory_space_1_sr_ack(7),
          maddr => memory_space_1_sr_addr(47 downto 42),
          mdata => memory_space_1_sr_data(63 downto 56),
          mtag => memory_space_1_sr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(7),
          mack => memory_space_1_sc_ack(7),
          mtag => memory_space_1_sc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_156_store_1 ptr_deref_235_store_1 ptr_deref_210_store_1 ptr_deref_375_store_1 ptr_deref_285_store_1 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(29 downto 0);
      signal data_in: std_logic_vector(39 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= ptr_deref_156_store_1_req_0;
      reqL(3) <= ptr_deref_235_store_1_req_0;
      reqL(2) <= ptr_deref_210_store_1_req_0;
      reqL(1) <= ptr_deref_375_store_1_req_0;
      reqL(0) <= ptr_deref_285_store_1_req_0;
      ptr_deref_156_store_1_ack_0 <= ackL(4);
      ptr_deref_235_store_1_ack_0 <= ackL(3);
      ptr_deref_210_store_1_ack_0 <= ackL(2);
      ptr_deref_375_store_1_ack_0 <= ackL(1);
      ptr_deref_285_store_1_ack_0 <= ackL(0);
      reqR(4) <= ptr_deref_156_store_1_req_1;
      reqR(3) <= ptr_deref_235_store_1_req_1;
      reqR(2) <= ptr_deref_210_store_1_req_1;
      reqR(1) <= ptr_deref_375_store_1_req_1;
      reqR(0) <= ptr_deref_285_store_1_req_1;
      ptr_deref_156_store_1_ack_1 <= ackR(4);
      ptr_deref_235_store_1_ack_1 <= ackR(3);
      ptr_deref_210_store_1_ack_1 <= ackR(2);
      ptr_deref_375_store_1_ack_1 <= ackR(1);
      ptr_deref_285_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_156_word_address_1 & ptr_deref_235_word_address_1 & ptr_deref_210_word_address_1 & ptr_deref_375_word_address_1 & ptr_deref_285_word_address_1;
      data_in <= ptr_deref_156_data_1 & ptr_deref_235_data_1 & ptr_deref_210_data_1 & ptr_deref_375_data_1 & ptr_deref_285_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 5,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(6),
          mack => memory_space_1_sr_ack(6),
          maddr => memory_space_1_sr_addr(41 downto 36),
          mdata => memory_space_1_sr_data(55 downto 48),
          mtag => memory_space_1_sr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 5,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(6),
          mack => memory_space_1_sc_ack(6),
          mtag => memory_space_1_sc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_156_store_2 ptr_deref_210_store_2 ptr_deref_235_store_2 ptr_deref_285_store_2 ptr_deref_375_store_2 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(29 downto 0);
      signal data_in: std_logic_vector(39 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= ptr_deref_156_store_2_req_0;
      reqL(3) <= ptr_deref_210_store_2_req_0;
      reqL(2) <= ptr_deref_235_store_2_req_0;
      reqL(1) <= ptr_deref_285_store_2_req_0;
      reqL(0) <= ptr_deref_375_store_2_req_0;
      ptr_deref_156_store_2_ack_0 <= ackL(4);
      ptr_deref_210_store_2_ack_0 <= ackL(3);
      ptr_deref_235_store_2_ack_0 <= ackL(2);
      ptr_deref_285_store_2_ack_0 <= ackL(1);
      ptr_deref_375_store_2_ack_0 <= ackL(0);
      reqR(4) <= ptr_deref_156_store_2_req_1;
      reqR(3) <= ptr_deref_210_store_2_req_1;
      reqR(2) <= ptr_deref_235_store_2_req_1;
      reqR(1) <= ptr_deref_285_store_2_req_1;
      reqR(0) <= ptr_deref_375_store_2_req_1;
      ptr_deref_156_store_2_ack_1 <= ackR(4);
      ptr_deref_210_store_2_ack_1 <= ackR(3);
      ptr_deref_235_store_2_ack_1 <= ackR(2);
      ptr_deref_285_store_2_ack_1 <= ackR(1);
      ptr_deref_375_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_156_word_address_2 & ptr_deref_210_word_address_2 & ptr_deref_235_word_address_2 & ptr_deref_285_word_address_2 & ptr_deref_375_word_address_2;
      data_in <= ptr_deref_156_data_2 & ptr_deref_210_data_2 & ptr_deref_235_data_2 & ptr_deref_285_data_2 & ptr_deref_375_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 5,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(5),
          mack => memory_space_1_sr_ack(5),
          maddr => memory_space_1_sr_addr(35 downto 30),
          mdata => memory_space_1_sr_data(47 downto 40),
          mtag => memory_space_1_sr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 5,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(5),
          mack => memory_space_1_sc_ack(5),
          mtag => memory_space_1_sc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_156_store_3 ptr_deref_210_store_3 ptr_deref_235_store_3 ptr_deref_375_store_3 ptr_deref_285_store_3 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(29 downto 0);
      signal data_in: std_logic_vector(39 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= ptr_deref_156_store_3_req_0;
      reqL(3) <= ptr_deref_210_store_3_req_0;
      reqL(2) <= ptr_deref_235_store_3_req_0;
      reqL(1) <= ptr_deref_375_store_3_req_0;
      reqL(0) <= ptr_deref_285_store_3_req_0;
      ptr_deref_156_store_3_ack_0 <= ackL(4);
      ptr_deref_210_store_3_ack_0 <= ackL(3);
      ptr_deref_235_store_3_ack_0 <= ackL(2);
      ptr_deref_375_store_3_ack_0 <= ackL(1);
      ptr_deref_285_store_3_ack_0 <= ackL(0);
      reqR(4) <= ptr_deref_156_store_3_req_1;
      reqR(3) <= ptr_deref_210_store_3_req_1;
      reqR(2) <= ptr_deref_235_store_3_req_1;
      reqR(1) <= ptr_deref_375_store_3_req_1;
      reqR(0) <= ptr_deref_285_store_3_req_1;
      ptr_deref_156_store_3_ack_1 <= ackR(4);
      ptr_deref_210_store_3_ack_1 <= ackR(3);
      ptr_deref_235_store_3_ack_1 <= ackR(2);
      ptr_deref_375_store_3_ack_1 <= ackR(1);
      ptr_deref_285_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_156_word_address_3 & ptr_deref_210_word_address_3 & ptr_deref_235_word_address_3 & ptr_deref_375_word_address_3 & ptr_deref_285_word_address_3;
      data_in <= ptr_deref_156_data_3 & ptr_deref_210_data_3 & ptr_deref_235_data_3 & ptr_deref_375_data_3 & ptr_deref_285_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 5,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(4),
          mack => memory_space_1_sr_ack(4),
          maddr => memory_space_1_sr_addr(29 downto 24),
          mdata => memory_space_1_sr_data(39 downto 32),
          mtag => memory_space_1_sr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 5,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(4),
          mack => memory_space_1_sc_ack(4),
          mtag => memory_space_1_sc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_223_store_0 ptr_deref_391_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_223_store_0_req_0;
      reqL(0) <= ptr_deref_391_store_0_req_0;
      ptr_deref_223_store_0_ack_0 <= ackL(1);
      ptr_deref_391_store_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_223_store_0_req_1;
      reqR(0) <= ptr_deref_391_store_0_req_1;
      ptr_deref_223_store_0_ack_1 <= ackR(1);
      ptr_deref_391_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_223_word_address_0 & ptr_deref_391_word_address_0;
      data_in <= ptr_deref_223_data_0 & ptr_deref_391_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(3),
          mack => memory_space_1_sr_ack(3),
          maddr => memory_space_1_sr_addr(23 downto 18),
          mdata => memory_space_1_sr_data(31 downto 24),
          mtag => memory_space_1_sr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(3),
          mack => memory_space_1_sc_ack(3),
          mtag => memory_space_1_sc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_223_store_1 ptr_deref_391_store_1 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_223_store_1_req_0;
      reqL(0) <= ptr_deref_391_store_1_req_0;
      ptr_deref_223_store_1_ack_0 <= ackL(1);
      ptr_deref_391_store_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_223_store_1_req_1;
      reqR(0) <= ptr_deref_391_store_1_req_1;
      ptr_deref_223_store_1_ack_1 <= ackR(1);
      ptr_deref_391_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_223_word_address_1 & ptr_deref_391_word_address_1;
      data_in <= ptr_deref_223_data_1 & ptr_deref_391_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(2),
          mack => memory_space_1_sr_ack(2),
          maddr => memory_space_1_sr_addr(17 downto 12),
          mdata => memory_space_1_sr_data(23 downto 16),
          mtag => memory_space_1_sr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(2),
          mack => memory_space_1_sc_ack(2),
          mtag => memory_space_1_sc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_223_store_2 ptr_deref_391_store_2 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_223_store_2_req_0;
      reqL(0) <= ptr_deref_391_store_2_req_0;
      ptr_deref_223_store_2_ack_0 <= ackL(1);
      ptr_deref_391_store_2_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_223_store_2_req_1;
      reqR(0) <= ptr_deref_391_store_2_req_1;
      ptr_deref_223_store_2_ack_1 <= ackR(1);
      ptr_deref_391_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_223_word_address_2 & ptr_deref_391_word_address_2;
      data_in <= ptr_deref_223_data_2 & ptr_deref_391_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(1),
          mack => memory_space_1_sr_ack(1),
          maddr => memory_space_1_sr_addr(11 downto 6),
          mdata => memory_space_1_sr_data(15 downto 8),
          mtag => memory_space_1_sr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(1),
          mack => memory_space_1_sc_ack(1),
          mtag => memory_space_1_sc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_223_store_3 ptr_deref_391_store_3 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_223_store_3_req_0;
      reqL(0) <= ptr_deref_391_store_3_req_0;
      ptr_deref_223_store_3_ack_0 <= ackL(1);
      ptr_deref_391_store_3_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_223_store_3_req_1;
      reqR(0) <= ptr_deref_391_store_3_req_1;
      ptr_deref_223_store_3_ack_1 <= ackR(1);
      ptr_deref_391_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_223_word_address_3 & ptr_deref_391_word_address_3;
      data_in <= ptr_deref_223_data_3 & ptr_deref_391_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(5 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared store operator group (8) : simple_obj_ref_243_store_0 simple_obj_ref_317_store_0 simple_obj_ref_398_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= simple_obj_ref_243_store_0_req_0;
      reqL(1) <= simple_obj_ref_317_store_0_req_0;
      reqL(0) <= simple_obj_ref_398_store_0_req_0;
      simple_obj_ref_243_store_0_ack_0 <= ackL(2);
      simple_obj_ref_317_store_0_ack_0 <= ackL(1);
      simple_obj_ref_398_store_0_ack_0 <= ackL(0);
      reqR(2) <= simple_obj_ref_243_store_0_req_1;
      reqR(1) <= simple_obj_ref_317_store_0_req_1;
      reqR(0) <= simple_obj_ref_398_store_0_req_1;
      simple_obj_ref_243_store_0_ack_1 <= ackR(2);
      simple_obj_ref_317_store_0_ack_1 <= ackR(1);
      simple_obj_ref_398_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_243_word_address_0 & simple_obj_ref_317_word_address_0 & simple_obj_ref_398_word_address_0;
      data_in <= simple_obj_ref_243_data_0 & simple_obj_ref_317_data_0 & simple_obj_ref_398_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    -- shared inport operator group (0) : simple_obj_ref_254_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_254_inst_req_0;
      simple_obj_ref_254_inst_ack_0 <= ack(0);
      simple_obj_ref_254_wire <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_request_pipe_read_req(0),
          oack => free_queue_request_pipe_read_ack(0),
          odata => free_queue_request_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_367_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_367_inst_req_0;
      simple_obj_ref_367_inst_ack_0 <= ack(0);
      simple_obj_ref_367_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_put_pipe_read_req(0),
          oack => free_queue_put_pipe_read_ack(0),
          odata => free_queue_put_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_335_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_335_inst_req_0;
      simple_obj_ref_335_inst_ack_0 <= ack(0);
      data_in <= type_cast_337_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_get_pipe_write_req(0),
          oack => free_queue_get_pipe_write_ack(0),
          odata => free_queue_get_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity input_module is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(11 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(11 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(71 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(35 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(11 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(11 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(95 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(35 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(47 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(23 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(7 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(23 downto 0);
    free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_data_pipe_read_data : in   std_logic_vector(31 downto 0);
    foo_in_pipe_write_req : out  std_logic_vector(0 downto 0);
    foo_in_pipe_write_ack : in   std_logic_vector(0 downto 0);
    foo_in_pipe_write_data : out  std_logic_vector(31 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity input_module;
architecture Default of input_module is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_494_load_0_req_1 : boolean;
  signal ptr_deref_494_load_2_req_1 : boolean;
  signal simple_obj_ref_505_inst_ack_0 : boolean;
  signal simple_obj_ref_505_inst_req_0 : boolean;
  signal ptr_deref_494_load_0_ack_1 : boolean;
  signal type_cast_507_inst_req_0 : boolean;
  signal ptr_deref_494_load_1_ack_1 : boolean;
  signal ptr_deref_494_load_1_req_1 : boolean;
  signal ptr_deref_494_load_2_ack_1 : boolean;
  signal type_cast_507_inst_ack_0 : boolean;
  signal ptr_deref_494_load_3_req_1 : boolean;
  signal type_cast_498_inst_req_0 : boolean;
  signal ptr_deref_494_load_3_ack_1 : boolean;
  signal type_cast_498_inst_ack_0 : boolean;
  signal ptr_deref_494_gather_scatter_req_0 : boolean;
  signal ptr_deref_494_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_423_inst_req_0 : boolean;
  signal simple_obj_ref_423_inst_ack_0 : boolean;
  signal simple_obj_ref_433_inst_req_0 : boolean;
  signal simple_obj_ref_433_inst_ack_0 : boolean;
  signal type_cast_434_inst_req_0 : boolean;
  signal type_cast_434_inst_ack_0 : boolean;
  signal type_cast_438_inst_req_0 : boolean;
  signal type_cast_438_inst_ack_0 : boolean;
  signal ptr_deref_441_gather_scatter_req_0 : boolean;
  signal ptr_deref_441_gather_scatter_ack_0 : boolean;
  signal ptr_deref_441_store_0_req_0 : boolean;
  signal ptr_deref_441_store_0_ack_0 : boolean;
  signal ptr_deref_441_store_1_req_0 : boolean;
  signal ptr_deref_441_store_1_ack_0 : boolean;
  signal ptr_deref_441_store_2_req_0 : boolean;
  signal ptr_deref_441_store_2_ack_0 : boolean;
  signal ptr_deref_441_store_3_req_0 : boolean;
  signal ptr_deref_441_store_3_ack_0 : boolean;
  signal ptr_deref_441_store_0_req_1 : boolean;
  signal ptr_deref_441_store_0_ack_1 : boolean;
  signal ptr_deref_441_store_1_req_1 : boolean;
  signal ptr_deref_441_store_1_ack_1 : boolean;
  signal ptr_deref_441_store_2_req_1 : boolean;
  signal ptr_deref_441_store_2_ack_1 : boolean;
  signal ptr_deref_441_store_3_req_1 : boolean;
  signal ptr_deref_441_store_3_ack_1 : boolean;
  signal ptr_deref_446_load_0_req_0 : boolean;
  signal ptr_deref_446_load_0_ack_0 : boolean;
  signal ptr_deref_446_load_1_req_0 : boolean;
  signal ptr_deref_446_load_1_ack_0 : boolean;
  signal ptr_deref_446_load_2_req_0 : boolean;
  signal ptr_deref_446_load_2_ack_0 : boolean;
  signal ptr_deref_446_load_3_req_0 : boolean;
  signal ptr_deref_446_load_3_ack_0 : boolean;
  signal ptr_deref_446_load_0_req_1 : boolean;
  signal ptr_deref_446_load_0_ack_1 : boolean;
  signal ptr_deref_446_load_1_req_1 : boolean;
  signal ptr_deref_446_load_1_ack_1 : boolean;
  signal ptr_deref_446_load_2_req_1 : boolean;
  signal ptr_deref_446_load_2_ack_1 : boolean;
  signal ptr_deref_446_load_3_req_1 : boolean;
  signal ptr_deref_446_load_3_ack_1 : boolean;
  signal ptr_deref_446_gather_scatter_req_0 : boolean;
  signal ptr_deref_446_gather_scatter_ack_0 : boolean;
  signal type_cast_450_inst_req_0 : boolean;
  signal type_cast_450_inst_ack_0 : boolean;
  signal type_cast_450_inst_req_1 : boolean;
  signal type_cast_450_inst_ack_1 : boolean;
  signal binary_453_inst_req_0 : boolean;
  signal binary_453_inst_ack_0 : boolean;
  signal binary_453_inst_req_1 : boolean;
  signal binary_453_inst_ack_1 : boolean;
  signal if_stmt_455_branch_req_0 : boolean;
  signal if_stmt_455_branch_ack_1 : boolean;
  signal if_stmt_455_branch_ack_0 : boolean;
  signal simple_obj_ref_468_inst_req_0 : boolean;
  signal simple_obj_ref_468_inst_ack_0 : boolean;
  signal type_cast_469_inst_req_0 : boolean;
  signal type_cast_469_inst_ack_0 : boolean;
  signal ptr_deref_472_gather_scatter_req_0 : boolean;
  signal ptr_deref_472_gather_scatter_ack_0 : boolean;
  signal ptr_deref_472_store_0_req_0 : boolean;
  signal ptr_deref_472_store_0_ack_0 : boolean;
  signal ptr_deref_472_store_1_req_0 : boolean;
  signal ptr_deref_472_store_1_ack_0 : boolean;
  signal ptr_deref_472_store_2_req_0 : boolean;
  signal ptr_deref_472_store_2_ack_0 : boolean;
  signal ptr_deref_472_store_3_req_0 : boolean;
  signal ptr_deref_472_store_3_ack_0 : boolean;
  signal ptr_deref_472_store_0_req_1 : boolean;
  signal ptr_deref_472_store_0_ack_1 : boolean;
  signal ptr_deref_472_store_1_req_1 : boolean;
  signal ptr_deref_472_store_1_ack_1 : boolean;
  signal ptr_deref_472_store_2_req_1 : boolean;
  signal ptr_deref_472_store_2_ack_1 : boolean;
  signal ptr_deref_472_store_3_req_1 : boolean;
  signal ptr_deref_472_store_3_ack_1 : boolean;
  signal ptr_deref_477_load_0_req_0 : boolean;
  signal ptr_deref_477_load_0_ack_0 : boolean;
  signal ptr_deref_477_load_1_req_0 : boolean;
  signal ptr_deref_477_load_1_ack_0 : boolean;
  signal ptr_deref_477_load_2_req_0 : boolean;
  signal ptr_deref_477_load_2_ack_0 : boolean;
  signal ptr_deref_477_load_3_req_0 : boolean;
  signal ptr_deref_477_load_3_ack_0 : boolean;
  signal ptr_deref_477_load_0_req_1 : boolean;
  signal ptr_deref_477_load_0_ack_1 : boolean;
  signal ptr_deref_477_load_1_req_1 : boolean;
  signal ptr_deref_477_load_1_ack_1 : boolean;
  signal ptr_deref_477_load_2_req_1 : boolean;
  signal ptr_deref_477_load_2_ack_1 : boolean;
  signal ptr_deref_477_load_3_req_1 : boolean;
  signal ptr_deref_477_load_3_ack_1 : boolean;
  signal ptr_deref_477_gather_scatter_req_0 : boolean;
  signal ptr_deref_477_gather_scatter_ack_0 : boolean;
  signal ptr_deref_481_load_0_req_0 : boolean;
  signal ptr_deref_481_load_0_ack_0 : boolean;
  signal ptr_deref_481_load_1_req_0 : boolean;
  signal ptr_deref_481_load_1_ack_0 : boolean;
  signal ptr_deref_481_load_2_req_0 : boolean;
  signal ptr_deref_481_load_2_ack_0 : boolean;
  signal ptr_deref_481_load_3_req_0 : boolean;
  signal ptr_deref_481_load_3_ack_0 : boolean;
  signal ptr_deref_481_load_0_req_1 : boolean;
  signal ptr_deref_481_load_0_ack_1 : boolean;
  signal ptr_deref_481_load_1_req_1 : boolean;
  signal ptr_deref_481_load_1_ack_1 : boolean;
  signal ptr_deref_481_load_2_req_1 : boolean;
  signal ptr_deref_481_load_2_ack_1 : boolean;
  signal ptr_deref_481_load_3_req_1 : boolean;
  signal ptr_deref_481_load_3_ack_1 : boolean;
  signal ptr_deref_481_gather_scatter_req_0 : boolean;
  signal ptr_deref_481_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_486_base_resize_req_0 : boolean;
  signal array_obj_ref_486_base_resize_ack_0 : boolean;
  signal array_obj_ref_486_root_address_inst_req_0 : boolean;
  signal array_obj_ref_486_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_486_root_address_inst_req_1 : boolean;
  signal array_obj_ref_486_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_486_final_reg_req_0 : boolean;
  signal array_obj_ref_486_final_reg_ack_0 : boolean;
  signal ptr_deref_489_base_resize_req_0 : boolean;
  signal ptr_deref_489_base_resize_ack_0 : boolean;
  signal ptr_deref_489_root_address_inst_req_0 : boolean;
  signal ptr_deref_489_root_address_inst_ack_0 : boolean;
  signal ptr_deref_489_addr_0_req_0 : boolean;
  signal ptr_deref_489_addr_0_ack_0 : boolean;
  signal ptr_deref_489_addr_0_req_1 : boolean;
  signal ptr_deref_489_addr_0_ack_1 : boolean;
  signal ptr_deref_489_addr_1_req_0 : boolean;
  signal ptr_deref_489_addr_1_ack_0 : boolean;
  signal ptr_deref_489_addr_1_req_1 : boolean;
  signal ptr_deref_489_addr_1_ack_1 : boolean;
  signal ptr_deref_489_addr_2_req_0 : boolean;
  signal ptr_deref_489_addr_2_ack_0 : boolean;
  signal ptr_deref_489_addr_2_req_1 : boolean;
  signal ptr_deref_489_addr_2_ack_1 : boolean;
  signal ptr_deref_489_addr_3_req_0 : boolean;
  signal ptr_deref_489_addr_3_ack_0 : boolean;
  signal ptr_deref_489_addr_3_req_1 : boolean;
  signal ptr_deref_489_addr_3_ack_1 : boolean;
  signal ptr_deref_489_gather_scatter_req_0 : boolean;
  signal ptr_deref_489_gather_scatter_ack_0 : boolean;
  signal ptr_deref_489_store_0_req_0 : boolean;
  signal ptr_deref_489_store_0_ack_0 : boolean;
  signal ptr_deref_489_store_1_req_0 : boolean;
  signal ptr_deref_489_store_1_ack_0 : boolean;
  signal ptr_deref_489_store_2_req_0 : boolean;
  signal ptr_deref_489_store_2_ack_0 : boolean;
  signal ptr_deref_489_store_3_req_0 : boolean;
  signal ptr_deref_489_store_3_ack_0 : boolean;
  signal ptr_deref_489_store_0_req_1 : boolean;
  signal ptr_deref_489_store_0_ack_1 : boolean;
  signal ptr_deref_489_store_1_req_1 : boolean;
  signal ptr_deref_489_store_1_ack_1 : boolean;
  signal ptr_deref_489_store_2_req_1 : boolean;
  signal ptr_deref_489_store_2_ack_1 : boolean;
  signal ptr_deref_489_store_3_req_1 : boolean;
  signal ptr_deref_489_store_3_ack_1 : boolean;
  signal ptr_deref_494_load_0_req_0 : boolean;
  signal ptr_deref_494_load_0_ack_0 : boolean;
  signal ptr_deref_494_load_1_req_0 : boolean;
  signal ptr_deref_494_load_1_ack_0 : boolean;
  signal ptr_deref_494_load_2_req_0 : boolean;
  signal ptr_deref_494_load_2_ack_0 : boolean;
  signal ptr_deref_494_load_3_req_0 : boolean;
  signal ptr_deref_494_load_3_ack_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  input_module_CP_2574: Block -- control-path 
    signal input_module_CP_2574_start: Boolean;
    signal Xentry_2575_symbol: Boolean;
    signal Xexit_2576_symbol: Boolean;
    signal branch_block_stmt_405_2577_symbol : Boolean;
    -- 
  begin -- 
    input_module_CP_2574_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_2575_symbol  <= input_module_CP_2574_start; -- transition $entry
    branch_block_stmt_405_2577: Block -- branch_block_stmt_405 
      signal branch_block_stmt_405_2577_start: Boolean;
      signal Xentry_2578_symbol: Boolean;
      signal Xexit_2579_symbol: Boolean;
      signal branch_block_stmt_405_x_xentry_x_xx_x2580_symbol : Boolean;
      signal branch_block_stmt_405_x_xexit_x_xx_x2581_symbol : Boolean;
      signal assign_stmt_411_to_assign_stmt_415_x_xentry_x_xx_x2582_symbol : Boolean;
      signal assign_stmt_411_to_assign_stmt_415_x_xexit_x_xx_x2583_symbol : Boolean;
      signal bb_0_bb_1_2584_symbol : Boolean;
      signal merge_stmt_417_x_xexit_x_xx_x2585_symbol : Boolean;
      signal assign_stmt_422_x_xentry_x_xx_x2586_symbol : Boolean;
      signal assign_stmt_422_x_xexit_x_xx_x2587_symbol : Boolean;
      signal assign_stmt_426_x_xentry_x_xx_x2588_symbol : Boolean;
      signal assign_stmt_426_x_xexit_x_xx_x2589_symbol : Boolean;
      signal assign_stmt_431_x_xentry_x_xx_x2590_symbol : Boolean;
      signal assign_stmt_431_x_xexit_x_xx_x2591_symbol : Boolean;
      signal assign_stmt_435_x_xentry_x_xx_x2592_symbol : Boolean;
      signal assign_stmt_435_x_xexit_x_xx_x2593_symbol : Boolean;
      signal assign_stmt_439_to_assign_stmt_454_x_xentry_x_xx_x2594_symbol : Boolean;
      signal assign_stmt_439_to_assign_stmt_454_x_xexit_x_xx_x2595_symbol : Boolean;
      signal if_stmt_455_x_xentry_x_xx_x2596_symbol : Boolean;
      signal if_stmt_455_x_xexit_x_xx_x2597_symbol : Boolean;
      signal merge_stmt_461_x_xentry_x_xx_x2598_symbol : Boolean;
      signal merge_stmt_461_x_xexit_x_xx_x2599_symbol : Boolean;
      signal assign_stmt_466_x_xentry_x_xx_x2600_symbol : Boolean;
      signal assign_stmt_466_x_xexit_x_xx_x2601_symbol : Boolean;
      signal assign_stmt_470_x_xentry_x_xx_x2602_symbol : Boolean;
      signal assign_stmt_470_x_xexit_x_xx_x2603_symbol : Boolean;
      signal assign_stmt_474_to_assign_stmt_504_x_xentry_x_xx_x2604_symbol : Boolean;
      signal assign_stmt_474_to_assign_stmt_504_x_xexit_x_xx_x2605_symbol : Boolean;
      signal assign_stmt_508_x_xentry_x_xx_x2606_symbol : Boolean;
      signal assign_stmt_508_x_xexit_x_xx_x2607_symbol : Boolean;
      signal bb_2_bb_1_2608_symbol : Boolean;
      signal assign_stmt_411_to_assign_stmt_415_2609_symbol : Boolean;
      signal assign_stmt_422_2612_symbol : Boolean;
      signal assign_stmt_426_2615_symbol : Boolean;
      signal assign_stmt_431_2626_symbol : Boolean;
      signal assign_stmt_435_2629_symbol : Boolean;
      signal assign_stmt_439_to_assign_stmt_454_2647_symbol : Boolean;
      signal if_stmt_455_dead_link_2804_symbol : Boolean;
      signal if_stmt_455_eval_test_2808_symbol : Boolean;
      signal simple_obj_ref_456_place_2812_symbol : Boolean;
      signal if_stmt_455_if_link_2813_symbol : Boolean;
      signal if_stmt_455_else_link_2817_symbol : Boolean;
      signal bb_1_bb_2_2821_symbol : Boolean;
      signal bb_1_bb_1_2822_symbol : Boolean;
      signal assign_stmt_466_2823_symbol : Boolean;
      signal assign_stmt_470_2826_symbol : Boolean;
      signal assign_stmt_474_to_assign_stmt_504_2844_symbol : Boolean;
      signal assign_stmt_508_3232_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_3251_symbol : Boolean;
      signal bb_1_bb_1_PhiReq_3254_symbol : Boolean;
      signal bb_2_bb_1_PhiReq_3257_symbol : Boolean;
      signal merge_stmt_417_PhiReqMerge_3260_symbol : Boolean;
      signal merge_stmt_417_PhiAck_3261_symbol : Boolean;
      signal merge_stmt_461_dead_link_3265_symbol : Boolean;
      signal bb_1_bb_2_PhiReq_3269_symbol : Boolean;
      signal merge_stmt_461_PhiReqMerge_3272_symbol : Boolean;
      signal merge_stmt_461_PhiAck_3273_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_405_2577_start <= Xentry_2575_symbol; -- control passed to block
      Xentry_2578_symbol  <= branch_block_stmt_405_2577_start; -- transition branch_block_stmt_405/$entry
      branch_block_stmt_405_x_xentry_x_xx_x2580_symbol  <=  Xentry_2578_symbol; -- place branch_block_stmt_405/branch_block_stmt_405__entry__ (optimized away) 
      branch_block_stmt_405_x_xexit_x_xx_x2581_symbol  <=   false ; -- place branch_block_stmt_405/branch_block_stmt_405__exit__ (optimized away) 
      assign_stmt_411_to_assign_stmt_415_x_xentry_x_xx_x2582_symbol  <=  branch_block_stmt_405_x_xentry_x_xx_x2580_symbol; -- place branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415__entry__ (optimized away) 
      assign_stmt_411_to_assign_stmt_415_x_xexit_x_xx_x2583_symbol  <=  assign_stmt_411_to_assign_stmt_415_2609_symbol; -- place branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415__exit__ (optimized away) 
      bb_0_bb_1_2584_symbol  <=  assign_stmt_411_to_assign_stmt_415_x_xexit_x_xx_x2583_symbol; -- place branch_block_stmt_405/bb_0_bb_1 (optimized away) 
      merge_stmt_417_x_xexit_x_xx_x2585_symbol  <=  merge_stmt_417_PhiAck_3261_symbol; -- place branch_block_stmt_405/merge_stmt_417__exit__ (optimized away) 
      assign_stmt_422_x_xentry_x_xx_x2586_symbol  <=  merge_stmt_417_x_xexit_x_xx_x2585_symbol; -- place branch_block_stmt_405/assign_stmt_422__entry__ (optimized away) 
      assign_stmt_422_x_xexit_x_xx_x2587_symbol  <=  assign_stmt_422_2612_symbol; -- place branch_block_stmt_405/assign_stmt_422__exit__ (optimized away) 
      assign_stmt_426_x_xentry_x_xx_x2588_symbol  <=  assign_stmt_422_x_xexit_x_xx_x2587_symbol; -- place branch_block_stmt_405/assign_stmt_426__entry__ (optimized away) 
      assign_stmt_426_x_xexit_x_xx_x2589_symbol  <=  assign_stmt_426_2615_symbol; -- place branch_block_stmt_405/assign_stmt_426__exit__ (optimized away) 
      assign_stmt_431_x_xentry_x_xx_x2590_symbol  <=  assign_stmt_426_x_xexit_x_xx_x2589_symbol; -- place branch_block_stmt_405/assign_stmt_431__entry__ (optimized away) 
      assign_stmt_431_x_xexit_x_xx_x2591_symbol  <=  assign_stmt_431_2626_symbol; -- place branch_block_stmt_405/assign_stmt_431__exit__ (optimized away) 
      assign_stmt_435_x_xentry_x_xx_x2592_symbol  <=  assign_stmt_431_x_xexit_x_xx_x2591_symbol; -- place branch_block_stmt_405/assign_stmt_435__entry__ (optimized away) 
      assign_stmt_435_x_xexit_x_xx_x2593_symbol  <=  assign_stmt_435_2629_symbol; -- place branch_block_stmt_405/assign_stmt_435__exit__ (optimized away) 
      assign_stmt_439_to_assign_stmt_454_x_xentry_x_xx_x2594_symbol  <=  assign_stmt_435_x_xexit_x_xx_x2593_symbol; -- place branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454__entry__ (optimized away) 
      assign_stmt_439_to_assign_stmt_454_x_xexit_x_xx_x2595_symbol  <=  assign_stmt_439_to_assign_stmt_454_2647_symbol; -- place branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454__exit__ (optimized away) 
      if_stmt_455_x_xentry_x_xx_x2596_symbol  <=  assign_stmt_439_to_assign_stmt_454_x_xexit_x_xx_x2595_symbol; -- place branch_block_stmt_405/if_stmt_455__entry__ (optimized away) 
      if_stmt_455_x_xexit_x_xx_x2597_symbol  <=  if_stmt_455_dead_link_2804_symbol; -- place branch_block_stmt_405/if_stmt_455__exit__ (optimized away) 
      merge_stmt_461_x_xentry_x_xx_x2598_symbol  <=  if_stmt_455_x_xexit_x_xx_x2597_symbol; -- place branch_block_stmt_405/merge_stmt_461__entry__ (optimized away) 
      merge_stmt_461_x_xexit_x_xx_x2599_symbol  <=  merge_stmt_461_dead_link_3265_symbol or merge_stmt_461_PhiAck_3273_symbol; -- place branch_block_stmt_405/merge_stmt_461__exit__ (optimized away) 
      assign_stmt_466_x_xentry_x_xx_x2600_symbol  <=  merge_stmt_461_x_xexit_x_xx_x2599_symbol; -- place branch_block_stmt_405/assign_stmt_466__entry__ (optimized away) 
      assign_stmt_466_x_xexit_x_xx_x2601_symbol  <=  assign_stmt_466_2823_symbol; -- place branch_block_stmt_405/assign_stmt_466__exit__ (optimized away) 
      assign_stmt_470_x_xentry_x_xx_x2602_symbol  <=  assign_stmt_466_x_xexit_x_xx_x2601_symbol; -- place branch_block_stmt_405/assign_stmt_470__entry__ (optimized away) 
      assign_stmt_470_x_xexit_x_xx_x2603_symbol  <=  assign_stmt_470_2826_symbol; -- place branch_block_stmt_405/assign_stmt_470__exit__ (optimized away) 
      assign_stmt_474_to_assign_stmt_504_x_xentry_x_xx_x2604_symbol  <=  assign_stmt_470_x_xexit_x_xx_x2603_symbol; -- place branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504__entry__ (optimized away) 
      assign_stmt_474_to_assign_stmt_504_x_xexit_x_xx_x2605_symbol  <=  assign_stmt_474_to_assign_stmt_504_2844_symbol; -- place branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504__exit__ (optimized away) 
      assign_stmt_508_x_xentry_x_xx_x2606_symbol  <=  assign_stmt_474_to_assign_stmt_504_x_xexit_x_xx_x2605_symbol; -- place branch_block_stmt_405/assign_stmt_508__entry__ (optimized away) 
      assign_stmt_508_x_xexit_x_xx_x2607_symbol  <=  assign_stmt_508_3232_symbol; -- place branch_block_stmt_405/assign_stmt_508__exit__ (optimized away) 
      bb_2_bb_1_2608_symbol  <=  assign_stmt_508_x_xexit_x_xx_x2607_symbol; -- place branch_block_stmt_405/bb_2_bb_1 (optimized away) 
      assign_stmt_411_to_assign_stmt_415_2609: Block -- branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415 
        signal assign_stmt_411_to_assign_stmt_415_2609_start: Boolean;
        signal Xentry_2610_symbol: Boolean;
        signal Xexit_2611_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_411_to_assign_stmt_415_2609_start <= assign_stmt_411_to_assign_stmt_415_x_xentry_x_xx_x2582_symbol; -- control passed to block
        Xentry_2610_symbol  <= assign_stmt_411_to_assign_stmt_415_2609_start; -- transition branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415/$entry
        Xexit_2611_symbol <= Xentry_2610_symbol; -- transition branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415/$exit
        assign_stmt_411_to_assign_stmt_415_2609_symbol <= Xexit_2611_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415
      assign_stmt_422_2612: Block -- branch_block_stmt_405/assign_stmt_422 
        signal assign_stmt_422_2612_start: Boolean;
        signal Xentry_2613_symbol: Boolean;
        signal Xexit_2614_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_422_2612_start <= assign_stmt_422_x_xentry_x_xx_x2586_symbol; -- control passed to block
        Xentry_2613_symbol  <= assign_stmt_422_2612_start; -- transition branch_block_stmt_405/assign_stmt_422/$entry
        Xexit_2614_symbol <= Xentry_2613_symbol; -- transition branch_block_stmt_405/assign_stmt_422/$exit
        assign_stmt_422_2612_symbol <= Xexit_2614_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_422
      assign_stmt_426_2615: Block -- branch_block_stmt_405/assign_stmt_426 
        signal assign_stmt_426_2615_start: Boolean;
        signal Xentry_2616_symbol: Boolean;
        signal Xexit_2617_symbol: Boolean;
        signal assign_stmt_426_active_x_x2618_symbol : Boolean;
        signal assign_stmt_426_completed_x_x2619_symbol : Boolean;
        signal simple_obj_ref_423_trigger_x_x2620_symbol : Boolean;
        signal simple_obj_ref_423_complete_2621_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_426_2615_start <= assign_stmt_426_x_xentry_x_xx_x2588_symbol; -- control passed to block
        Xentry_2616_symbol  <= assign_stmt_426_2615_start; -- transition branch_block_stmt_405/assign_stmt_426/$entry
        assign_stmt_426_active_x_x2618_symbol <= Xentry_2616_symbol; -- transition branch_block_stmt_405/assign_stmt_426/assign_stmt_426_active_
        assign_stmt_426_completed_x_x2619_symbol <= simple_obj_ref_423_complete_2621_symbol; -- transition branch_block_stmt_405/assign_stmt_426/assign_stmt_426_completed_
        simple_obj_ref_423_trigger_x_x2620_symbol <= assign_stmt_426_active_x_x2618_symbol; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_trigger_
        simple_obj_ref_423_complete_2621: Block -- branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete 
          signal simple_obj_ref_423_complete_2621_start: Boolean;
          signal Xentry_2622_symbol: Boolean;
          signal Xexit_2623_symbol: Boolean;
          signal pipe_wreq_2624_symbol : Boolean;
          signal pipe_wack_2625_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_423_complete_2621_start <= simple_obj_ref_423_trigger_x_x2620_symbol; -- control passed to block
          Xentry_2622_symbol  <= simple_obj_ref_423_complete_2621_start; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/$entry
          pipe_wreq_2624_symbol <= Xentry_2622_symbol; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/pipe_wreq
          simple_obj_ref_423_inst_req_0 <= pipe_wreq_2624_symbol; -- link to DP
          pipe_wack_2625_symbol <= simple_obj_ref_423_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/pipe_wack
          Xexit_2623_symbol <= pipe_wack_2625_symbol; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/$exit
          simple_obj_ref_423_complete_2621_symbol <= Xexit_2623_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete
        Xexit_2617_symbol <= assign_stmt_426_completed_x_x2619_symbol; -- transition branch_block_stmt_405/assign_stmt_426/$exit
        assign_stmt_426_2615_symbol <= Xexit_2617_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_426
      assign_stmt_431_2626: Block -- branch_block_stmt_405/assign_stmt_431 
        signal assign_stmt_431_2626_start: Boolean;
        signal Xentry_2627_symbol: Boolean;
        signal Xexit_2628_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_431_2626_start <= assign_stmt_431_x_xentry_x_xx_x2590_symbol; -- control passed to block
        Xentry_2627_symbol  <= assign_stmt_431_2626_start; -- transition branch_block_stmt_405/assign_stmt_431/$entry
        Xexit_2628_symbol <= Xentry_2627_symbol; -- transition branch_block_stmt_405/assign_stmt_431/$exit
        assign_stmt_431_2626_symbol <= Xexit_2628_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_431
      assign_stmt_435_2629: Block -- branch_block_stmt_405/assign_stmt_435 
        signal assign_stmt_435_2629_start: Boolean;
        signal Xentry_2630_symbol: Boolean;
        signal Xexit_2631_symbol: Boolean;
        signal assign_stmt_435_active_x_x2632_symbol : Boolean;
        signal assign_stmt_435_completed_x_x2633_symbol : Boolean;
        signal type_cast_434_active_x_x2634_symbol : Boolean;
        signal type_cast_434_trigger_x_x2635_symbol : Boolean;
        signal simple_obj_ref_433_trigger_x_x2636_symbol : Boolean;
        signal simple_obj_ref_433_complete_2637_symbol : Boolean;
        signal type_cast_434_complete_2642_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_435_2629_start <= assign_stmt_435_x_xentry_x_xx_x2592_symbol; -- control passed to block
        Xentry_2630_symbol  <= assign_stmt_435_2629_start; -- transition branch_block_stmt_405/assign_stmt_435/$entry
        assign_stmt_435_active_x_x2632_symbol <= type_cast_434_complete_2642_symbol; -- transition branch_block_stmt_405/assign_stmt_435/assign_stmt_435_active_
        assign_stmt_435_completed_x_x2633_symbol <= assign_stmt_435_active_x_x2632_symbol; -- transition branch_block_stmt_405/assign_stmt_435/assign_stmt_435_completed_
        type_cast_434_active_x_x2634_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_435/type_cast_434_active_ 
          signal type_cast_434_active_x_x2634_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_434_active_x_x2634_predecessors(0) <= type_cast_434_trigger_x_x2635_symbol;
          type_cast_434_active_x_x2634_predecessors(1) <= simple_obj_ref_433_complete_2637_symbol;
          type_cast_434_active_x_x2634_join: join -- 
            port map( -- 
              preds => type_cast_434_active_x_x2634_predecessors,
              symbol_out => type_cast_434_active_x_x2634_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_435/type_cast_434_active_
        type_cast_434_trigger_x_x2635_symbol <= Xentry_2630_symbol; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_trigger_
        simple_obj_ref_433_trigger_x_x2636_symbol <= Xentry_2630_symbol; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_trigger_
        simple_obj_ref_433_complete_2637: Block -- branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete 
          signal simple_obj_ref_433_complete_2637_start: Boolean;
          signal Xentry_2638_symbol: Boolean;
          signal Xexit_2639_symbol: Boolean;
          signal req_2640_symbol : Boolean;
          signal ack_2641_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_433_complete_2637_start <= simple_obj_ref_433_trigger_x_x2636_symbol; -- control passed to block
          Xentry_2638_symbol  <= simple_obj_ref_433_complete_2637_start; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/$entry
          req_2640_symbol <= Xentry_2638_symbol; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/req
          simple_obj_ref_433_inst_req_0 <= req_2640_symbol; -- link to DP
          ack_2641_symbol <= simple_obj_ref_433_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/ack
          Xexit_2639_symbol <= ack_2641_symbol; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/$exit
          simple_obj_ref_433_complete_2637_symbol <= Xexit_2639_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete
        type_cast_434_complete_2642: Block -- branch_block_stmt_405/assign_stmt_435/type_cast_434_complete 
          signal type_cast_434_complete_2642_start: Boolean;
          signal Xentry_2643_symbol: Boolean;
          signal Xexit_2644_symbol: Boolean;
          signal req_2645_symbol : Boolean;
          signal ack_2646_symbol : Boolean;
          -- 
        begin -- 
          type_cast_434_complete_2642_start <= type_cast_434_active_x_x2634_symbol; -- control passed to block
          Xentry_2643_symbol  <= type_cast_434_complete_2642_start; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/$entry
          req_2645_symbol <= Xentry_2643_symbol; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/req
          type_cast_434_inst_req_0 <= req_2645_symbol; -- link to DP
          ack_2646_symbol <= type_cast_434_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/ack
          Xexit_2644_symbol <= ack_2646_symbol; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/$exit
          type_cast_434_complete_2642_symbol <= Xexit_2644_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_435/type_cast_434_complete
        Xexit_2631_symbol <= assign_stmt_435_completed_x_x2633_symbol; -- transition branch_block_stmt_405/assign_stmt_435/$exit
        assign_stmt_435_2629_symbol <= Xexit_2631_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_435
      assign_stmt_439_to_assign_stmt_454_2647: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454 
        signal assign_stmt_439_to_assign_stmt_454_2647_start: Boolean;
        signal Xentry_2648_symbol: Boolean;
        signal Xexit_2649_symbol: Boolean;
        signal assign_stmt_439_active_x_x2650_symbol : Boolean;
        signal assign_stmt_439_completed_x_x2651_symbol : Boolean;
        signal type_cast_438_active_x_x2652_symbol : Boolean;
        signal type_cast_438_trigger_x_x2653_symbol : Boolean;
        signal simple_obj_ref_437_complete_2654_symbol : Boolean;
        signal type_cast_438_complete_2655_symbol : Boolean;
        signal assign_stmt_443_active_x_x2660_symbol : Boolean;
        signal assign_stmt_443_completed_x_x2661_symbol : Boolean;
        signal simple_obj_ref_442_complete_2662_symbol : Boolean;
        signal ptr_deref_441_trigger_x_x2663_symbol : Boolean;
        signal ptr_deref_441_active_x_x2664_symbol : Boolean;
        signal ptr_deref_441_base_address_calculated_2665_symbol : Boolean;
        signal ptr_deref_441_root_address_calculated_2666_symbol : Boolean;
        signal ptr_deref_441_word_address_calculated_2667_symbol : Boolean;
        signal ptr_deref_441_request_2668_symbol : Boolean;
        signal ptr_deref_441_complete_2696_symbol : Boolean;
        signal assign_stmt_447_active_x_x2722_symbol : Boolean;
        signal assign_stmt_447_completed_x_x2723_symbol : Boolean;
        signal ptr_deref_446_trigger_x_x2724_symbol : Boolean;
        signal ptr_deref_446_active_x_x2725_symbol : Boolean;
        signal ptr_deref_446_base_address_calculated_2726_symbol : Boolean;
        signal ptr_deref_446_root_address_calculated_2727_symbol : Boolean;
        signal ptr_deref_446_word_address_calculated_2728_symbol : Boolean;
        signal ptr_deref_446_request_2729_symbol : Boolean;
        signal ptr_deref_446_complete_2755_symbol : Boolean;
        signal assign_stmt_454_active_x_x2783_symbol : Boolean;
        signal assign_stmt_454_completed_x_x2784_symbol : Boolean;
        signal binary_453_active_x_x2785_symbol : Boolean;
        signal binary_453_trigger_x_x2786_symbol : Boolean;
        signal type_cast_450_active_x_x2787_symbol : Boolean;
        signal type_cast_450_trigger_x_x2788_symbol : Boolean;
        signal simple_obj_ref_449_complete_2789_symbol : Boolean;
        signal type_cast_450_complete_2790_symbol : Boolean;
        signal binary_453_complete_2797_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_439_to_assign_stmt_454_2647_start <= assign_stmt_439_to_assign_stmt_454_x_xentry_x_xx_x2594_symbol; -- control passed to block
        Xentry_2648_symbol  <= assign_stmt_439_to_assign_stmt_454_2647_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/$entry
        assign_stmt_439_active_x_x2650_symbol <= type_cast_438_complete_2655_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_439_active_
        assign_stmt_439_completed_x_x2651_symbol <= assign_stmt_439_active_x_x2650_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_439_completed_
        type_cast_438_active_x_x2652_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_active_ 
          signal type_cast_438_active_x_x2652_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_438_active_x_x2652_predecessors(0) <= type_cast_438_trigger_x_x2653_symbol;
          type_cast_438_active_x_x2652_predecessors(1) <= simple_obj_ref_437_complete_2654_symbol;
          type_cast_438_active_x_x2652_join: join -- 
            port map( -- 
              preds => type_cast_438_active_x_x2652_predecessors,
              symbol_out => type_cast_438_active_x_x2652_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_active_
        type_cast_438_trigger_x_x2653_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_trigger_
        simple_obj_ref_437_complete_2654_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/simple_obj_ref_437_complete
        type_cast_438_complete_2655: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete 
          signal type_cast_438_complete_2655_start: Boolean;
          signal Xentry_2656_symbol: Boolean;
          signal Xexit_2657_symbol: Boolean;
          signal req_2658_symbol : Boolean;
          signal ack_2659_symbol : Boolean;
          -- 
        begin -- 
          type_cast_438_complete_2655_start <= type_cast_438_active_x_x2652_symbol; -- control passed to block
          Xentry_2656_symbol  <= type_cast_438_complete_2655_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/$entry
          req_2658_symbol <= Xentry_2656_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/req
          type_cast_438_inst_req_0 <= req_2658_symbol; -- link to DP
          ack_2659_symbol <= type_cast_438_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/ack
          Xexit_2657_symbol <= ack_2659_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/$exit
          type_cast_438_complete_2655_symbol <= Xexit_2657_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete
        assign_stmt_443_active_x_x2660_symbol <= simple_obj_ref_442_complete_2662_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_443_active_
        assign_stmt_443_completed_x_x2661_symbol <= ptr_deref_441_complete_2696_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_443_completed_
        simple_obj_ref_442_complete_2662_symbol <= assign_stmt_439_completed_x_x2651_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/simple_obj_ref_442_complete
        ptr_deref_441_trigger_x_x2663_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_trigger_ 
          signal ptr_deref_441_trigger_x_x2663_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_441_trigger_x_x2663_predecessors(0) <= ptr_deref_441_word_address_calculated_2667_symbol;
          ptr_deref_441_trigger_x_x2663_predecessors(1) <= assign_stmt_443_active_x_x2660_symbol;
          ptr_deref_441_trigger_x_x2663_join: join -- 
            port map( -- 
              preds => ptr_deref_441_trigger_x_x2663_predecessors,
              symbol_out => ptr_deref_441_trigger_x_x2663_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_trigger_
        ptr_deref_441_active_x_x2664_symbol <= ptr_deref_441_request_2668_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_active_
        ptr_deref_441_base_address_calculated_2665_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_base_address_calculated
        ptr_deref_441_root_address_calculated_2666_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_root_address_calculated
        ptr_deref_441_word_address_calculated_2667_symbol <= ptr_deref_441_root_address_calculated_2666_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_word_address_calculated
        ptr_deref_441_request_2668: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request 
          signal ptr_deref_441_request_2668_start: Boolean;
          signal Xentry_2669_symbol: Boolean;
          signal Xexit_2670_symbol: Boolean;
          signal split_req_2671_symbol : Boolean;
          signal split_ack_2672_symbol : Boolean;
          signal word_access_2673_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_441_request_2668_start <= ptr_deref_441_trigger_x_x2663_symbol; -- control passed to block
          Xentry_2669_symbol  <= ptr_deref_441_request_2668_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/$entry
          split_req_2671_symbol <= Xentry_2669_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/split_req
          ptr_deref_441_gather_scatter_req_0 <= split_req_2671_symbol; -- link to DP
          split_ack_2672_symbol <= ptr_deref_441_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/split_ack
          word_access_2673: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access 
            signal word_access_2673_start: Boolean;
            signal Xentry_2674_symbol: Boolean;
            signal Xexit_2675_symbol: Boolean;
            signal word_access_0_2676_symbol : Boolean;
            signal word_access_1_2681_symbol : Boolean;
            signal word_access_2_2686_symbol : Boolean;
            signal word_access_3_2691_symbol : Boolean;
            -- 
          begin -- 
            word_access_2673_start <= split_ack_2672_symbol; -- control passed to block
            Xentry_2674_symbol  <= word_access_2673_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/$entry
            word_access_0_2676: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0 
              signal word_access_0_2676_start: Boolean;
              signal Xentry_2677_symbol: Boolean;
              signal Xexit_2678_symbol: Boolean;
              signal rr_2679_symbol : Boolean;
              signal ra_2680_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2676_start <= Xentry_2674_symbol; -- control passed to block
              Xentry_2677_symbol  <= word_access_0_2676_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/$entry
              rr_2679_symbol <= Xentry_2677_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/rr
              ptr_deref_441_store_0_req_0 <= rr_2679_symbol; -- link to DP
              ra_2680_symbol <= ptr_deref_441_store_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/ra
              Xexit_2678_symbol <= ra_2680_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/$exit
              word_access_0_2676_symbol <= Xexit_2678_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0
            word_access_1_2681: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_1 
              signal word_access_1_2681_start: Boolean;
              signal Xentry_2682_symbol: Boolean;
              signal Xexit_2683_symbol: Boolean;
              signal rr_2684_symbol : Boolean;
              signal ra_2685_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2681_start <= Xentry_2674_symbol; -- control passed to block
              Xentry_2682_symbol  <= word_access_1_2681_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_1/$entry
              rr_2684_symbol <= Xentry_2682_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_1/rr
              ptr_deref_441_store_1_req_0 <= rr_2684_symbol; -- link to DP
              ra_2685_symbol <= ptr_deref_441_store_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_1/ra
              Xexit_2683_symbol <= ra_2685_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_1/$exit
              word_access_1_2681_symbol <= Xexit_2683_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_1
            word_access_2_2686: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_2 
              signal word_access_2_2686_start: Boolean;
              signal Xentry_2687_symbol: Boolean;
              signal Xexit_2688_symbol: Boolean;
              signal rr_2689_symbol : Boolean;
              signal ra_2690_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2686_start <= Xentry_2674_symbol; -- control passed to block
              Xentry_2687_symbol  <= word_access_2_2686_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_2/$entry
              rr_2689_symbol <= Xentry_2687_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_2/rr
              ptr_deref_441_store_2_req_0 <= rr_2689_symbol; -- link to DP
              ra_2690_symbol <= ptr_deref_441_store_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_2/ra
              Xexit_2688_symbol <= ra_2690_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_2/$exit
              word_access_2_2686_symbol <= Xexit_2688_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_2
            word_access_3_2691: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_3 
              signal word_access_3_2691_start: Boolean;
              signal Xentry_2692_symbol: Boolean;
              signal Xexit_2693_symbol: Boolean;
              signal rr_2694_symbol : Boolean;
              signal ra_2695_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2691_start <= Xentry_2674_symbol; -- control passed to block
              Xentry_2692_symbol  <= word_access_3_2691_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_3/$entry
              rr_2694_symbol <= Xentry_2692_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_3/rr
              ptr_deref_441_store_3_req_0 <= rr_2694_symbol; -- link to DP
              ra_2695_symbol <= ptr_deref_441_store_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_3/ra
              Xexit_2693_symbol <= ra_2695_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_3/$exit
              word_access_3_2691_symbol <= Xexit_2693_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_3
            Xexit_2675_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/$exit 
              signal Xexit_2675_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2675_predecessors(0) <= word_access_0_2676_symbol;
              Xexit_2675_predecessors(1) <= word_access_1_2681_symbol;
              Xexit_2675_predecessors(2) <= word_access_2_2686_symbol;
              Xexit_2675_predecessors(3) <= word_access_3_2691_symbol;
              Xexit_2675_join: join -- 
                port map( -- 
                  preds => Xexit_2675_predecessors,
                  symbol_out => Xexit_2675_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/$exit
            word_access_2673_symbol <= Xexit_2675_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access
          Xexit_2670_symbol <= word_access_2673_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/$exit
          ptr_deref_441_request_2668_symbol <= Xexit_2670_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request
        ptr_deref_441_complete_2696: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete 
          signal ptr_deref_441_complete_2696_start: Boolean;
          signal Xentry_2697_symbol: Boolean;
          signal Xexit_2698_symbol: Boolean;
          signal word_access_2699_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_441_complete_2696_start <= ptr_deref_441_active_x_x2664_symbol; -- control passed to block
          Xentry_2697_symbol  <= ptr_deref_441_complete_2696_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/$entry
          word_access_2699: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access 
            signal word_access_2699_start: Boolean;
            signal Xentry_2700_symbol: Boolean;
            signal Xexit_2701_symbol: Boolean;
            signal word_access_0_2702_symbol : Boolean;
            signal word_access_1_2707_symbol : Boolean;
            signal word_access_2_2712_symbol : Boolean;
            signal word_access_3_2717_symbol : Boolean;
            -- 
          begin -- 
            word_access_2699_start <= Xentry_2697_symbol; -- control passed to block
            Xentry_2700_symbol  <= word_access_2699_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/$entry
            word_access_0_2702: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0 
              signal word_access_0_2702_start: Boolean;
              signal Xentry_2703_symbol: Boolean;
              signal Xexit_2704_symbol: Boolean;
              signal cr_2705_symbol : Boolean;
              signal ca_2706_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2702_start <= Xentry_2700_symbol; -- control passed to block
              Xentry_2703_symbol  <= word_access_0_2702_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/$entry
              cr_2705_symbol <= Xentry_2703_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/cr
              ptr_deref_441_store_0_req_1 <= cr_2705_symbol; -- link to DP
              ca_2706_symbol <= ptr_deref_441_store_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/ca
              Xexit_2704_symbol <= ca_2706_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/$exit
              word_access_0_2702_symbol <= Xexit_2704_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0
            word_access_1_2707: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_1 
              signal word_access_1_2707_start: Boolean;
              signal Xentry_2708_symbol: Boolean;
              signal Xexit_2709_symbol: Boolean;
              signal cr_2710_symbol : Boolean;
              signal ca_2711_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2707_start <= Xentry_2700_symbol; -- control passed to block
              Xentry_2708_symbol  <= word_access_1_2707_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_1/$entry
              cr_2710_symbol <= Xentry_2708_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_1/cr
              ptr_deref_441_store_1_req_1 <= cr_2710_symbol; -- link to DP
              ca_2711_symbol <= ptr_deref_441_store_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_1/ca
              Xexit_2709_symbol <= ca_2711_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_1/$exit
              word_access_1_2707_symbol <= Xexit_2709_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_1
            word_access_2_2712: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_2 
              signal word_access_2_2712_start: Boolean;
              signal Xentry_2713_symbol: Boolean;
              signal Xexit_2714_symbol: Boolean;
              signal cr_2715_symbol : Boolean;
              signal ca_2716_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2712_start <= Xentry_2700_symbol; -- control passed to block
              Xentry_2713_symbol  <= word_access_2_2712_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_2/$entry
              cr_2715_symbol <= Xentry_2713_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_2/cr
              ptr_deref_441_store_2_req_1 <= cr_2715_symbol; -- link to DP
              ca_2716_symbol <= ptr_deref_441_store_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_2/ca
              Xexit_2714_symbol <= ca_2716_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_2/$exit
              word_access_2_2712_symbol <= Xexit_2714_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_2
            word_access_3_2717: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_3 
              signal word_access_3_2717_start: Boolean;
              signal Xentry_2718_symbol: Boolean;
              signal Xexit_2719_symbol: Boolean;
              signal cr_2720_symbol : Boolean;
              signal ca_2721_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2717_start <= Xentry_2700_symbol; -- control passed to block
              Xentry_2718_symbol  <= word_access_3_2717_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_3/$entry
              cr_2720_symbol <= Xentry_2718_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_3/cr
              ptr_deref_441_store_3_req_1 <= cr_2720_symbol; -- link to DP
              ca_2721_symbol <= ptr_deref_441_store_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_3/ca
              Xexit_2719_symbol <= ca_2721_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_3/$exit
              word_access_3_2717_symbol <= Xexit_2719_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_3
            Xexit_2701_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/$exit 
              signal Xexit_2701_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2701_predecessors(0) <= word_access_0_2702_symbol;
              Xexit_2701_predecessors(1) <= word_access_1_2707_symbol;
              Xexit_2701_predecessors(2) <= word_access_2_2712_symbol;
              Xexit_2701_predecessors(3) <= word_access_3_2717_symbol;
              Xexit_2701_join: join -- 
                port map( -- 
                  preds => Xexit_2701_predecessors,
                  symbol_out => Xexit_2701_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/$exit
            word_access_2699_symbol <= Xexit_2701_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access
          Xexit_2698_symbol <= word_access_2699_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/$exit
          ptr_deref_441_complete_2696_symbol <= Xexit_2698_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete
        assign_stmt_447_active_x_x2722_symbol <= ptr_deref_446_complete_2755_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_447_active_
        assign_stmt_447_completed_x_x2723_symbol <= assign_stmt_447_active_x_x2722_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_447_completed_
        ptr_deref_446_trigger_x_x2724_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_trigger_ 
          signal ptr_deref_446_trigger_x_x2724_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_446_trigger_x_x2724_predecessors(0) <= ptr_deref_446_word_address_calculated_2728_symbol;
          ptr_deref_446_trigger_x_x2724_predecessors(1) <= ptr_deref_441_active_x_x2664_symbol;
          ptr_deref_446_trigger_x_x2724_join: join -- 
            port map( -- 
              preds => ptr_deref_446_trigger_x_x2724_predecessors,
              symbol_out => ptr_deref_446_trigger_x_x2724_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_trigger_
        ptr_deref_446_active_x_x2725_symbol <= ptr_deref_446_request_2729_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_active_
        ptr_deref_446_base_address_calculated_2726_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_base_address_calculated
        ptr_deref_446_root_address_calculated_2727_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_root_address_calculated
        ptr_deref_446_word_address_calculated_2728_symbol <= ptr_deref_446_root_address_calculated_2727_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_word_address_calculated
        ptr_deref_446_request_2729: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request 
          signal ptr_deref_446_request_2729_start: Boolean;
          signal Xentry_2730_symbol: Boolean;
          signal Xexit_2731_symbol: Boolean;
          signal word_access_2732_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_446_request_2729_start <= ptr_deref_446_trigger_x_x2724_symbol; -- control passed to block
          Xentry_2730_symbol  <= ptr_deref_446_request_2729_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/$entry
          word_access_2732: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access 
            signal word_access_2732_start: Boolean;
            signal Xentry_2733_symbol: Boolean;
            signal Xexit_2734_symbol: Boolean;
            signal word_access_0_2735_symbol : Boolean;
            signal word_access_1_2740_symbol : Boolean;
            signal word_access_2_2745_symbol : Boolean;
            signal word_access_3_2750_symbol : Boolean;
            -- 
          begin -- 
            word_access_2732_start <= Xentry_2730_symbol; -- control passed to block
            Xentry_2733_symbol  <= word_access_2732_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/$entry
            word_access_0_2735: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0 
              signal word_access_0_2735_start: Boolean;
              signal Xentry_2736_symbol: Boolean;
              signal Xexit_2737_symbol: Boolean;
              signal rr_2738_symbol : Boolean;
              signal ra_2739_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2735_start <= Xentry_2733_symbol; -- control passed to block
              Xentry_2736_symbol  <= word_access_0_2735_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/$entry
              rr_2738_symbol <= Xentry_2736_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/rr
              ptr_deref_446_load_0_req_0 <= rr_2738_symbol; -- link to DP
              ra_2739_symbol <= ptr_deref_446_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/ra
              Xexit_2737_symbol <= ra_2739_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/$exit
              word_access_0_2735_symbol <= Xexit_2737_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0
            word_access_1_2740: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_1 
              signal word_access_1_2740_start: Boolean;
              signal Xentry_2741_symbol: Boolean;
              signal Xexit_2742_symbol: Boolean;
              signal rr_2743_symbol : Boolean;
              signal ra_2744_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2740_start <= Xentry_2733_symbol; -- control passed to block
              Xentry_2741_symbol  <= word_access_1_2740_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_1/$entry
              rr_2743_symbol <= Xentry_2741_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_1/rr
              ptr_deref_446_load_1_req_0 <= rr_2743_symbol; -- link to DP
              ra_2744_symbol <= ptr_deref_446_load_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_1/ra
              Xexit_2742_symbol <= ra_2744_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_1/$exit
              word_access_1_2740_symbol <= Xexit_2742_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_1
            word_access_2_2745: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_2 
              signal word_access_2_2745_start: Boolean;
              signal Xentry_2746_symbol: Boolean;
              signal Xexit_2747_symbol: Boolean;
              signal rr_2748_symbol : Boolean;
              signal ra_2749_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2745_start <= Xentry_2733_symbol; -- control passed to block
              Xentry_2746_symbol  <= word_access_2_2745_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_2/$entry
              rr_2748_symbol <= Xentry_2746_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_2/rr
              ptr_deref_446_load_2_req_0 <= rr_2748_symbol; -- link to DP
              ra_2749_symbol <= ptr_deref_446_load_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_2/ra
              Xexit_2747_symbol <= ra_2749_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_2/$exit
              word_access_2_2745_symbol <= Xexit_2747_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_2
            word_access_3_2750: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_3 
              signal word_access_3_2750_start: Boolean;
              signal Xentry_2751_symbol: Boolean;
              signal Xexit_2752_symbol: Boolean;
              signal rr_2753_symbol : Boolean;
              signal ra_2754_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2750_start <= Xentry_2733_symbol; -- control passed to block
              Xentry_2751_symbol  <= word_access_3_2750_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_3/$entry
              rr_2753_symbol <= Xentry_2751_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_3/rr
              ptr_deref_446_load_3_req_0 <= rr_2753_symbol; -- link to DP
              ra_2754_symbol <= ptr_deref_446_load_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_3/ra
              Xexit_2752_symbol <= ra_2754_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_3/$exit
              word_access_3_2750_symbol <= Xexit_2752_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_3
            Xexit_2734_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/$exit 
              signal Xexit_2734_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2734_predecessors(0) <= word_access_0_2735_symbol;
              Xexit_2734_predecessors(1) <= word_access_1_2740_symbol;
              Xexit_2734_predecessors(2) <= word_access_2_2745_symbol;
              Xexit_2734_predecessors(3) <= word_access_3_2750_symbol;
              Xexit_2734_join: join -- 
                port map( -- 
                  preds => Xexit_2734_predecessors,
                  symbol_out => Xexit_2734_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/$exit
            word_access_2732_symbol <= Xexit_2734_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access
          Xexit_2731_symbol <= word_access_2732_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/$exit
          ptr_deref_446_request_2729_symbol <= Xexit_2731_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request
        ptr_deref_446_complete_2755: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete 
          signal ptr_deref_446_complete_2755_start: Boolean;
          signal Xentry_2756_symbol: Boolean;
          signal Xexit_2757_symbol: Boolean;
          signal word_access_2758_symbol : Boolean;
          signal merge_req_2781_symbol : Boolean;
          signal merge_ack_2782_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_446_complete_2755_start <= ptr_deref_446_active_x_x2725_symbol; -- control passed to block
          Xentry_2756_symbol  <= ptr_deref_446_complete_2755_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/$entry
          word_access_2758: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access 
            signal word_access_2758_start: Boolean;
            signal Xentry_2759_symbol: Boolean;
            signal Xexit_2760_symbol: Boolean;
            signal word_access_0_2761_symbol : Boolean;
            signal word_access_1_2766_symbol : Boolean;
            signal word_access_2_2771_symbol : Boolean;
            signal word_access_3_2776_symbol : Boolean;
            -- 
          begin -- 
            word_access_2758_start <= Xentry_2756_symbol; -- control passed to block
            Xentry_2759_symbol  <= word_access_2758_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/$entry
            word_access_0_2761: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0 
              signal word_access_0_2761_start: Boolean;
              signal Xentry_2762_symbol: Boolean;
              signal Xexit_2763_symbol: Boolean;
              signal cr_2764_symbol : Boolean;
              signal ca_2765_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2761_start <= Xentry_2759_symbol; -- control passed to block
              Xentry_2762_symbol  <= word_access_0_2761_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/$entry
              cr_2764_symbol <= Xentry_2762_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/cr
              ptr_deref_446_load_0_req_1 <= cr_2764_symbol; -- link to DP
              ca_2765_symbol <= ptr_deref_446_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/ca
              Xexit_2763_symbol <= ca_2765_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/$exit
              word_access_0_2761_symbol <= Xexit_2763_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0
            word_access_1_2766: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_1 
              signal word_access_1_2766_start: Boolean;
              signal Xentry_2767_symbol: Boolean;
              signal Xexit_2768_symbol: Boolean;
              signal cr_2769_symbol : Boolean;
              signal ca_2770_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2766_start <= Xentry_2759_symbol; -- control passed to block
              Xentry_2767_symbol  <= word_access_1_2766_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_1/$entry
              cr_2769_symbol <= Xentry_2767_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_1/cr
              ptr_deref_446_load_1_req_1 <= cr_2769_symbol; -- link to DP
              ca_2770_symbol <= ptr_deref_446_load_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_1/ca
              Xexit_2768_symbol <= ca_2770_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_1/$exit
              word_access_1_2766_symbol <= Xexit_2768_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_1
            word_access_2_2771: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_2 
              signal word_access_2_2771_start: Boolean;
              signal Xentry_2772_symbol: Boolean;
              signal Xexit_2773_symbol: Boolean;
              signal cr_2774_symbol : Boolean;
              signal ca_2775_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2771_start <= Xentry_2759_symbol; -- control passed to block
              Xentry_2772_symbol  <= word_access_2_2771_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_2/$entry
              cr_2774_symbol <= Xentry_2772_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_2/cr
              ptr_deref_446_load_2_req_1 <= cr_2774_symbol; -- link to DP
              ca_2775_symbol <= ptr_deref_446_load_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_2/ca
              Xexit_2773_symbol <= ca_2775_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_2/$exit
              word_access_2_2771_symbol <= Xexit_2773_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_2
            word_access_3_2776: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_3 
              signal word_access_3_2776_start: Boolean;
              signal Xentry_2777_symbol: Boolean;
              signal Xexit_2778_symbol: Boolean;
              signal cr_2779_symbol : Boolean;
              signal ca_2780_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2776_start <= Xentry_2759_symbol; -- control passed to block
              Xentry_2777_symbol  <= word_access_3_2776_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_3/$entry
              cr_2779_symbol <= Xentry_2777_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_3/cr
              ptr_deref_446_load_3_req_1 <= cr_2779_symbol; -- link to DP
              ca_2780_symbol <= ptr_deref_446_load_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_3/ca
              Xexit_2778_symbol <= ca_2780_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_3/$exit
              word_access_3_2776_symbol <= Xexit_2778_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_3
            Xexit_2760_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/$exit 
              signal Xexit_2760_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2760_predecessors(0) <= word_access_0_2761_symbol;
              Xexit_2760_predecessors(1) <= word_access_1_2766_symbol;
              Xexit_2760_predecessors(2) <= word_access_2_2771_symbol;
              Xexit_2760_predecessors(3) <= word_access_3_2776_symbol;
              Xexit_2760_join: join -- 
                port map( -- 
                  preds => Xexit_2760_predecessors,
                  symbol_out => Xexit_2760_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/$exit
            word_access_2758_symbol <= Xexit_2760_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access
          merge_req_2781_symbol <= word_access_2758_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/merge_req
          ptr_deref_446_gather_scatter_req_0 <= merge_req_2781_symbol; -- link to DP
          merge_ack_2782_symbol <= ptr_deref_446_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/merge_ack
          Xexit_2757_symbol <= merge_ack_2782_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/$exit
          ptr_deref_446_complete_2755_symbol <= Xexit_2757_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete
        assign_stmt_454_active_x_x2783_symbol <= binary_453_complete_2797_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_454_active_
        assign_stmt_454_completed_x_x2784_symbol <= assign_stmt_454_active_x_x2783_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_454_completed_
        binary_453_active_x_x2785_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_active_ 
          signal binary_453_active_x_x2785_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_453_active_x_x2785_predecessors(0) <= binary_453_trigger_x_x2786_symbol;
          binary_453_active_x_x2785_predecessors(1) <= type_cast_450_complete_2790_symbol;
          binary_453_active_x_x2785_join: join -- 
            port map( -- 
              preds => binary_453_active_x_x2785_predecessors,
              symbol_out => binary_453_active_x_x2785_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_active_
        binary_453_trigger_x_x2786_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_trigger_
        type_cast_450_active_x_x2787_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_active_ 
          signal type_cast_450_active_x_x2787_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_450_active_x_x2787_predecessors(0) <= type_cast_450_trigger_x_x2788_symbol;
          type_cast_450_active_x_x2787_predecessors(1) <= simple_obj_ref_449_complete_2789_symbol;
          type_cast_450_active_x_x2787_join: join -- 
            port map( -- 
              preds => type_cast_450_active_x_x2787_predecessors,
              symbol_out => type_cast_450_active_x_x2787_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_active_
        type_cast_450_trigger_x_x2788_symbol <= Xentry_2648_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_trigger_
        simple_obj_ref_449_complete_2789_symbol <= assign_stmt_447_completed_x_x2723_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/simple_obj_ref_449_complete
        type_cast_450_complete_2790: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete 
          signal type_cast_450_complete_2790_start: Boolean;
          signal Xentry_2791_symbol: Boolean;
          signal Xexit_2792_symbol: Boolean;
          signal rr_2793_symbol : Boolean;
          signal ra_2794_symbol : Boolean;
          signal cr_2795_symbol : Boolean;
          signal ca_2796_symbol : Boolean;
          -- 
        begin -- 
          type_cast_450_complete_2790_start <= type_cast_450_active_x_x2787_symbol; -- control passed to block
          Xentry_2791_symbol  <= type_cast_450_complete_2790_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/$entry
          rr_2793_symbol <= Xentry_2791_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/rr
          type_cast_450_inst_req_0 <= rr_2793_symbol; -- link to DP
          ra_2794_symbol <= type_cast_450_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/ra
          cr_2795_symbol <= ra_2794_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/cr
          type_cast_450_inst_req_1 <= cr_2795_symbol; -- link to DP
          ca_2796_symbol <= type_cast_450_inst_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/ca
          Xexit_2792_symbol <= ca_2796_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/$exit
          type_cast_450_complete_2790_symbol <= Xexit_2792_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete
        binary_453_complete_2797: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete 
          signal binary_453_complete_2797_start: Boolean;
          signal Xentry_2798_symbol: Boolean;
          signal Xexit_2799_symbol: Boolean;
          signal rr_2800_symbol : Boolean;
          signal ra_2801_symbol : Boolean;
          signal cr_2802_symbol : Boolean;
          signal ca_2803_symbol : Boolean;
          -- 
        begin -- 
          binary_453_complete_2797_start <= binary_453_active_x_x2785_symbol; -- control passed to block
          Xentry_2798_symbol  <= binary_453_complete_2797_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/$entry
          rr_2800_symbol <= Xentry_2798_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/rr
          binary_453_inst_req_0 <= rr_2800_symbol; -- link to DP
          ra_2801_symbol <= binary_453_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/ra
          cr_2802_symbol <= ra_2801_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/cr
          binary_453_inst_req_1 <= cr_2802_symbol; -- link to DP
          ca_2803_symbol <= binary_453_inst_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/ca
          Xexit_2799_symbol <= ca_2803_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/$exit
          binary_453_complete_2797_symbol <= Xexit_2799_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete
        Xexit_2649_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/$exit 
          signal Xexit_2649_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          Xexit_2649_predecessors(0) <= assign_stmt_443_completed_x_x2661_symbol;
          Xexit_2649_predecessors(1) <= ptr_deref_441_base_address_calculated_2665_symbol;
          Xexit_2649_predecessors(2) <= ptr_deref_446_base_address_calculated_2726_symbol;
          Xexit_2649_predecessors(3) <= assign_stmt_454_completed_x_x2784_symbol;
          Xexit_2649_join: join -- 
            port map( -- 
              preds => Xexit_2649_predecessors,
              symbol_out => Xexit_2649_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/$exit
        assign_stmt_439_to_assign_stmt_454_2647_symbol <= Xexit_2649_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454
      if_stmt_455_dead_link_2804: Block -- branch_block_stmt_405/if_stmt_455_dead_link 
        signal if_stmt_455_dead_link_2804_start: Boolean;
        signal Xentry_2805_symbol: Boolean;
        signal Xexit_2806_symbol: Boolean;
        signal dead_transition_2807_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_dead_link_2804_start <= if_stmt_455_x_xentry_x_xx_x2596_symbol; -- control passed to block
        Xentry_2805_symbol  <= if_stmt_455_dead_link_2804_start; -- transition branch_block_stmt_405/if_stmt_455_dead_link/$entry
        dead_transition_2807_symbol <= false;
        Xexit_2806_symbol <= dead_transition_2807_symbol; -- transition branch_block_stmt_405/if_stmt_455_dead_link/$exit
        if_stmt_455_dead_link_2804_symbol <= Xexit_2806_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_dead_link
      if_stmt_455_eval_test_2808: Block -- branch_block_stmt_405/if_stmt_455_eval_test 
        signal if_stmt_455_eval_test_2808_start: Boolean;
        signal Xentry_2809_symbol: Boolean;
        signal Xexit_2810_symbol: Boolean;
        signal branch_req_2811_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_eval_test_2808_start <= if_stmt_455_x_xentry_x_xx_x2596_symbol; -- control passed to block
        Xentry_2809_symbol  <= if_stmt_455_eval_test_2808_start; -- transition branch_block_stmt_405/if_stmt_455_eval_test/$entry
        branch_req_2811_symbol <= Xentry_2809_symbol; -- transition branch_block_stmt_405/if_stmt_455_eval_test/branch_req
        if_stmt_455_branch_req_0 <= branch_req_2811_symbol; -- link to DP
        Xexit_2810_symbol <= branch_req_2811_symbol; -- transition branch_block_stmt_405/if_stmt_455_eval_test/$exit
        if_stmt_455_eval_test_2808_symbol <= Xexit_2810_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_eval_test
      simple_obj_ref_456_place_2812_symbol  <=  if_stmt_455_eval_test_2808_symbol; -- place branch_block_stmt_405/simple_obj_ref_456_place (optimized away) 
      if_stmt_455_if_link_2813: Block -- branch_block_stmt_405/if_stmt_455_if_link 
        signal if_stmt_455_if_link_2813_start: Boolean;
        signal Xentry_2814_symbol: Boolean;
        signal Xexit_2815_symbol: Boolean;
        signal if_choice_transition_2816_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_if_link_2813_start <= simple_obj_ref_456_place_2812_symbol; -- control passed to block
        Xentry_2814_symbol  <= if_stmt_455_if_link_2813_start; -- transition branch_block_stmt_405/if_stmt_455_if_link/$entry
        if_choice_transition_2816_symbol <= if_stmt_455_branch_ack_1; -- transition branch_block_stmt_405/if_stmt_455_if_link/if_choice_transition
        Xexit_2815_symbol <= if_choice_transition_2816_symbol; -- transition branch_block_stmt_405/if_stmt_455_if_link/$exit
        if_stmt_455_if_link_2813_symbol <= Xexit_2815_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_if_link
      if_stmt_455_else_link_2817: Block -- branch_block_stmt_405/if_stmt_455_else_link 
        signal if_stmt_455_else_link_2817_start: Boolean;
        signal Xentry_2818_symbol: Boolean;
        signal Xexit_2819_symbol: Boolean;
        signal else_choice_transition_2820_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_else_link_2817_start <= simple_obj_ref_456_place_2812_symbol; -- control passed to block
        Xentry_2818_symbol  <= if_stmt_455_else_link_2817_start; -- transition branch_block_stmt_405/if_stmt_455_else_link/$entry
        else_choice_transition_2820_symbol <= if_stmt_455_branch_ack_0; -- transition branch_block_stmt_405/if_stmt_455_else_link/else_choice_transition
        Xexit_2819_symbol <= else_choice_transition_2820_symbol; -- transition branch_block_stmt_405/if_stmt_455_else_link/$exit
        if_stmt_455_else_link_2817_symbol <= Xexit_2819_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_else_link
      bb_1_bb_2_2821_symbol  <=  if_stmt_455_if_link_2813_symbol; -- place branch_block_stmt_405/bb_1_bb_2 (optimized away) 
      bb_1_bb_1_2822_symbol  <=  if_stmt_455_else_link_2817_symbol; -- place branch_block_stmt_405/bb_1_bb_1 (optimized away) 
      assign_stmt_466_2823: Block -- branch_block_stmt_405/assign_stmt_466 
        signal assign_stmt_466_2823_start: Boolean;
        signal Xentry_2824_symbol: Boolean;
        signal Xexit_2825_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_466_2823_start <= assign_stmt_466_x_xentry_x_xx_x2600_symbol; -- control passed to block
        Xentry_2824_symbol  <= assign_stmt_466_2823_start; -- transition branch_block_stmt_405/assign_stmt_466/$entry
        Xexit_2825_symbol <= Xentry_2824_symbol; -- transition branch_block_stmt_405/assign_stmt_466/$exit
        assign_stmt_466_2823_symbol <= Xexit_2825_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_466
      assign_stmt_470_2826: Block -- branch_block_stmt_405/assign_stmt_470 
        signal assign_stmt_470_2826_start: Boolean;
        signal Xentry_2827_symbol: Boolean;
        signal Xexit_2828_symbol: Boolean;
        signal assign_stmt_470_active_x_x2829_symbol : Boolean;
        signal assign_stmt_470_completed_x_x2830_symbol : Boolean;
        signal type_cast_469_active_x_x2831_symbol : Boolean;
        signal type_cast_469_trigger_x_x2832_symbol : Boolean;
        signal simple_obj_ref_468_trigger_x_x2833_symbol : Boolean;
        signal simple_obj_ref_468_complete_2834_symbol : Boolean;
        signal type_cast_469_complete_2839_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_470_2826_start <= assign_stmt_470_x_xentry_x_xx_x2602_symbol; -- control passed to block
        Xentry_2827_symbol  <= assign_stmt_470_2826_start; -- transition branch_block_stmt_405/assign_stmt_470/$entry
        assign_stmt_470_active_x_x2829_symbol <= type_cast_469_complete_2839_symbol; -- transition branch_block_stmt_405/assign_stmt_470/assign_stmt_470_active_
        assign_stmt_470_completed_x_x2830_symbol <= assign_stmt_470_active_x_x2829_symbol; -- transition branch_block_stmt_405/assign_stmt_470/assign_stmt_470_completed_
        type_cast_469_active_x_x2831_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_470/type_cast_469_active_ 
          signal type_cast_469_active_x_x2831_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_469_active_x_x2831_predecessors(0) <= type_cast_469_trigger_x_x2832_symbol;
          type_cast_469_active_x_x2831_predecessors(1) <= simple_obj_ref_468_complete_2834_symbol;
          type_cast_469_active_x_x2831_join: join -- 
            port map( -- 
              preds => type_cast_469_active_x_x2831_predecessors,
              symbol_out => type_cast_469_active_x_x2831_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_470/type_cast_469_active_
        type_cast_469_trigger_x_x2832_symbol <= Xentry_2827_symbol; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_trigger_
        simple_obj_ref_468_trigger_x_x2833_symbol <= Xentry_2827_symbol; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_trigger_
        simple_obj_ref_468_complete_2834: Block -- branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete 
          signal simple_obj_ref_468_complete_2834_start: Boolean;
          signal Xentry_2835_symbol: Boolean;
          signal Xexit_2836_symbol: Boolean;
          signal req_2837_symbol : Boolean;
          signal ack_2838_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_468_complete_2834_start <= simple_obj_ref_468_trigger_x_x2833_symbol; -- control passed to block
          Xentry_2835_symbol  <= simple_obj_ref_468_complete_2834_start; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/$entry
          req_2837_symbol <= Xentry_2835_symbol; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/req
          simple_obj_ref_468_inst_req_0 <= req_2837_symbol; -- link to DP
          ack_2838_symbol <= simple_obj_ref_468_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/ack
          Xexit_2836_symbol <= ack_2838_symbol; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/$exit
          simple_obj_ref_468_complete_2834_symbol <= Xexit_2836_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete
        type_cast_469_complete_2839: Block -- branch_block_stmt_405/assign_stmt_470/type_cast_469_complete 
          signal type_cast_469_complete_2839_start: Boolean;
          signal Xentry_2840_symbol: Boolean;
          signal Xexit_2841_symbol: Boolean;
          signal req_2842_symbol : Boolean;
          signal ack_2843_symbol : Boolean;
          -- 
        begin -- 
          type_cast_469_complete_2839_start <= type_cast_469_active_x_x2831_symbol; -- control passed to block
          Xentry_2840_symbol  <= type_cast_469_complete_2839_start; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/$entry
          req_2842_symbol <= Xentry_2840_symbol; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/req
          type_cast_469_inst_req_0 <= req_2842_symbol; -- link to DP
          ack_2843_symbol <= type_cast_469_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/ack
          Xexit_2841_symbol <= ack_2843_symbol; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/$exit
          type_cast_469_complete_2839_symbol <= Xexit_2841_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_470/type_cast_469_complete
        Xexit_2828_symbol <= assign_stmt_470_completed_x_x2830_symbol; -- transition branch_block_stmt_405/assign_stmt_470/$exit
        assign_stmt_470_2826_symbol <= Xexit_2828_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_470
      assign_stmt_474_to_assign_stmt_504_2844: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504 
        signal assign_stmt_474_to_assign_stmt_504_2844_start: Boolean;
        signal Xentry_2845_symbol: Boolean;
        signal Xexit_2846_symbol: Boolean;
        signal assign_stmt_474_active_x_x2847_symbol : Boolean;
        signal assign_stmt_474_completed_x_x2848_symbol : Boolean;
        signal simple_obj_ref_473_complete_2849_symbol : Boolean;
        signal ptr_deref_472_trigger_x_x2850_symbol : Boolean;
        signal ptr_deref_472_active_x_x2851_symbol : Boolean;
        signal ptr_deref_472_base_address_calculated_2852_symbol : Boolean;
        signal ptr_deref_472_root_address_calculated_2853_symbol : Boolean;
        signal ptr_deref_472_word_address_calculated_2854_symbol : Boolean;
        signal ptr_deref_472_request_2855_symbol : Boolean;
        signal ptr_deref_472_complete_2883_symbol : Boolean;
        signal assign_stmt_478_active_x_x2909_symbol : Boolean;
        signal assign_stmt_478_completed_x_x2910_symbol : Boolean;
        signal ptr_deref_477_trigger_x_x2911_symbol : Boolean;
        signal ptr_deref_477_active_x_x2912_symbol : Boolean;
        signal ptr_deref_477_base_address_calculated_2913_symbol : Boolean;
        signal ptr_deref_477_root_address_calculated_2914_symbol : Boolean;
        signal ptr_deref_477_word_address_calculated_2915_symbol : Boolean;
        signal ptr_deref_477_request_2916_symbol : Boolean;
        signal ptr_deref_477_complete_2942_symbol : Boolean;
        signal assign_stmt_482_active_x_x2970_symbol : Boolean;
        signal assign_stmt_482_completed_x_x2971_symbol : Boolean;
        signal ptr_deref_481_trigger_x_x2972_symbol : Boolean;
        signal ptr_deref_481_active_x_x2973_symbol : Boolean;
        signal ptr_deref_481_base_address_calculated_2974_symbol : Boolean;
        signal ptr_deref_481_root_address_calculated_2975_symbol : Boolean;
        signal ptr_deref_481_word_address_calculated_2976_symbol : Boolean;
        signal ptr_deref_481_request_2977_symbol : Boolean;
        signal ptr_deref_481_complete_3003_symbol : Boolean;
        signal assign_stmt_487_active_x_x3031_symbol : Boolean;
        signal assign_stmt_487_completed_x_x3032_symbol : Boolean;
        signal array_obj_ref_486_trigger_x_x3033_symbol : Boolean;
        signal array_obj_ref_486_active_x_x3034_symbol : Boolean;
        signal array_obj_ref_486_base_address_calculated_3035_symbol : Boolean;
        signal array_obj_ref_486_root_address_calculated_3036_symbol : Boolean;
        signal array_obj_ref_486_base_address_resized_3037_symbol : Boolean;
        signal array_obj_ref_486_base_addr_resize_3038_symbol : Boolean;
        signal array_obj_ref_486_base_plus_offset_trigger_3043_symbol : Boolean;
        signal array_obj_ref_486_base_plus_offset_3044_symbol : Boolean;
        signal array_obj_ref_486_complete_3051_symbol : Boolean;
        signal assign_stmt_491_active_x_x3056_symbol : Boolean;
        signal assign_stmt_491_completed_x_x3057_symbol : Boolean;
        signal simple_obj_ref_490_complete_3058_symbol : Boolean;
        signal ptr_deref_489_trigger_x_x3059_symbol : Boolean;
        signal ptr_deref_489_active_x_x3060_symbol : Boolean;
        signal ptr_deref_489_base_address_calculated_3061_symbol : Boolean;
        signal simple_obj_ref_488_complete_3062_symbol : Boolean;
        signal ptr_deref_489_root_address_calculated_3063_symbol : Boolean;
        signal ptr_deref_489_word_address_calculated_3064_symbol : Boolean;
        signal ptr_deref_489_base_address_resized_3065_symbol : Boolean;
        signal ptr_deref_489_base_addr_resize_3066_symbol : Boolean;
        signal ptr_deref_489_base_plus_offset_3071_symbol : Boolean;
        signal ptr_deref_489_word_addrgen_3076_symbol : Boolean;
        signal ptr_deref_489_request_3107_symbol : Boolean;
        signal ptr_deref_489_complete_3135_symbol : Boolean;
        signal assign_stmt_495_active_x_x3161_symbol : Boolean;
        signal assign_stmt_495_completed_x_x3162_symbol : Boolean;
        signal ptr_deref_494_trigger_x_x3163_symbol : Boolean;
        signal ptr_deref_494_active_x_x3164_symbol : Boolean;
        signal ptr_deref_494_base_address_calculated_3165_symbol : Boolean;
        signal ptr_deref_494_root_address_calculated_3166_symbol : Boolean;
        signal ptr_deref_494_word_address_calculated_3167_symbol : Boolean;
        signal ptr_deref_494_request_3168_symbol : Boolean;
        signal ptr_deref_494_complete_3194_symbol : Boolean;
        signal assign_stmt_499_active_x_x3222_symbol : Boolean;
        signal assign_stmt_499_completed_x_x3223_symbol : Boolean;
        signal type_cast_498_active_x_x3224_symbol : Boolean;
        signal type_cast_498_trigger_x_x3225_symbol : Boolean;
        signal simple_obj_ref_497_complete_3226_symbol : Boolean;
        signal type_cast_498_complete_3227_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_474_to_assign_stmt_504_2844_start <= assign_stmt_474_to_assign_stmt_504_x_xentry_x_xx_x2604_symbol; -- control passed to block
        Xentry_2845_symbol  <= assign_stmt_474_to_assign_stmt_504_2844_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/$entry
        assign_stmt_474_active_x_x2847_symbol <= simple_obj_ref_473_complete_2849_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_474_active_
        assign_stmt_474_completed_x_x2848_symbol <= ptr_deref_472_complete_2883_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_474_completed_
        simple_obj_ref_473_complete_2849_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_473_complete
        ptr_deref_472_trigger_x_x2850_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_trigger_ 
          signal ptr_deref_472_trigger_x_x2850_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_472_trigger_x_x2850_predecessors(0) <= ptr_deref_472_word_address_calculated_2854_symbol;
          ptr_deref_472_trigger_x_x2850_predecessors(1) <= assign_stmt_474_active_x_x2847_symbol;
          ptr_deref_472_trigger_x_x2850_join: join -- 
            port map( -- 
              preds => ptr_deref_472_trigger_x_x2850_predecessors,
              symbol_out => ptr_deref_472_trigger_x_x2850_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_trigger_
        ptr_deref_472_active_x_x2851_symbol <= ptr_deref_472_request_2855_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_active_
        ptr_deref_472_base_address_calculated_2852_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_base_address_calculated
        ptr_deref_472_root_address_calculated_2853_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_root_address_calculated
        ptr_deref_472_word_address_calculated_2854_symbol <= ptr_deref_472_root_address_calculated_2853_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_word_address_calculated
        ptr_deref_472_request_2855: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request 
          signal ptr_deref_472_request_2855_start: Boolean;
          signal Xentry_2856_symbol: Boolean;
          signal Xexit_2857_symbol: Boolean;
          signal split_req_2858_symbol : Boolean;
          signal split_ack_2859_symbol : Boolean;
          signal word_access_2860_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_472_request_2855_start <= ptr_deref_472_trigger_x_x2850_symbol; -- control passed to block
          Xentry_2856_symbol  <= ptr_deref_472_request_2855_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/$entry
          split_req_2858_symbol <= Xentry_2856_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/split_req
          ptr_deref_472_gather_scatter_req_0 <= split_req_2858_symbol; -- link to DP
          split_ack_2859_symbol <= ptr_deref_472_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/split_ack
          word_access_2860: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access 
            signal word_access_2860_start: Boolean;
            signal Xentry_2861_symbol: Boolean;
            signal Xexit_2862_symbol: Boolean;
            signal word_access_0_2863_symbol : Boolean;
            signal word_access_1_2868_symbol : Boolean;
            signal word_access_2_2873_symbol : Boolean;
            signal word_access_3_2878_symbol : Boolean;
            -- 
          begin -- 
            word_access_2860_start <= split_ack_2859_symbol; -- control passed to block
            Xentry_2861_symbol  <= word_access_2860_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/$entry
            word_access_0_2863: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0 
              signal word_access_0_2863_start: Boolean;
              signal Xentry_2864_symbol: Boolean;
              signal Xexit_2865_symbol: Boolean;
              signal rr_2866_symbol : Boolean;
              signal ra_2867_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2863_start <= Xentry_2861_symbol; -- control passed to block
              Xentry_2864_symbol  <= word_access_0_2863_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/$entry
              rr_2866_symbol <= Xentry_2864_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/rr
              ptr_deref_472_store_0_req_0 <= rr_2866_symbol; -- link to DP
              ra_2867_symbol <= ptr_deref_472_store_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/ra
              Xexit_2865_symbol <= ra_2867_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/$exit
              word_access_0_2863_symbol <= Xexit_2865_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0
            word_access_1_2868: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_1 
              signal word_access_1_2868_start: Boolean;
              signal Xentry_2869_symbol: Boolean;
              signal Xexit_2870_symbol: Boolean;
              signal rr_2871_symbol : Boolean;
              signal ra_2872_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2868_start <= Xentry_2861_symbol; -- control passed to block
              Xentry_2869_symbol  <= word_access_1_2868_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_1/$entry
              rr_2871_symbol <= Xentry_2869_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_1/rr
              ptr_deref_472_store_1_req_0 <= rr_2871_symbol; -- link to DP
              ra_2872_symbol <= ptr_deref_472_store_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_1/ra
              Xexit_2870_symbol <= ra_2872_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_1/$exit
              word_access_1_2868_symbol <= Xexit_2870_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_1
            word_access_2_2873: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_2 
              signal word_access_2_2873_start: Boolean;
              signal Xentry_2874_symbol: Boolean;
              signal Xexit_2875_symbol: Boolean;
              signal rr_2876_symbol : Boolean;
              signal ra_2877_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2873_start <= Xentry_2861_symbol; -- control passed to block
              Xentry_2874_symbol  <= word_access_2_2873_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_2/$entry
              rr_2876_symbol <= Xentry_2874_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_2/rr
              ptr_deref_472_store_2_req_0 <= rr_2876_symbol; -- link to DP
              ra_2877_symbol <= ptr_deref_472_store_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_2/ra
              Xexit_2875_symbol <= ra_2877_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_2/$exit
              word_access_2_2873_symbol <= Xexit_2875_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_2
            word_access_3_2878: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_3 
              signal word_access_3_2878_start: Boolean;
              signal Xentry_2879_symbol: Boolean;
              signal Xexit_2880_symbol: Boolean;
              signal rr_2881_symbol : Boolean;
              signal ra_2882_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2878_start <= Xentry_2861_symbol; -- control passed to block
              Xentry_2879_symbol  <= word_access_3_2878_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_3/$entry
              rr_2881_symbol <= Xentry_2879_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_3/rr
              ptr_deref_472_store_3_req_0 <= rr_2881_symbol; -- link to DP
              ra_2882_symbol <= ptr_deref_472_store_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_3/ra
              Xexit_2880_symbol <= ra_2882_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_3/$exit
              word_access_3_2878_symbol <= Xexit_2880_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_3
            Xexit_2862_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/$exit 
              signal Xexit_2862_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2862_predecessors(0) <= word_access_0_2863_symbol;
              Xexit_2862_predecessors(1) <= word_access_1_2868_symbol;
              Xexit_2862_predecessors(2) <= word_access_2_2873_symbol;
              Xexit_2862_predecessors(3) <= word_access_3_2878_symbol;
              Xexit_2862_join: join -- 
                port map( -- 
                  preds => Xexit_2862_predecessors,
                  symbol_out => Xexit_2862_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/$exit
            word_access_2860_symbol <= Xexit_2862_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access
          Xexit_2857_symbol <= word_access_2860_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/$exit
          ptr_deref_472_request_2855_symbol <= Xexit_2857_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request
        ptr_deref_472_complete_2883: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete 
          signal ptr_deref_472_complete_2883_start: Boolean;
          signal Xentry_2884_symbol: Boolean;
          signal Xexit_2885_symbol: Boolean;
          signal word_access_2886_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_472_complete_2883_start <= ptr_deref_472_active_x_x2851_symbol; -- control passed to block
          Xentry_2884_symbol  <= ptr_deref_472_complete_2883_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/$entry
          word_access_2886: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access 
            signal word_access_2886_start: Boolean;
            signal Xentry_2887_symbol: Boolean;
            signal Xexit_2888_symbol: Boolean;
            signal word_access_0_2889_symbol : Boolean;
            signal word_access_1_2894_symbol : Boolean;
            signal word_access_2_2899_symbol : Boolean;
            signal word_access_3_2904_symbol : Boolean;
            -- 
          begin -- 
            word_access_2886_start <= Xentry_2884_symbol; -- control passed to block
            Xentry_2887_symbol  <= word_access_2886_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/$entry
            word_access_0_2889: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0 
              signal word_access_0_2889_start: Boolean;
              signal Xentry_2890_symbol: Boolean;
              signal Xexit_2891_symbol: Boolean;
              signal cr_2892_symbol : Boolean;
              signal ca_2893_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2889_start <= Xentry_2887_symbol; -- control passed to block
              Xentry_2890_symbol  <= word_access_0_2889_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/$entry
              cr_2892_symbol <= Xentry_2890_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/cr
              ptr_deref_472_store_0_req_1 <= cr_2892_symbol; -- link to DP
              ca_2893_symbol <= ptr_deref_472_store_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/ca
              Xexit_2891_symbol <= ca_2893_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/$exit
              word_access_0_2889_symbol <= Xexit_2891_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0
            word_access_1_2894: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_1 
              signal word_access_1_2894_start: Boolean;
              signal Xentry_2895_symbol: Boolean;
              signal Xexit_2896_symbol: Boolean;
              signal cr_2897_symbol : Boolean;
              signal ca_2898_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2894_start <= Xentry_2887_symbol; -- control passed to block
              Xentry_2895_symbol  <= word_access_1_2894_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_1/$entry
              cr_2897_symbol <= Xentry_2895_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_1/cr
              ptr_deref_472_store_1_req_1 <= cr_2897_symbol; -- link to DP
              ca_2898_symbol <= ptr_deref_472_store_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_1/ca
              Xexit_2896_symbol <= ca_2898_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_1/$exit
              word_access_1_2894_symbol <= Xexit_2896_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_1
            word_access_2_2899: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_2 
              signal word_access_2_2899_start: Boolean;
              signal Xentry_2900_symbol: Boolean;
              signal Xexit_2901_symbol: Boolean;
              signal cr_2902_symbol : Boolean;
              signal ca_2903_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2899_start <= Xentry_2887_symbol; -- control passed to block
              Xentry_2900_symbol  <= word_access_2_2899_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_2/$entry
              cr_2902_symbol <= Xentry_2900_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_2/cr
              ptr_deref_472_store_2_req_1 <= cr_2902_symbol; -- link to DP
              ca_2903_symbol <= ptr_deref_472_store_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_2/ca
              Xexit_2901_symbol <= ca_2903_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_2/$exit
              word_access_2_2899_symbol <= Xexit_2901_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_2
            word_access_3_2904: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_3 
              signal word_access_3_2904_start: Boolean;
              signal Xentry_2905_symbol: Boolean;
              signal Xexit_2906_symbol: Boolean;
              signal cr_2907_symbol : Boolean;
              signal ca_2908_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2904_start <= Xentry_2887_symbol; -- control passed to block
              Xentry_2905_symbol  <= word_access_3_2904_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_3/$entry
              cr_2907_symbol <= Xentry_2905_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_3/cr
              ptr_deref_472_store_3_req_1 <= cr_2907_symbol; -- link to DP
              ca_2908_symbol <= ptr_deref_472_store_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_3/ca
              Xexit_2906_symbol <= ca_2908_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_3/$exit
              word_access_3_2904_symbol <= Xexit_2906_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_3
            Xexit_2888_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/$exit 
              signal Xexit_2888_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2888_predecessors(0) <= word_access_0_2889_symbol;
              Xexit_2888_predecessors(1) <= word_access_1_2894_symbol;
              Xexit_2888_predecessors(2) <= word_access_2_2899_symbol;
              Xexit_2888_predecessors(3) <= word_access_3_2904_symbol;
              Xexit_2888_join: join -- 
                port map( -- 
                  preds => Xexit_2888_predecessors,
                  symbol_out => Xexit_2888_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/$exit
            word_access_2886_symbol <= Xexit_2888_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access
          Xexit_2885_symbol <= word_access_2886_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/$exit
          ptr_deref_472_complete_2883_symbol <= Xexit_2885_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete
        assign_stmt_478_active_x_x2909_symbol <= ptr_deref_477_complete_2942_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_478_active_
        assign_stmt_478_completed_x_x2910_symbol <= assign_stmt_478_active_x_x2909_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_478_completed_
        ptr_deref_477_trigger_x_x2911_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_trigger_ 
          signal ptr_deref_477_trigger_x_x2911_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_477_trigger_x_x2911_predecessors(0) <= ptr_deref_477_word_address_calculated_2915_symbol;
          ptr_deref_477_trigger_x_x2911_predecessors(1) <= ptr_deref_472_active_x_x2851_symbol;
          ptr_deref_477_trigger_x_x2911_join: join -- 
            port map( -- 
              preds => ptr_deref_477_trigger_x_x2911_predecessors,
              symbol_out => ptr_deref_477_trigger_x_x2911_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_trigger_
        ptr_deref_477_active_x_x2912_symbol <= ptr_deref_477_request_2916_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_active_
        ptr_deref_477_base_address_calculated_2913_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_base_address_calculated
        ptr_deref_477_root_address_calculated_2914_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_root_address_calculated
        ptr_deref_477_word_address_calculated_2915_symbol <= ptr_deref_477_root_address_calculated_2914_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_word_address_calculated
        ptr_deref_477_request_2916: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request 
          signal ptr_deref_477_request_2916_start: Boolean;
          signal Xentry_2917_symbol: Boolean;
          signal Xexit_2918_symbol: Boolean;
          signal word_access_2919_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_477_request_2916_start <= ptr_deref_477_trigger_x_x2911_symbol; -- control passed to block
          Xentry_2917_symbol  <= ptr_deref_477_request_2916_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/$entry
          word_access_2919: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access 
            signal word_access_2919_start: Boolean;
            signal Xentry_2920_symbol: Boolean;
            signal Xexit_2921_symbol: Boolean;
            signal word_access_0_2922_symbol : Boolean;
            signal word_access_1_2927_symbol : Boolean;
            signal word_access_2_2932_symbol : Boolean;
            signal word_access_3_2937_symbol : Boolean;
            -- 
          begin -- 
            word_access_2919_start <= Xentry_2917_symbol; -- control passed to block
            Xentry_2920_symbol  <= word_access_2919_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/$entry
            word_access_0_2922: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0 
              signal word_access_0_2922_start: Boolean;
              signal Xentry_2923_symbol: Boolean;
              signal Xexit_2924_symbol: Boolean;
              signal rr_2925_symbol : Boolean;
              signal ra_2926_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2922_start <= Xentry_2920_symbol; -- control passed to block
              Xentry_2923_symbol  <= word_access_0_2922_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/$entry
              rr_2925_symbol <= Xentry_2923_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/rr
              ptr_deref_477_load_0_req_0 <= rr_2925_symbol; -- link to DP
              ra_2926_symbol <= ptr_deref_477_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/ra
              Xexit_2924_symbol <= ra_2926_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/$exit
              word_access_0_2922_symbol <= Xexit_2924_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0
            word_access_1_2927: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_1 
              signal word_access_1_2927_start: Boolean;
              signal Xentry_2928_symbol: Boolean;
              signal Xexit_2929_symbol: Boolean;
              signal rr_2930_symbol : Boolean;
              signal ra_2931_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2927_start <= Xentry_2920_symbol; -- control passed to block
              Xentry_2928_symbol  <= word_access_1_2927_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_1/$entry
              rr_2930_symbol <= Xentry_2928_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_1/rr
              ptr_deref_477_load_1_req_0 <= rr_2930_symbol; -- link to DP
              ra_2931_symbol <= ptr_deref_477_load_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_1/ra
              Xexit_2929_symbol <= ra_2931_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_1/$exit
              word_access_1_2927_symbol <= Xexit_2929_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_1
            word_access_2_2932: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_2 
              signal word_access_2_2932_start: Boolean;
              signal Xentry_2933_symbol: Boolean;
              signal Xexit_2934_symbol: Boolean;
              signal rr_2935_symbol : Boolean;
              signal ra_2936_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2932_start <= Xentry_2920_symbol; -- control passed to block
              Xentry_2933_symbol  <= word_access_2_2932_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_2/$entry
              rr_2935_symbol <= Xentry_2933_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_2/rr
              ptr_deref_477_load_2_req_0 <= rr_2935_symbol; -- link to DP
              ra_2936_symbol <= ptr_deref_477_load_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_2/ra
              Xexit_2934_symbol <= ra_2936_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_2/$exit
              word_access_2_2932_symbol <= Xexit_2934_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_2
            word_access_3_2937: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_3 
              signal word_access_3_2937_start: Boolean;
              signal Xentry_2938_symbol: Boolean;
              signal Xexit_2939_symbol: Boolean;
              signal rr_2940_symbol : Boolean;
              signal ra_2941_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2937_start <= Xentry_2920_symbol; -- control passed to block
              Xentry_2938_symbol  <= word_access_3_2937_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_3/$entry
              rr_2940_symbol <= Xentry_2938_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_3/rr
              ptr_deref_477_load_3_req_0 <= rr_2940_symbol; -- link to DP
              ra_2941_symbol <= ptr_deref_477_load_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_3/ra
              Xexit_2939_symbol <= ra_2941_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_3/$exit
              word_access_3_2937_symbol <= Xexit_2939_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_3
            Xexit_2921_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/$exit 
              signal Xexit_2921_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2921_predecessors(0) <= word_access_0_2922_symbol;
              Xexit_2921_predecessors(1) <= word_access_1_2927_symbol;
              Xexit_2921_predecessors(2) <= word_access_2_2932_symbol;
              Xexit_2921_predecessors(3) <= word_access_3_2937_symbol;
              Xexit_2921_join: join -- 
                port map( -- 
                  preds => Xexit_2921_predecessors,
                  symbol_out => Xexit_2921_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/$exit
            word_access_2919_symbol <= Xexit_2921_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access
          Xexit_2918_symbol <= word_access_2919_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/$exit
          ptr_deref_477_request_2916_symbol <= Xexit_2918_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request
        ptr_deref_477_complete_2942: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete 
          signal ptr_deref_477_complete_2942_start: Boolean;
          signal Xentry_2943_symbol: Boolean;
          signal Xexit_2944_symbol: Boolean;
          signal word_access_2945_symbol : Boolean;
          signal merge_req_2968_symbol : Boolean;
          signal merge_ack_2969_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_477_complete_2942_start <= ptr_deref_477_active_x_x2912_symbol; -- control passed to block
          Xentry_2943_symbol  <= ptr_deref_477_complete_2942_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/$entry
          word_access_2945: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access 
            signal word_access_2945_start: Boolean;
            signal Xentry_2946_symbol: Boolean;
            signal Xexit_2947_symbol: Boolean;
            signal word_access_0_2948_symbol : Boolean;
            signal word_access_1_2953_symbol : Boolean;
            signal word_access_2_2958_symbol : Boolean;
            signal word_access_3_2963_symbol : Boolean;
            -- 
          begin -- 
            word_access_2945_start <= Xentry_2943_symbol; -- control passed to block
            Xentry_2946_symbol  <= word_access_2945_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/$entry
            word_access_0_2948: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0 
              signal word_access_0_2948_start: Boolean;
              signal Xentry_2949_symbol: Boolean;
              signal Xexit_2950_symbol: Boolean;
              signal cr_2951_symbol : Boolean;
              signal ca_2952_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2948_start <= Xentry_2946_symbol; -- control passed to block
              Xentry_2949_symbol  <= word_access_0_2948_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/$entry
              cr_2951_symbol <= Xentry_2949_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/cr
              ptr_deref_477_load_0_req_1 <= cr_2951_symbol; -- link to DP
              ca_2952_symbol <= ptr_deref_477_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/ca
              Xexit_2950_symbol <= ca_2952_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/$exit
              word_access_0_2948_symbol <= Xexit_2950_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0
            word_access_1_2953: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_1 
              signal word_access_1_2953_start: Boolean;
              signal Xentry_2954_symbol: Boolean;
              signal Xexit_2955_symbol: Boolean;
              signal cr_2956_symbol : Boolean;
              signal ca_2957_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2953_start <= Xentry_2946_symbol; -- control passed to block
              Xentry_2954_symbol  <= word_access_1_2953_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_1/$entry
              cr_2956_symbol <= Xentry_2954_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_1/cr
              ptr_deref_477_load_1_req_1 <= cr_2956_symbol; -- link to DP
              ca_2957_symbol <= ptr_deref_477_load_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_1/ca
              Xexit_2955_symbol <= ca_2957_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_1/$exit
              word_access_1_2953_symbol <= Xexit_2955_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_1
            word_access_2_2958: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_2 
              signal word_access_2_2958_start: Boolean;
              signal Xentry_2959_symbol: Boolean;
              signal Xexit_2960_symbol: Boolean;
              signal cr_2961_symbol : Boolean;
              signal ca_2962_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2958_start <= Xentry_2946_symbol; -- control passed to block
              Xentry_2959_symbol  <= word_access_2_2958_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_2/$entry
              cr_2961_symbol <= Xentry_2959_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_2/cr
              ptr_deref_477_load_2_req_1 <= cr_2961_symbol; -- link to DP
              ca_2962_symbol <= ptr_deref_477_load_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_2/ca
              Xexit_2960_symbol <= ca_2962_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_2/$exit
              word_access_2_2958_symbol <= Xexit_2960_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_2
            word_access_3_2963: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_3 
              signal word_access_3_2963_start: Boolean;
              signal Xentry_2964_symbol: Boolean;
              signal Xexit_2965_symbol: Boolean;
              signal cr_2966_symbol : Boolean;
              signal ca_2967_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2963_start <= Xentry_2946_symbol; -- control passed to block
              Xentry_2964_symbol  <= word_access_3_2963_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_3/$entry
              cr_2966_symbol <= Xentry_2964_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_3/cr
              ptr_deref_477_load_3_req_1 <= cr_2966_symbol; -- link to DP
              ca_2967_symbol <= ptr_deref_477_load_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_3/ca
              Xexit_2965_symbol <= ca_2967_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_3/$exit
              word_access_3_2963_symbol <= Xexit_2965_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_3
            Xexit_2947_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/$exit 
              signal Xexit_2947_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2947_predecessors(0) <= word_access_0_2948_symbol;
              Xexit_2947_predecessors(1) <= word_access_1_2953_symbol;
              Xexit_2947_predecessors(2) <= word_access_2_2958_symbol;
              Xexit_2947_predecessors(3) <= word_access_3_2963_symbol;
              Xexit_2947_join: join -- 
                port map( -- 
                  preds => Xexit_2947_predecessors,
                  symbol_out => Xexit_2947_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/$exit
            word_access_2945_symbol <= Xexit_2947_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access
          merge_req_2968_symbol <= word_access_2945_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/merge_req
          ptr_deref_477_gather_scatter_req_0 <= merge_req_2968_symbol; -- link to DP
          merge_ack_2969_symbol <= ptr_deref_477_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/merge_ack
          Xexit_2944_symbol <= merge_ack_2969_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/$exit
          ptr_deref_477_complete_2942_symbol <= Xexit_2944_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete
        assign_stmt_482_active_x_x2970_symbol <= ptr_deref_481_complete_3003_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_482_active_
        assign_stmt_482_completed_x_x2971_symbol <= assign_stmt_482_active_x_x2970_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_482_completed_
        ptr_deref_481_trigger_x_x2972_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_trigger_ 
          signal ptr_deref_481_trigger_x_x2972_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_481_trigger_x_x2972_predecessors(0) <= ptr_deref_481_word_address_calculated_2976_symbol;
          ptr_deref_481_trigger_x_x2972_predecessors(1) <= ptr_deref_472_active_x_x2851_symbol;
          ptr_deref_481_trigger_x_x2972_join: join -- 
            port map( -- 
              preds => ptr_deref_481_trigger_x_x2972_predecessors,
              symbol_out => ptr_deref_481_trigger_x_x2972_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_trigger_
        ptr_deref_481_active_x_x2973_symbol <= ptr_deref_481_request_2977_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_active_
        ptr_deref_481_base_address_calculated_2974_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_base_address_calculated
        ptr_deref_481_root_address_calculated_2975_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_root_address_calculated
        ptr_deref_481_word_address_calculated_2976_symbol <= ptr_deref_481_root_address_calculated_2975_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_word_address_calculated
        ptr_deref_481_request_2977: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request 
          signal ptr_deref_481_request_2977_start: Boolean;
          signal Xentry_2978_symbol: Boolean;
          signal Xexit_2979_symbol: Boolean;
          signal word_access_2980_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_481_request_2977_start <= ptr_deref_481_trigger_x_x2972_symbol; -- control passed to block
          Xentry_2978_symbol  <= ptr_deref_481_request_2977_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/$entry
          word_access_2980: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access 
            signal word_access_2980_start: Boolean;
            signal Xentry_2981_symbol: Boolean;
            signal Xexit_2982_symbol: Boolean;
            signal word_access_0_2983_symbol : Boolean;
            signal word_access_1_2988_symbol : Boolean;
            signal word_access_2_2993_symbol : Boolean;
            signal word_access_3_2998_symbol : Boolean;
            -- 
          begin -- 
            word_access_2980_start <= Xentry_2978_symbol; -- control passed to block
            Xentry_2981_symbol  <= word_access_2980_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/$entry
            word_access_0_2983: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0 
              signal word_access_0_2983_start: Boolean;
              signal Xentry_2984_symbol: Boolean;
              signal Xexit_2985_symbol: Boolean;
              signal rr_2986_symbol : Boolean;
              signal ra_2987_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2983_start <= Xentry_2981_symbol; -- control passed to block
              Xentry_2984_symbol  <= word_access_0_2983_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/$entry
              rr_2986_symbol <= Xentry_2984_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/rr
              ptr_deref_481_load_0_req_0 <= rr_2986_symbol; -- link to DP
              ra_2987_symbol <= ptr_deref_481_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/ra
              Xexit_2985_symbol <= ra_2987_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/$exit
              word_access_0_2983_symbol <= Xexit_2985_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0
            word_access_1_2988: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_1 
              signal word_access_1_2988_start: Boolean;
              signal Xentry_2989_symbol: Boolean;
              signal Xexit_2990_symbol: Boolean;
              signal rr_2991_symbol : Boolean;
              signal ra_2992_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_2988_start <= Xentry_2981_symbol; -- control passed to block
              Xentry_2989_symbol  <= word_access_1_2988_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_1/$entry
              rr_2991_symbol <= Xentry_2989_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_1/rr
              ptr_deref_481_load_1_req_0 <= rr_2991_symbol; -- link to DP
              ra_2992_symbol <= ptr_deref_481_load_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_1/ra
              Xexit_2990_symbol <= ra_2992_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_1/$exit
              word_access_1_2988_symbol <= Xexit_2990_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_1
            word_access_2_2993: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_2 
              signal word_access_2_2993_start: Boolean;
              signal Xentry_2994_symbol: Boolean;
              signal Xexit_2995_symbol: Boolean;
              signal rr_2996_symbol : Boolean;
              signal ra_2997_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_2993_start <= Xentry_2981_symbol; -- control passed to block
              Xentry_2994_symbol  <= word_access_2_2993_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_2/$entry
              rr_2996_symbol <= Xentry_2994_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_2/rr
              ptr_deref_481_load_2_req_0 <= rr_2996_symbol; -- link to DP
              ra_2997_symbol <= ptr_deref_481_load_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_2/ra
              Xexit_2995_symbol <= ra_2997_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_2/$exit
              word_access_2_2993_symbol <= Xexit_2995_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_2
            word_access_3_2998: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_3 
              signal word_access_3_2998_start: Boolean;
              signal Xentry_2999_symbol: Boolean;
              signal Xexit_3000_symbol: Boolean;
              signal rr_3001_symbol : Boolean;
              signal ra_3002_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_2998_start <= Xentry_2981_symbol; -- control passed to block
              Xentry_2999_symbol  <= word_access_3_2998_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_3/$entry
              rr_3001_symbol <= Xentry_2999_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_3/rr
              ptr_deref_481_load_3_req_0 <= rr_3001_symbol; -- link to DP
              ra_3002_symbol <= ptr_deref_481_load_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_3/ra
              Xexit_3000_symbol <= ra_3002_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_3/$exit
              word_access_3_2998_symbol <= Xexit_3000_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_3
            Xexit_2982_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/$exit 
              signal Xexit_2982_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_2982_predecessors(0) <= word_access_0_2983_symbol;
              Xexit_2982_predecessors(1) <= word_access_1_2988_symbol;
              Xexit_2982_predecessors(2) <= word_access_2_2993_symbol;
              Xexit_2982_predecessors(3) <= word_access_3_2998_symbol;
              Xexit_2982_join: join -- 
                port map( -- 
                  preds => Xexit_2982_predecessors,
                  symbol_out => Xexit_2982_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/$exit
            word_access_2980_symbol <= Xexit_2982_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access
          Xexit_2979_symbol <= word_access_2980_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/$exit
          ptr_deref_481_request_2977_symbol <= Xexit_2979_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request
        ptr_deref_481_complete_3003: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete 
          signal ptr_deref_481_complete_3003_start: Boolean;
          signal Xentry_3004_symbol: Boolean;
          signal Xexit_3005_symbol: Boolean;
          signal word_access_3006_symbol : Boolean;
          signal merge_req_3029_symbol : Boolean;
          signal merge_ack_3030_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_481_complete_3003_start <= ptr_deref_481_active_x_x2973_symbol; -- control passed to block
          Xentry_3004_symbol  <= ptr_deref_481_complete_3003_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/$entry
          word_access_3006: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access 
            signal word_access_3006_start: Boolean;
            signal Xentry_3007_symbol: Boolean;
            signal Xexit_3008_symbol: Boolean;
            signal word_access_0_3009_symbol : Boolean;
            signal word_access_1_3014_symbol : Boolean;
            signal word_access_2_3019_symbol : Boolean;
            signal word_access_3_3024_symbol : Boolean;
            -- 
          begin -- 
            word_access_3006_start <= Xentry_3004_symbol; -- control passed to block
            Xentry_3007_symbol  <= word_access_3006_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/$entry
            word_access_0_3009: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0 
              signal word_access_0_3009_start: Boolean;
              signal Xentry_3010_symbol: Boolean;
              signal Xexit_3011_symbol: Boolean;
              signal cr_3012_symbol : Boolean;
              signal ca_3013_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3009_start <= Xentry_3007_symbol; -- control passed to block
              Xentry_3010_symbol  <= word_access_0_3009_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/$entry
              cr_3012_symbol <= Xentry_3010_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/cr
              ptr_deref_481_load_0_req_1 <= cr_3012_symbol; -- link to DP
              ca_3013_symbol <= ptr_deref_481_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/ca
              Xexit_3011_symbol <= ca_3013_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/$exit
              word_access_0_3009_symbol <= Xexit_3011_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0
            word_access_1_3014: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_1 
              signal word_access_1_3014_start: Boolean;
              signal Xentry_3015_symbol: Boolean;
              signal Xexit_3016_symbol: Boolean;
              signal cr_3017_symbol : Boolean;
              signal ca_3018_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3014_start <= Xentry_3007_symbol; -- control passed to block
              Xentry_3015_symbol  <= word_access_1_3014_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_1/$entry
              cr_3017_symbol <= Xentry_3015_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_1/cr
              ptr_deref_481_load_1_req_1 <= cr_3017_symbol; -- link to DP
              ca_3018_symbol <= ptr_deref_481_load_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_1/ca
              Xexit_3016_symbol <= ca_3018_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_1/$exit
              word_access_1_3014_symbol <= Xexit_3016_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_1
            word_access_2_3019: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_2 
              signal word_access_2_3019_start: Boolean;
              signal Xentry_3020_symbol: Boolean;
              signal Xexit_3021_symbol: Boolean;
              signal cr_3022_symbol : Boolean;
              signal ca_3023_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3019_start <= Xentry_3007_symbol; -- control passed to block
              Xentry_3020_symbol  <= word_access_2_3019_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_2/$entry
              cr_3022_symbol <= Xentry_3020_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_2/cr
              ptr_deref_481_load_2_req_1 <= cr_3022_symbol; -- link to DP
              ca_3023_symbol <= ptr_deref_481_load_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_2/ca
              Xexit_3021_symbol <= ca_3023_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_2/$exit
              word_access_2_3019_symbol <= Xexit_3021_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_2
            word_access_3_3024: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_3 
              signal word_access_3_3024_start: Boolean;
              signal Xentry_3025_symbol: Boolean;
              signal Xexit_3026_symbol: Boolean;
              signal cr_3027_symbol : Boolean;
              signal ca_3028_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3024_start <= Xentry_3007_symbol; -- control passed to block
              Xentry_3025_symbol  <= word_access_3_3024_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_3/$entry
              cr_3027_symbol <= Xentry_3025_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_3/cr
              ptr_deref_481_load_3_req_1 <= cr_3027_symbol; -- link to DP
              ca_3028_symbol <= ptr_deref_481_load_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_3/ca
              Xexit_3026_symbol <= ca_3028_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_3/$exit
              word_access_3_3024_symbol <= Xexit_3026_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_3
            Xexit_3008_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/$exit 
              signal Xexit_3008_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3008_predecessors(0) <= word_access_0_3009_symbol;
              Xexit_3008_predecessors(1) <= word_access_1_3014_symbol;
              Xexit_3008_predecessors(2) <= word_access_2_3019_symbol;
              Xexit_3008_predecessors(3) <= word_access_3_3024_symbol;
              Xexit_3008_join: join -- 
                port map( -- 
                  preds => Xexit_3008_predecessors,
                  symbol_out => Xexit_3008_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/$exit
            word_access_3006_symbol <= Xexit_3008_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access
          merge_req_3029_symbol <= word_access_3006_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/merge_req
          ptr_deref_481_gather_scatter_req_0 <= merge_req_3029_symbol; -- link to DP
          merge_ack_3030_symbol <= ptr_deref_481_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/merge_ack
          Xexit_3005_symbol <= merge_ack_3030_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/$exit
          ptr_deref_481_complete_3003_symbol <= Xexit_3005_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete
        assign_stmt_487_active_x_x3031_symbol <= array_obj_ref_486_complete_3051_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_487_active_
        assign_stmt_487_completed_x_x3032_symbol <= assign_stmt_487_active_x_x3031_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_487_completed_
        array_obj_ref_486_trigger_x_x3033_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_trigger_
        array_obj_ref_486_active_x_x3034_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_active_ 
          signal array_obj_ref_486_active_x_x3034_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_486_active_x_x3034_predecessors(0) <= array_obj_ref_486_trigger_x_x3033_symbol;
          array_obj_ref_486_active_x_x3034_predecessors(1) <= array_obj_ref_486_root_address_calculated_3036_symbol;
          array_obj_ref_486_active_x_x3034_join: join -- 
            port map( -- 
              preds => array_obj_ref_486_active_x_x3034_predecessors,
              symbol_out => array_obj_ref_486_active_x_x3034_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_active_
        array_obj_ref_486_base_address_calculated_3035_symbol <= assign_stmt_482_completed_x_x2971_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_address_calculated
        array_obj_ref_486_root_address_calculated_3036_symbol <= array_obj_ref_486_base_plus_offset_3044_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_root_address_calculated
        array_obj_ref_486_base_address_resized_3037_symbol <= array_obj_ref_486_base_addr_resize_3038_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_address_resized
        array_obj_ref_486_base_addr_resize_3038: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize 
          signal array_obj_ref_486_base_addr_resize_3038_start: Boolean;
          signal Xentry_3039_symbol: Boolean;
          signal Xexit_3040_symbol: Boolean;
          signal base_resize_req_3041_symbol : Boolean;
          signal base_resize_ack_3042_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_486_base_addr_resize_3038_start <= array_obj_ref_486_base_address_calculated_3035_symbol; -- control passed to block
          Xentry_3039_symbol  <= array_obj_ref_486_base_addr_resize_3038_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/$entry
          base_resize_req_3041_symbol <= Xentry_3039_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/base_resize_req
          array_obj_ref_486_base_resize_req_0 <= base_resize_req_3041_symbol; -- link to DP
          base_resize_ack_3042_symbol <= array_obj_ref_486_base_resize_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/base_resize_ack
          Xexit_3040_symbol <= base_resize_ack_3042_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/$exit
          array_obj_ref_486_base_addr_resize_3038_symbol <= Xexit_3040_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize
        array_obj_ref_486_base_plus_offset_trigger_3043_symbol <= array_obj_ref_486_base_address_resized_3037_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset_trigger
        array_obj_ref_486_base_plus_offset_3044: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset 
          signal array_obj_ref_486_base_plus_offset_3044_start: Boolean;
          signal Xentry_3045_symbol: Boolean;
          signal Xexit_3046_symbol: Boolean;
          signal plus_base_rr_3047_symbol : Boolean;
          signal plus_base_ra_3048_symbol : Boolean;
          signal plus_base_cr_3049_symbol : Boolean;
          signal plus_base_ca_3050_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_486_base_plus_offset_3044_start <= array_obj_ref_486_base_plus_offset_trigger_3043_symbol; -- control passed to block
          Xentry_3045_symbol  <= array_obj_ref_486_base_plus_offset_3044_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/$entry
          plus_base_rr_3047_symbol <= Xentry_3045_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_rr
          array_obj_ref_486_root_address_inst_req_0 <= plus_base_rr_3047_symbol; -- link to DP
          plus_base_ra_3048_symbol <= array_obj_ref_486_root_address_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_ra
          plus_base_cr_3049_symbol <= plus_base_ra_3048_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_cr
          array_obj_ref_486_root_address_inst_req_1 <= plus_base_cr_3049_symbol; -- link to DP
          plus_base_ca_3050_symbol <= array_obj_ref_486_root_address_inst_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_ca
          Xexit_3046_symbol <= plus_base_ca_3050_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/$exit
          array_obj_ref_486_base_plus_offset_3044_symbol <= Xexit_3046_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset
        array_obj_ref_486_complete_3051: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete 
          signal array_obj_ref_486_complete_3051_start: Boolean;
          signal Xentry_3052_symbol: Boolean;
          signal Xexit_3053_symbol: Boolean;
          signal final_reg_req_3054_symbol : Boolean;
          signal final_reg_ack_3055_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_486_complete_3051_start <= array_obj_ref_486_active_x_x3034_symbol; -- control passed to block
          Xentry_3052_symbol  <= array_obj_ref_486_complete_3051_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/$entry
          final_reg_req_3054_symbol <= Xentry_3052_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/final_reg_req
          array_obj_ref_486_final_reg_req_0 <= final_reg_req_3054_symbol; -- link to DP
          final_reg_ack_3055_symbol <= array_obj_ref_486_final_reg_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/final_reg_ack
          Xexit_3053_symbol <= final_reg_ack_3055_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/$exit
          array_obj_ref_486_complete_3051_symbol <= Xexit_3053_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete
        assign_stmt_491_active_x_x3056_symbol <= simple_obj_ref_490_complete_3058_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_491_active_
        assign_stmt_491_completed_x_x3057_symbol <= ptr_deref_489_complete_3135_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_491_completed_
        simple_obj_ref_490_complete_3058_symbol <= assign_stmt_478_completed_x_x2910_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_490_complete
        ptr_deref_489_trigger_x_x3059_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_trigger_ 
          signal ptr_deref_489_trigger_x_x3059_predecessors: BooleanArray(4 downto 0);
          -- 
        begin -- 
          ptr_deref_489_trigger_x_x3059_predecessors(0) <= ptr_deref_489_word_address_calculated_3064_symbol;
          ptr_deref_489_trigger_x_x3059_predecessors(1) <= ptr_deref_489_base_address_calculated_3061_symbol;
          ptr_deref_489_trigger_x_x3059_predecessors(2) <= assign_stmt_491_active_x_x3056_symbol;
          ptr_deref_489_trigger_x_x3059_predecessors(3) <= ptr_deref_477_active_x_x2912_symbol;
          ptr_deref_489_trigger_x_x3059_predecessors(4) <= ptr_deref_481_active_x_x2973_symbol;
          ptr_deref_489_trigger_x_x3059_join: join -- 
            port map( -- 
              preds => ptr_deref_489_trigger_x_x3059_predecessors,
              symbol_out => ptr_deref_489_trigger_x_x3059_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_trigger_
        ptr_deref_489_active_x_x3060_symbol <= ptr_deref_489_request_3107_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_active_
        ptr_deref_489_base_address_calculated_3061_symbol <= simple_obj_ref_488_complete_3062_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_address_calculated
        simple_obj_ref_488_complete_3062_symbol <= assign_stmt_487_completed_x_x3032_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_488_complete
        ptr_deref_489_root_address_calculated_3063_symbol <= ptr_deref_489_base_plus_offset_3071_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_root_address_calculated
        ptr_deref_489_word_address_calculated_3064_symbol <= ptr_deref_489_word_addrgen_3076_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_address_calculated
        ptr_deref_489_base_address_resized_3065_symbol <= ptr_deref_489_base_addr_resize_3066_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_address_resized
        ptr_deref_489_base_addr_resize_3066: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize 
          signal ptr_deref_489_base_addr_resize_3066_start: Boolean;
          signal Xentry_3067_symbol: Boolean;
          signal Xexit_3068_symbol: Boolean;
          signal base_resize_req_3069_symbol : Boolean;
          signal base_resize_ack_3070_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_base_addr_resize_3066_start <= ptr_deref_489_base_address_calculated_3061_symbol; -- control passed to block
          Xentry_3067_symbol  <= ptr_deref_489_base_addr_resize_3066_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/$entry
          base_resize_req_3069_symbol <= Xentry_3067_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/base_resize_req
          ptr_deref_489_base_resize_req_0 <= base_resize_req_3069_symbol; -- link to DP
          base_resize_ack_3070_symbol <= ptr_deref_489_base_resize_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/base_resize_ack
          Xexit_3068_symbol <= base_resize_ack_3070_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/$exit
          ptr_deref_489_base_addr_resize_3066_symbol <= Xexit_3068_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize
        ptr_deref_489_base_plus_offset_3071: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset 
          signal ptr_deref_489_base_plus_offset_3071_start: Boolean;
          signal Xentry_3072_symbol: Boolean;
          signal Xexit_3073_symbol: Boolean;
          signal sum_rename_req_3074_symbol : Boolean;
          signal sum_rename_ack_3075_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_base_plus_offset_3071_start <= ptr_deref_489_base_address_resized_3065_symbol; -- control passed to block
          Xentry_3072_symbol  <= ptr_deref_489_base_plus_offset_3071_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/$entry
          sum_rename_req_3074_symbol <= Xentry_3072_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/sum_rename_req
          ptr_deref_489_root_address_inst_req_0 <= sum_rename_req_3074_symbol; -- link to DP
          sum_rename_ack_3075_symbol <= ptr_deref_489_root_address_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/sum_rename_ack
          Xexit_3073_symbol <= sum_rename_ack_3075_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/$exit
          ptr_deref_489_base_plus_offset_3071_symbol <= Xexit_3073_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset
        ptr_deref_489_word_addrgen_3076: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen 
          signal ptr_deref_489_word_addrgen_3076_start: Boolean;
          signal Xentry_3077_symbol: Boolean;
          signal Xexit_3078_symbol: Boolean;
          signal word_0_3079_symbol : Boolean;
          signal word_1_3086_symbol : Boolean;
          signal word_2_3093_symbol : Boolean;
          signal word_3_3100_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_word_addrgen_3076_start <= ptr_deref_489_root_address_calculated_3063_symbol; -- control passed to block
          Xentry_3077_symbol  <= ptr_deref_489_word_addrgen_3076_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/$entry
          word_0_3079: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0 
            signal word_0_3079_start: Boolean;
            signal Xentry_3080_symbol: Boolean;
            signal Xexit_3081_symbol: Boolean;
            signal rr_3082_symbol : Boolean;
            signal ra_3083_symbol : Boolean;
            signal cr_3084_symbol : Boolean;
            signal ca_3085_symbol : Boolean;
            -- 
          begin -- 
            word_0_3079_start <= Xentry_3077_symbol; -- control passed to block
            Xentry_3080_symbol  <= word_0_3079_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0/$entry
            rr_3082_symbol <= Xentry_3080_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0/rr
            ptr_deref_489_addr_0_req_0 <= rr_3082_symbol; -- link to DP
            ra_3083_symbol <= ptr_deref_489_addr_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0/ra
            cr_3084_symbol <= ra_3083_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0/cr
            ptr_deref_489_addr_0_req_1 <= cr_3084_symbol; -- link to DP
            ca_3085_symbol <= ptr_deref_489_addr_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0/ca
            Xexit_3081_symbol <= ca_3085_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0/$exit
            word_0_3079_symbol <= Xexit_3081_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_0
          word_1_3086: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1 
            signal word_1_3086_start: Boolean;
            signal Xentry_3087_symbol: Boolean;
            signal Xexit_3088_symbol: Boolean;
            signal rr_3089_symbol : Boolean;
            signal ra_3090_symbol : Boolean;
            signal cr_3091_symbol : Boolean;
            signal ca_3092_symbol : Boolean;
            -- 
          begin -- 
            word_1_3086_start <= Xentry_3077_symbol; -- control passed to block
            Xentry_3087_symbol  <= word_1_3086_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1/$entry
            rr_3089_symbol <= Xentry_3087_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1/rr
            ptr_deref_489_addr_1_req_0 <= rr_3089_symbol; -- link to DP
            ra_3090_symbol <= ptr_deref_489_addr_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1/ra
            cr_3091_symbol <= ra_3090_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1/cr
            ptr_deref_489_addr_1_req_1 <= cr_3091_symbol; -- link to DP
            ca_3092_symbol <= ptr_deref_489_addr_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1/ca
            Xexit_3088_symbol <= ca_3092_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1/$exit
            word_1_3086_symbol <= Xexit_3088_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_1
          word_2_3093: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2 
            signal word_2_3093_start: Boolean;
            signal Xentry_3094_symbol: Boolean;
            signal Xexit_3095_symbol: Boolean;
            signal rr_3096_symbol : Boolean;
            signal ra_3097_symbol : Boolean;
            signal cr_3098_symbol : Boolean;
            signal ca_3099_symbol : Boolean;
            -- 
          begin -- 
            word_2_3093_start <= Xentry_3077_symbol; -- control passed to block
            Xentry_3094_symbol  <= word_2_3093_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2/$entry
            rr_3096_symbol <= Xentry_3094_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2/rr
            ptr_deref_489_addr_2_req_0 <= rr_3096_symbol; -- link to DP
            ra_3097_symbol <= ptr_deref_489_addr_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2/ra
            cr_3098_symbol <= ra_3097_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2/cr
            ptr_deref_489_addr_2_req_1 <= cr_3098_symbol; -- link to DP
            ca_3099_symbol <= ptr_deref_489_addr_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2/ca
            Xexit_3095_symbol <= ca_3099_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2/$exit
            word_2_3093_symbol <= Xexit_3095_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_2
          word_3_3100: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3 
            signal word_3_3100_start: Boolean;
            signal Xentry_3101_symbol: Boolean;
            signal Xexit_3102_symbol: Boolean;
            signal rr_3103_symbol : Boolean;
            signal ra_3104_symbol : Boolean;
            signal cr_3105_symbol : Boolean;
            signal ca_3106_symbol : Boolean;
            -- 
          begin -- 
            word_3_3100_start <= Xentry_3077_symbol; -- control passed to block
            Xentry_3101_symbol  <= word_3_3100_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3/$entry
            rr_3103_symbol <= Xentry_3101_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3/rr
            ptr_deref_489_addr_3_req_0 <= rr_3103_symbol; -- link to DP
            ra_3104_symbol <= ptr_deref_489_addr_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3/ra
            cr_3105_symbol <= ra_3104_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3/cr
            ptr_deref_489_addr_3_req_1 <= cr_3105_symbol; -- link to DP
            ca_3106_symbol <= ptr_deref_489_addr_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3/ca
            Xexit_3102_symbol <= ca_3106_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3/$exit
            word_3_3100_symbol <= Xexit_3102_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/word_3
          Xexit_3078_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/$exit 
            signal Xexit_3078_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_3078_predecessors(0) <= word_0_3079_symbol;
            Xexit_3078_predecessors(1) <= word_1_3086_symbol;
            Xexit_3078_predecessors(2) <= word_2_3093_symbol;
            Xexit_3078_predecessors(3) <= word_3_3100_symbol;
            Xexit_3078_join: join -- 
              port map( -- 
                preds => Xexit_3078_predecessors,
                symbol_out => Xexit_3078_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/$exit
          ptr_deref_489_word_addrgen_3076_symbol <= Xexit_3078_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen
        ptr_deref_489_request_3107: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request 
          signal ptr_deref_489_request_3107_start: Boolean;
          signal Xentry_3108_symbol: Boolean;
          signal Xexit_3109_symbol: Boolean;
          signal split_req_3110_symbol : Boolean;
          signal split_ack_3111_symbol : Boolean;
          signal word_access_3112_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_request_3107_start <= ptr_deref_489_trigger_x_x3059_symbol; -- control passed to block
          Xentry_3108_symbol  <= ptr_deref_489_request_3107_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/$entry
          split_req_3110_symbol <= Xentry_3108_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/split_req
          ptr_deref_489_gather_scatter_req_0 <= split_req_3110_symbol; -- link to DP
          split_ack_3111_symbol <= ptr_deref_489_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/split_ack
          word_access_3112: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access 
            signal word_access_3112_start: Boolean;
            signal Xentry_3113_symbol: Boolean;
            signal Xexit_3114_symbol: Boolean;
            signal word_access_0_3115_symbol : Boolean;
            signal word_access_1_3120_symbol : Boolean;
            signal word_access_2_3125_symbol : Boolean;
            signal word_access_3_3130_symbol : Boolean;
            -- 
          begin -- 
            word_access_3112_start <= split_ack_3111_symbol; -- control passed to block
            Xentry_3113_symbol  <= word_access_3112_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/$entry
            word_access_0_3115: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0 
              signal word_access_0_3115_start: Boolean;
              signal Xentry_3116_symbol: Boolean;
              signal Xexit_3117_symbol: Boolean;
              signal rr_3118_symbol : Boolean;
              signal ra_3119_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3115_start <= Xentry_3113_symbol; -- control passed to block
              Xentry_3116_symbol  <= word_access_0_3115_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/$entry
              rr_3118_symbol <= Xentry_3116_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/rr
              ptr_deref_489_store_0_req_0 <= rr_3118_symbol; -- link to DP
              ra_3119_symbol <= ptr_deref_489_store_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/ra
              Xexit_3117_symbol <= ra_3119_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/$exit
              word_access_0_3115_symbol <= Xexit_3117_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0
            word_access_1_3120: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_1 
              signal word_access_1_3120_start: Boolean;
              signal Xentry_3121_symbol: Boolean;
              signal Xexit_3122_symbol: Boolean;
              signal rr_3123_symbol : Boolean;
              signal ra_3124_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3120_start <= Xentry_3113_symbol; -- control passed to block
              Xentry_3121_symbol  <= word_access_1_3120_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_1/$entry
              rr_3123_symbol <= Xentry_3121_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_1/rr
              ptr_deref_489_store_1_req_0 <= rr_3123_symbol; -- link to DP
              ra_3124_symbol <= ptr_deref_489_store_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_1/ra
              Xexit_3122_symbol <= ra_3124_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_1/$exit
              word_access_1_3120_symbol <= Xexit_3122_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_1
            word_access_2_3125: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_2 
              signal word_access_2_3125_start: Boolean;
              signal Xentry_3126_symbol: Boolean;
              signal Xexit_3127_symbol: Boolean;
              signal rr_3128_symbol : Boolean;
              signal ra_3129_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3125_start <= Xentry_3113_symbol; -- control passed to block
              Xentry_3126_symbol  <= word_access_2_3125_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_2/$entry
              rr_3128_symbol <= Xentry_3126_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_2/rr
              ptr_deref_489_store_2_req_0 <= rr_3128_symbol; -- link to DP
              ra_3129_symbol <= ptr_deref_489_store_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_2/ra
              Xexit_3127_symbol <= ra_3129_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_2/$exit
              word_access_2_3125_symbol <= Xexit_3127_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_2
            word_access_3_3130: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_3 
              signal word_access_3_3130_start: Boolean;
              signal Xentry_3131_symbol: Boolean;
              signal Xexit_3132_symbol: Boolean;
              signal rr_3133_symbol : Boolean;
              signal ra_3134_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3130_start <= Xentry_3113_symbol; -- control passed to block
              Xentry_3131_symbol  <= word_access_3_3130_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_3/$entry
              rr_3133_symbol <= Xentry_3131_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_3/rr
              ptr_deref_489_store_3_req_0 <= rr_3133_symbol; -- link to DP
              ra_3134_symbol <= ptr_deref_489_store_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_3/ra
              Xexit_3132_symbol <= ra_3134_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_3/$exit
              word_access_3_3130_symbol <= Xexit_3132_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_3
            Xexit_3114_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/$exit 
              signal Xexit_3114_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3114_predecessors(0) <= word_access_0_3115_symbol;
              Xexit_3114_predecessors(1) <= word_access_1_3120_symbol;
              Xexit_3114_predecessors(2) <= word_access_2_3125_symbol;
              Xexit_3114_predecessors(3) <= word_access_3_3130_symbol;
              Xexit_3114_join: join -- 
                port map( -- 
                  preds => Xexit_3114_predecessors,
                  symbol_out => Xexit_3114_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/$exit
            word_access_3112_symbol <= Xexit_3114_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access
          Xexit_3109_symbol <= word_access_3112_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/$exit
          ptr_deref_489_request_3107_symbol <= Xexit_3109_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request
        ptr_deref_489_complete_3135: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete 
          signal ptr_deref_489_complete_3135_start: Boolean;
          signal Xentry_3136_symbol: Boolean;
          signal Xexit_3137_symbol: Boolean;
          signal word_access_3138_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_complete_3135_start <= ptr_deref_489_active_x_x3060_symbol; -- control passed to block
          Xentry_3136_symbol  <= ptr_deref_489_complete_3135_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/$entry
          word_access_3138: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access 
            signal word_access_3138_start: Boolean;
            signal Xentry_3139_symbol: Boolean;
            signal Xexit_3140_symbol: Boolean;
            signal word_access_0_3141_symbol : Boolean;
            signal word_access_1_3146_symbol : Boolean;
            signal word_access_2_3151_symbol : Boolean;
            signal word_access_3_3156_symbol : Boolean;
            -- 
          begin -- 
            word_access_3138_start <= Xentry_3136_symbol; -- control passed to block
            Xentry_3139_symbol  <= word_access_3138_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/$entry
            word_access_0_3141: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0 
              signal word_access_0_3141_start: Boolean;
              signal Xentry_3142_symbol: Boolean;
              signal Xexit_3143_symbol: Boolean;
              signal cr_3144_symbol : Boolean;
              signal ca_3145_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3141_start <= Xentry_3139_symbol; -- control passed to block
              Xentry_3142_symbol  <= word_access_0_3141_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/$entry
              cr_3144_symbol <= Xentry_3142_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/cr
              ptr_deref_489_store_0_req_1 <= cr_3144_symbol; -- link to DP
              ca_3145_symbol <= ptr_deref_489_store_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/ca
              Xexit_3143_symbol <= ca_3145_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/$exit
              word_access_0_3141_symbol <= Xexit_3143_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0
            word_access_1_3146: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_1 
              signal word_access_1_3146_start: Boolean;
              signal Xentry_3147_symbol: Boolean;
              signal Xexit_3148_symbol: Boolean;
              signal cr_3149_symbol : Boolean;
              signal ca_3150_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3146_start <= Xentry_3139_symbol; -- control passed to block
              Xentry_3147_symbol  <= word_access_1_3146_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_1/$entry
              cr_3149_symbol <= Xentry_3147_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_1/cr
              ptr_deref_489_store_1_req_1 <= cr_3149_symbol; -- link to DP
              ca_3150_symbol <= ptr_deref_489_store_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_1/ca
              Xexit_3148_symbol <= ca_3150_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_1/$exit
              word_access_1_3146_symbol <= Xexit_3148_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_1
            word_access_2_3151: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_2 
              signal word_access_2_3151_start: Boolean;
              signal Xentry_3152_symbol: Boolean;
              signal Xexit_3153_symbol: Boolean;
              signal cr_3154_symbol : Boolean;
              signal ca_3155_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3151_start <= Xentry_3139_symbol; -- control passed to block
              Xentry_3152_symbol  <= word_access_2_3151_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_2/$entry
              cr_3154_symbol <= Xentry_3152_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_2/cr
              ptr_deref_489_store_2_req_1 <= cr_3154_symbol; -- link to DP
              ca_3155_symbol <= ptr_deref_489_store_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_2/ca
              Xexit_3153_symbol <= ca_3155_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_2/$exit
              word_access_2_3151_symbol <= Xexit_3153_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_2
            word_access_3_3156: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_3 
              signal word_access_3_3156_start: Boolean;
              signal Xentry_3157_symbol: Boolean;
              signal Xexit_3158_symbol: Boolean;
              signal cr_3159_symbol : Boolean;
              signal ca_3160_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3156_start <= Xentry_3139_symbol; -- control passed to block
              Xentry_3157_symbol  <= word_access_3_3156_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_3/$entry
              cr_3159_symbol <= Xentry_3157_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_3/cr
              ptr_deref_489_store_3_req_1 <= cr_3159_symbol; -- link to DP
              ca_3160_symbol <= ptr_deref_489_store_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_3/ca
              Xexit_3158_symbol <= ca_3160_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_3/$exit
              word_access_3_3156_symbol <= Xexit_3158_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_3
            Xexit_3140_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/$exit 
              signal Xexit_3140_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3140_predecessors(0) <= word_access_0_3141_symbol;
              Xexit_3140_predecessors(1) <= word_access_1_3146_symbol;
              Xexit_3140_predecessors(2) <= word_access_2_3151_symbol;
              Xexit_3140_predecessors(3) <= word_access_3_3156_symbol;
              Xexit_3140_join: join -- 
                port map( -- 
                  preds => Xexit_3140_predecessors,
                  symbol_out => Xexit_3140_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/$exit
            word_access_3138_symbol <= Xexit_3140_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access
          Xexit_3137_symbol <= word_access_3138_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/$exit
          ptr_deref_489_complete_3135_symbol <= Xexit_3137_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete
        assign_stmt_495_active_x_x3161_symbol <= ptr_deref_494_complete_3194_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_495_active_
        assign_stmt_495_completed_x_x3162_symbol <= assign_stmt_495_active_x_x3161_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_495_completed_
        ptr_deref_494_trigger_x_x3163_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_trigger_ 
          signal ptr_deref_494_trigger_x_x3163_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_494_trigger_x_x3163_predecessors(0) <= ptr_deref_494_word_address_calculated_3167_symbol;
          ptr_deref_494_trigger_x_x3163_predecessors(1) <= ptr_deref_489_active_x_x3060_symbol;
          ptr_deref_494_trigger_x_x3163_join: join -- 
            port map( -- 
              preds => ptr_deref_494_trigger_x_x3163_predecessors,
              symbol_out => ptr_deref_494_trigger_x_x3163_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_trigger_
        ptr_deref_494_active_x_x3164_symbol <= ptr_deref_494_request_3168_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_active_
        ptr_deref_494_base_address_calculated_3165_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_base_address_calculated
        ptr_deref_494_root_address_calculated_3166_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_root_address_calculated
        ptr_deref_494_word_address_calculated_3167_symbol <= ptr_deref_494_root_address_calculated_3166_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_word_address_calculated
        ptr_deref_494_request_3168: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request 
          signal ptr_deref_494_request_3168_start: Boolean;
          signal Xentry_3169_symbol: Boolean;
          signal Xexit_3170_symbol: Boolean;
          signal word_access_3171_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_494_request_3168_start <= ptr_deref_494_trigger_x_x3163_symbol; -- control passed to block
          Xentry_3169_symbol  <= ptr_deref_494_request_3168_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/$entry
          word_access_3171: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access 
            signal word_access_3171_start: Boolean;
            signal Xentry_3172_symbol: Boolean;
            signal Xexit_3173_symbol: Boolean;
            signal word_access_0_3174_symbol : Boolean;
            signal word_access_1_3179_symbol : Boolean;
            signal word_access_2_3184_symbol : Boolean;
            signal word_access_3_3189_symbol : Boolean;
            -- 
          begin -- 
            word_access_3171_start <= Xentry_3169_symbol; -- control passed to block
            Xentry_3172_symbol  <= word_access_3171_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/$entry
            word_access_0_3174: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0 
              signal word_access_0_3174_start: Boolean;
              signal Xentry_3175_symbol: Boolean;
              signal Xexit_3176_symbol: Boolean;
              signal rr_3177_symbol : Boolean;
              signal ra_3178_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3174_start <= Xentry_3172_symbol; -- control passed to block
              Xentry_3175_symbol  <= word_access_0_3174_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/$entry
              rr_3177_symbol <= Xentry_3175_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/rr
              ptr_deref_494_load_0_req_0 <= rr_3177_symbol; -- link to DP
              ra_3178_symbol <= ptr_deref_494_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/ra
              Xexit_3176_symbol <= ra_3178_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/$exit
              word_access_0_3174_symbol <= Xexit_3176_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0
            word_access_1_3179: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_1 
              signal word_access_1_3179_start: Boolean;
              signal Xentry_3180_symbol: Boolean;
              signal Xexit_3181_symbol: Boolean;
              signal rr_3182_symbol : Boolean;
              signal ra_3183_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3179_start <= Xentry_3172_symbol; -- control passed to block
              Xentry_3180_symbol  <= word_access_1_3179_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_1/$entry
              rr_3182_symbol <= Xentry_3180_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_1/rr
              ptr_deref_494_load_1_req_0 <= rr_3182_symbol; -- link to DP
              ra_3183_symbol <= ptr_deref_494_load_1_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_1/ra
              Xexit_3181_symbol <= ra_3183_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_1/$exit
              word_access_1_3179_symbol <= Xexit_3181_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_1
            word_access_2_3184: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_2 
              signal word_access_2_3184_start: Boolean;
              signal Xentry_3185_symbol: Boolean;
              signal Xexit_3186_symbol: Boolean;
              signal rr_3187_symbol : Boolean;
              signal ra_3188_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3184_start <= Xentry_3172_symbol; -- control passed to block
              Xentry_3185_symbol  <= word_access_2_3184_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_2/$entry
              rr_3187_symbol <= Xentry_3185_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_2/rr
              ptr_deref_494_load_2_req_0 <= rr_3187_symbol; -- link to DP
              ra_3188_symbol <= ptr_deref_494_load_2_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_2/ra
              Xexit_3186_symbol <= ra_3188_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_2/$exit
              word_access_2_3184_symbol <= Xexit_3186_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_2
            word_access_3_3189: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_3 
              signal word_access_3_3189_start: Boolean;
              signal Xentry_3190_symbol: Boolean;
              signal Xexit_3191_symbol: Boolean;
              signal rr_3192_symbol : Boolean;
              signal ra_3193_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3189_start <= Xentry_3172_symbol; -- control passed to block
              Xentry_3190_symbol  <= word_access_3_3189_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_3/$entry
              rr_3192_symbol <= Xentry_3190_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_3/rr
              ptr_deref_494_load_3_req_0 <= rr_3192_symbol; -- link to DP
              ra_3193_symbol <= ptr_deref_494_load_3_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_3/ra
              Xexit_3191_symbol <= ra_3193_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_3/$exit
              word_access_3_3189_symbol <= Xexit_3191_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_3
            Xexit_3173_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/$exit 
              signal Xexit_3173_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3173_predecessors(0) <= word_access_0_3174_symbol;
              Xexit_3173_predecessors(1) <= word_access_1_3179_symbol;
              Xexit_3173_predecessors(2) <= word_access_2_3184_symbol;
              Xexit_3173_predecessors(3) <= word_access_3_3189_symbol;
              Xexit_3173_join: join -- 
                port map( -- 
                  preds => Xexit_3173_predecessors,
                  symbol_out => Xexit_3173_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/$exit
            word_access_3171_symbol <= Xexit_3173_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access
          Xexit_3170_symbol <= word_access_3171_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/$exit
          ptr_deref_494_request_3168_symbol <= Xexit_3170_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request
        ptr_deref_494_complete_3194: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete 
          signal ptr_deref_494_complete_3194_start: Boolean;
          signal Xentry_3195_symbol: Boolean;
          signal Xexit_3196_symbol: Boolean;
          signal word_access_3197_symbol : Boolean;
          signal merge_req_3220_symbol : Boolean;
          signal merge_ack_3221_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_494_complete_3194_start <= ptr_deref_494_active_x_x3164_symbol; -- control passed to block
          Xentry_3195_symbol  <= ptr_deref_494_complete_3194_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/$entry
          word_access_3197: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access 
            signal word_access_3197_start: Boolean;
            signal Xentry_3198_symbol: Boolean;
            signal Xexit_3199_symbol: Boolean;
            signal word_access_0_3200_symbol : Boolean;
            signal word_access_1_3205_symbol : Boolean;
            signal word_access_2_3210_symbol : Boolean;
            signal word_access_3_3215_symbol : Boolean;
            -- 
          begin -- 
            word_access_3197_start <= Xentry_3195_symbol; -- control passed to block
            Xentry_3198_symbol  <= word_access_3197_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/$entry
            word_access_0_3200: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0 
              signal word_access_0_3200_start: Boolean;
              signal Xentry_3201_symbol: Boolean;
              signal Xexit_3202_symbol: Boolean;
              signal cr_3203_symbol : Boolean;
              signal ca_3204_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3200_start <= Xentry_3198_symbol; -- control passed to block
              Xentry_3201_symbol  <= word_access_0_3200_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/$entry
              cr_3203_symbol <= Xentry_3201_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/cr
              ptr_deref_494_load_0_req_1 <= cr_3203_symbol; -- link to DP
              ca_3204_symbol <= ptr_deref_494_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/ca
              Xexit_3202_symbol <= ca_3204_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/$exit
              word_access_0_3200_symbol <= Xexit_3202_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0
            word_access_1_3205: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_1 
              signal word_access_1_3205_start: Boolean;
              signal Xentry_3206_symbol: Boolean;
              signal Xexit_3207_symbol: Boolean;
              signal cr_3208_symbol : Boolean;
              signal ca_3209_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3205_start <= Xentry_3198_symbol; -- control passed to block
              Xentry_3206_symbol  <= word_access_1_3205_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_1/$entry
              cr_3208_symbol <= Xentry_3206_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_1/cr
              ptr_deref_494_load_1_req_1 <= cr_3208_symbol; -- link to DP
              ca_3209_symbol <= ptr_deref_494_load_1_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_1/ca
              Xexit_3207_symbol <= ca_3209_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_1/$exit
              word_access_1_3205_symbol <= Xexit_3207_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_1
            word_access_2_3210: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_2 
              signal word_access_2_3210_start: Boolean;
              signal Xentry_3211_symbol: Boolean;
              signal Xexit_3212_symbol: Boolean;
              signal cr_3213_symbol : Boolean;
              signal ca_3214_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3210_start <= Xentry_3198_symbol; -- control passed to block
              Xentry_3211_symbol  <= word_access_2_3210_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_2/$entry
              cr_3213_symbol <= Xentry_3211_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_2/cr
              ptr_deref_494_load_2_req_1 <= cr_3213_symbol; -- link to DP
              ca_3214_symbol <= ptr_deref_494_load_2_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_2/ca
              Xexit_3212_symbol <= ca_3214_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_2/$exit
              word_access_2_3210_symbol <= Xexit_3212_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_2
            word_access_3_3215: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_3 
              signal word_access_3_3215_start: Boolean;
              signal Xentry_3216_symbol: Boolean;
              signal Xexit_3217_symbol: Boolean;
              signal cr_3218_symbol : Boolean;
              signal ca_3219_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3215_start <= Xentry_3198_symbol; -- control passed to block
              Xentry_3216_symbol  <= word_access_3_3215_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_3/$entry
              cr_3218_symbol <= Xentry_3216_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_3/cr
              ptr_deref_494_load_3_req_1 <= cr_3218_symbol; -- link to DP
              ca_3219_symbol <= ptr_deref_494_load_3_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_3/ca
              Xexit_3217_symbol <= ca_3219_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_3/$exit
              word_access_3_3215_symbol <= Xexit_3217_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_3
            Xexit_3199_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/$exit 
              signal Xexit_3199_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3199_predecessors(0) <= word_access_0_3200_symbol;
              Xexit_3199_predecessors(1) <= word_access_1_3205_symbol;
              Xexit_3199_predecessors(2) <= word_access_2_3210_symbol;
              Xexit_3199_predecessors(3) <= word_access_3_3215_symbol;
              Xexit_3199_join: join -- 
                port map( -- 
                  preds => Xexit_3199_predecessors,
                  symbol_out => Xexit_3199_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/$exit
            word_access_3197_symbol <= Xexit_3199_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access
          merge_req_3220_symbol <= word_access_3197_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/merge_req
          ptr_deref_494_gather_scatter_req_0 <= merge_req_3220_symbol; -- link to DP
          merge_ack_3221_symbol <= ptr_deref_494_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/merge_ack
          Xexit_3196_symbol <= merge_ack_3221_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/$exit
          ptr_deref_494_complete_3194_symbol <= Xexit_3196_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete
        assign_stmt_499_active_x_x3222_symbol <= type_cast_498_complete_3227_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_499_active_
        assign_stmt_499_completed_x_x3223_symbol <= assign_stmt_499_active_x_x3222_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_499_completed_
        type_cast_498_active_x_x3224_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_active_ 
          signal type_cast_498_active_x_x3224_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_498_active_x_x3224_predecessors(0) <= type_cast_498_trigger_x_x3225_symbol;
          type_cast_498_active_x_x3224_predecessors(1) <= simple_obj_ref_497_complete_3226_symbol;
          type_cast_498_active_x_x3224_join: join -- 
            port map( -- 
              preds => type_cast_498_active_x_x3224_predecessors,
              symbol_out => type_cast_498_active_x_x3224_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_active_
        type_cast_498_trigger_x_x3225_symbol <= Xentry_2845_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_trigger_
        simple_obj_ref_497_complete_3226_symbol <= assign_stmt_495_completed_x_x3162_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_497_complete
        type_cast_498_complete_3227: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete 
          signal type_cast_498_complete_3227_start: Boolean;
          signal Xentry_3228_symbol: Boolean;
          signal Xexit_3229_symbol: Boolean;
          signal req_3230_symbol : Boolean;
          signal ack_3231_symbol : Boolean;
          -- 
        begin -- 
          type_cast_498_complete_3227_start <= type_cast_498_active_x_x3224_symbol; -- control passed to block
          Xentry_3228_symbol  <= type_cast_498_complete_3227_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/$entry
          req_3230_symbol <= Xentry_3228_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/req
          type_cast_498_inst_req_0 <= req_3230_symbol; -- link to DP
          ack_3231_symbol <= type_cast_498_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/ack
          Xexit_3229_symbol <= ack_3231_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/$exit
          type_cast_498_complete_3227_symbol <= Xexit_3229_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete
        Xexit_2846_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/$exit 
          signal Xexit_2846_predecessors: BooleanArray(6 downto 0);
          -- 
        begin -- 
          Xexit_2846_predecessors(0) <= assign_stmt_474_completed_x_x2848_symbol;
          Xexit_2846_predecessors(1) <= ptr_deref_472_base_address_calculated_2852_symbol;
          Xexit_2846_predecessors(2) <= ptr_deref_477_base_address_calculated_2913_symbol;
          Xexit_2846_predecessors(3) <= ptr_deref_481_base_address_calculated_2974_symbol;
          Xexit_2846_predecessors(4) <= assign_stmt_491_completed_x_x3057_symbol;
          Xexit_2846_predecessors(5) <= ptr_deref_494_base_address_calculated_3165_symbol;
          Xexit_2846_predecessors(6) <= assign_stmt_499_completed_x_x3223_symbol;
          Xexit_2846_join: join -- 
            port map( -- 
              preds => Xexit_2846_predecessors,
              symbol_out => Xexit_2846_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/$exit
        assign_stmt_474_to_assign_stmt_504_2844_symbol <= Xexit_2846_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504
      assign_stmt_508_3232: Block -- branch_block_stmt_405/assign_stmt_508 
        signal assign_stmt_508_3232_start: Boolean;
        signal Xentry_3233_symbol: Boolean;
        signal Xexit_3234_symbol: Boolean;
        signal assign_stmt_508_active_x_x3235_symbol : Boolean;
        signal assign_stmt_508_completed_x_x3236_symbol : Boolean;
        signal type_cast_507_active_x_x3237_symbol : Boolean;
        signal type_cast_507_trigger_x_x3238_symbol : Boolean;
        signal simple_obj_ref_506_complete_3239_symbol : Boolean;
        signal type_cast_507_complete_3240_symbol : Boolean;
        signal simple_obj_ref_505_trigger_x_x3245_symbol : Boolean;
        signal simple_obj_ref_505_complete_3246_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_508_3232_start <= assign_stmt_508_x_xentry_x_xx_x2606_symbol; -- control passed to block
        Xentry_3233_symbol  <= assign_stmt_508_3232_start; -- transition branch_block_stmt_405/assign_stmt_508/$entry
        assign_stmt_508_active_x_x3235_symbol <= type_cast_507_complete_3240_symbol; -- transition branch_block_stmt_405/assign_stmt_508/assign_stmt_508_active_
        assign_stmt_508_completed_x_x3236_symbol <= simple_obj_ref_505_complete_3246_symbol; -- transition branch_block_stmt_405/assign_stmt_508/assign_stmt_508_completed_
        type_cast_507_active_x_x3237_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_508/type_cast_507_active_ 
          signal type_cast_507_active_x_x3237_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_507_active_x_x3237_predecessors(0) <= type_cast_507_trigger_x_x3238_symbol;
          type_cast_507_active_x_x3237_predecessors(1) <= simple_obj_ref_506_complete_3239_symbol;
          type_cast_507_active_x_x3237_join: join -- 
            port map( -- 
              preds => type_cast_507_active_x_x3237_predecessors,
              symbol_out => type_cast_507_active_x_x3237_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_508/type_cast_507_active_
        type_cast_507_trigger_x_x3238_symbol <= Xentry_3233_symbol; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_trigger_
        simple_obj_ref_506_complete_3239_symbol <= Xentry_3233_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_506_complete
        type_cast_507_complete_3240: Block -- branch_block_stmt_405/assign_stmt_508/type_cast_507_complete 
          signal type_cast_507_complete_3240_start: Boolean;
          signal Xentry_3241_symbol: Boolean;
          signal Xexit_3242_symbol: Boolean;
          signal req_3243_symbol : Boolean;
          signal ack_3244_symbol : Boolean;
          -- 
        begin -- 
          type_cast_507_complete_3240_start <= type_cast_507_active_x_x3237_symbol; -- control passed to block
          Xentry_3241_symbol  <= type_cast_507_complete_3240_start; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/$entry
          req_3243_symbol <= Xentry_3241_symbol; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/req
          type_cast_507_inst_req_0 <= req_3243_symbol; -- link to DP
          ack_3244_symbol <= type_cast_507_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/ack
          Xexit_3242_symbol <= ack_3244_symbol; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/$exit
          type_cast_507_complete_3240_symbol <= Xexit_3242_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_508/type_cast_507_complete
        simple_obj_ref_505_trigger_x_x3245_symbol <= assign_stmt_508_active_x_x3235_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_trigger_
        simple_obj_ref_505_complete_3246: Block -- branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete 
          signal simple_obj_ref_505_complete_3246_start: Boolean;
          signal Xentry_3247_symbol: Boolean;
          signal Xexit_3248_symbol: Boolean;
          signal pipe_wreq_3249_symbol : Boolean;
          signal pipe_wack_3250_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_505_complete_3246_start <= simple_obj_ref_505_trigger_x_x3245_symbol; -- control passed to block
          Xentry_3247_symbol  <= simple_obj_ref_505_complete_3246_start; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/$entry
          pipe_wreq_3249_symbol <= Xentry_3247_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/pipe_wreq
          simple_obj_ref_505_inst_req_0 <= pipe_wreq_3249_symbol; -- link to DP
          pipe_wack_3250_symbol <= simple_obj_ref_505_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/pipe_wack
          Xexit_3248_symbol <= pipe_wack_3250_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/$exit
          simple_obj_ref_505_complete_3246_symbol <= Xexit_3248_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete
        Xexit_3234_symbol <= assign_stmt_508_completed_x_x3236_symbol; -- transition branch_block_stmt_405/assign_stmt_508/$exit
        assign_stmt_508_3232_symbol <= Xexit_3234_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_508
      bb_0_bb_1_PhiReq_3251: Block -- branch_block_stmt_405/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_3251_start: Boolean;
        signal Xentry_3252_symbol: Boolean;
        signal Xexit_3253_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_3251_start <= bb_0_bb_1_2584_symbol; -- control passed to block
        Xentry_3252_symbol  <= bb_0_bb_1_PhiReq_3251_start; -- transition branch_block_stmt_405/bb_0_bb_1_PhiReq/$entry
        Xexit_3253_symbol <= Xentry_3252_symbol; -- transition branch_block_stmt_405/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_3251_symbol <= Xexit_3253_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_0_bb_1_PhiReq
      bb_1_bb_1_PhiReq_3254: Block -- branch_block_stmt_405/bb_1_bb_1_PhiReq 
        signal bb_1_bb_1_PhiReq_3254_start: Boolean;
        signal Xentry_3255_symbol: Boolean;
        signal Xexit_3256_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_1_PhiReq_3254_start <= bb_1_bb_1_2822_symbol; -- control passed to block
        Xentry_3255_symbol  <= bb_1_bb_1_PhiReq_3254_start; -- transition branch_block_stmt_405/bb_1_bb_1_PhiReq/$entry
        Xexit_3256_symbol <= Xentry_3255_symbol; -- transition branch_block_stmt_405/bb_1_bb_1_PhiReq/$exit
        bb_1_bb_1_PhiReq_3254_symbol <= Xexit_3256_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_1_bb_1_PhiReq
      bb_2_bb_1_PhiReq_3257: Block -- branch_block_stmt_405/bb_2_bb_1_PhiReq 
        signal bb_2_bb_1_PhiReq_3257_start: Boolean;
        signal Xentry_3258_symbol: Boolean;
        signal Xexit_3259_symbol: Boolean;
        -- 
      begin -- 
        bb_2_bb_1_PhiReq_3257_start <= bb_2_bb_1_2608_symbol; -- control passed to block
        Xentry_3258_symbol  <= bb_2_bb_1_PhiReq_3257_start; -- transition branch_block_stmt_405/bb_2_bb_1_PhiReq/$entry
        Xexit_3259_symbol <= Xentry_3258_symbol; -- transition branch_block_stmt_405/bb_2_bb_1_PhiReq/$exit
        bb_2_bb_1_PhiReq_3257_symbol <= Xexit_3259_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_2_bb_1_PhiReq
      merge_stmt_417_PhiReqMerge_3260_symbol  <=  bb_0_bb_1_PhiReq_3251_symbol or bb_1_bb_1_PhiReq_3254_symbol or bb_2_bb_1_PhiReq_3257_symbol; -- place branch_block_stmt_405/merge_stmt_417_PhiReqMerge (optimized away) 
      merge_stmt_417_PhiAck_3261: Block -- branch_block_stmt_405/merge_stmt_417_PhiAck 
        signal merge_stmt_417_PhiAck_3261_start: Boolean;
        signal Xentry_3262_symbol: Boolean;
        signal Xexit_3263_symbol: Boolean;
        signal dummy_3264_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_417_PhiAck_3261_start <= merge_stmt_417_PhiReqMerge_3260_symbol; -- control passed to block
        Xentry_3262_symbol  <= merge_stmt_417_PhiAck_3261_start; -- transition branch_block_stmt_405/merge_stmt_417_PhiAck/$entry
        dummy_3264_symbol <= Xentry_3262_symbol; -- transition branch_block_stmt_405/merge_stmt_417_PhiAck/dummy
        Xexit_3263_symbol <= dummy_3264_symbol; -- transition branch_block_stmt_405/merge_stmt_417_PhiAck/$exit
        merge_stmt_417_PhiAck_3261_symbol <= Xexit_3263_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/merge_stmt_417_PhiAck
      merge_stmt_461_dead_link_3265: Block -- branch_block_stmt_405/merge_stmt_461_dead_link 
        signal merge_stmt_461_dead_link_3265_start: Boolean;
        signal Xentry_3266_symbol: Boolean;
        signal Xexit_3267_symbol: Boolean;
        signal dead_transition_3268_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_461_dead_link_3265_start <= merge_stmt_461_x_xentry_x_xx_x2598_symbol; -- control passed to block
        Xentry_3266_symbol  <= merge_stmt_461_dead_link_3265_start; -- transition branch_block_stmt_405/merge_stmt_461_dead_link/$entry
        dead_transition_3268_symbol <= false;
        Xexit_3267_symbol <= dead_transition_3268_symbol; -- transition branch_block_stmt_405/merge_stmt_461_dead_link/$exit
        merge_stmt_461_dead_link_3265_symbol <= Xexit_3267_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/merge_stmt_461_dead_link
      bb_1_bb_2_PhiReq_3269: Block -- branch_block_stmt_405/bb_1_bb_2_PhiReq 
        signal bb_1_bb_2_PhiReq_3269_start: Boolean;
        signal Xentry_3270_symbol: Boolean;
        signal Xexit_3271_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_2_PhiReq_3269_start <= bb_1_bb_2_2821_symbol; -- control passed to block
        Xentry_3270_symbol  <= bb_1_bb_2_PhiReq_3269_start; -- transition branch_block_stmt_405/bb_1_bb_2_PhiReq/$entry
        Xexit_3271_symbol <= Xentry_3270_symbol; -- transition branch_block_stmt_405/bb_1_bb_2_PhiReq/$exit
        bb_1_bb_2_PhiReq_3269_symbol <= Xexit_3271_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_1_bb_2_PhiReq
      merge_stmt_461_PhiReqMerge_3272_symbol  <=  bb_1_bb_2_PhiReq_3269_symbol; -- place branch_block_stmt_405/merge_stmt_461_PhiReqMerge (optimized away) 
      merge_stmt_461_PhiAck_3273: Block -- branch_block_stmt_405/merge_stmt_461_PhiAck 
        signal merge_stmt_461_PhiAck_3273_start: Boolean;
        signal Xentry_3274_symbol: Boolean;
        signal Xexit_3275_symbol: Boolean;
        signal dummy_3276_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_461_PhiAck_3273_start <= merge_stmt_461_PhiReqMerge_3272_symbol; -- control passed to block
        Xentry_3274_symbol  <= merge_stmt_461_PhiAck_3273_start; -- transition branch_block_stmt_405/merge_stmt_461_PhiAck/$entry
        dummy_3276_symbol <= Xentry_3274_symbol; -- transition branch_block_stmt_405/merge_stmt_461_PhiAck/dummy
        Xexit_3275_symbol <= dummy_3276_symbol; -- transition branch_block_stmt_405/merge_stmt_461_PhiAck/$exit
        merge_stmt_461_PhiAck_3273_symbol <= Xexit_3275_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/merge_stmt_461_PhiAck
      Xexit_2579_symbol <= branch_block_stmt_405_x_xexit_x_xx_x2581_symbol; -- transition branch_block_stmt_405/$exit
      branch_block_stmt_405_2577_symbol <= Xexit_2579_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_405
    Xexit_2576_symbol <= branch_block_stmt_405_2577_symbol; -- transition $exit
    fin  <=  '1' when Xexit_2576_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_486_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_486_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_486_root_address : std_logic_vector(5 downto 0);
    signal iNsTr_10_466 : std_logic_vector(31 downto 0);
    signal iNsTr_11_470 : std_logic_vector(31 downto 0);
    signal iNsTr_13_478 : std_logic_vector(31 downto 0);
    signal iNsTr_14_482 : std_logic_vector(31 downto 0);
    signal iNsTr_15_487 : std_logic_vector(31 downto 0);
    signal iNsTr_17_495 : std_logic_vector(31 downto 0);
    signal iNsTr_18_499 : std_logic_vector(31 downto 0);
    signal iNsTr_19_504 : std_logic_vector(31 downto 0);
    signal iNsTr_1_422 : std_logic_vector(31 downto 0);
    signal iNsTr_3_431 : std_logic_vector(31 downto 0);
    signal iNsTr_4_435 : std_logic_vector(31 downto 0);
    signal iNsTr_5_439 : std_logic_vector(31 downto 0);
    signal iNsTr_7_447 : std_logic_vector(31 downto 0);
    signal iNsTr_8_454 : std_logic_vector(0 downto 0);
    signal lptr_411 : std_logic_vector(31 downto 0);
    signal nval_415 : std_logic_vector(31 downto 0);
    signal ptr_deref_441_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_441_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_441_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_441_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_441_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_441_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_441_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_441_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_441_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_446_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_446_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_446_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_446_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_446_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_446_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_446_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_446_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_472_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_472_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_472_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_472_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_472_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_472_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_472_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_472_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_472_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_477_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_477_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_477_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_477_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_477_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_477_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_477_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_477_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_481_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_481_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_481_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_481_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_481_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_481_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_481_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_481_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_489_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_489_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_489_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_489_word_offset_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_494_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_494_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_494_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_494_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_494_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_494_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_494_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_494_word_address_3 : std_logic_vector(5 downto 0);
    signal simple_obj_ref_433_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_468_wire : std_logic_vector(31 downto 0);
    signal type_cast_425_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_450_wire : std_logic_vector(31 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_507_wire : std_logic_vector(31 downto 0);
    signal xxinput_modulexxbodyxxlptr_alloc_base_address : std_logic_vector(5 downto 0);
    signal xxinput_modulexxbodyxxnval_alloc_base_address : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    array_obj_ref_486_final_offset <= "000100";
    iNsTr_10_466 <= "00000000000000000000000000000000";
    iNsTr_19_504 <= "00000000000000000000000000000000";
    iNsTr_1_422 <= "00000000000000000000000000000000";
    iNsTr_3_431 <= "00000000000000000000000000000000";
    lptr_411 <= "00000000000000000000000000101001";
    nval_415 <= "00000000000000000000000000101101";
    ptr_deref_441_word_address_0 <= "101001";
    ptr_deref_441_word_address_1 <= "101010";
    ptr_deref_441_word_address_2 <= "101011";
    ptr_deref_441_word_address_3 <= "101100";
    ptr_deref_446_word_address_0 <= "101001";
    ptr_deref_446_word_address_1 <= "101010";
    ptr_deref_446_word_address_2 <= "101011";
    ptr_deref_446_word_address_3 <= "101100";
    ptr_deref_472_word_address_0 <= "101101";
    ptr_deref_472_word_address_1 <= "101110";
    ptr_deref_472_word_address_2 <= "101111";
    ptr_deref_472_word_address_3 <= "110000";
    ptr_deref_477_word_address_0 <= "101101";
    ptr_deref_477_word_address_1 <= "101110";
    ptr_deref_477_word_address_2 <= "101111";
    ptr_deref_477_word_address_3 <= "110000";
    ptr_deref_481_word_address_0 <= "101001";
    ptr_deref_481_word_address_1 <= "101010";
    ptr_deref_481_word_address_2 <= "101011";
    ptr_deref_481_word_address_3 <= "101100";
    ptr_deref_489_word_offset_0 <= "000000";
    ptr_deref_489_word_offset_1 <= "000001";
    ptr_deref_489_word_offset_2 <= "000010";
    ptr_deref_489_word_offset_3 <= "000011";
    ptr_deref_494_word_address_0 <= "101001";
    ptr_deref_494_word_address_1 <= "101010";
    ptr_deref_494_word_address_2 <= "101011";
    ptr_deref_494_word_address_3 <= "101100";
    type_cast_425_wire_constant <= "00000010";
    type_cast_452_wire_constant <= "00000000000000000000000000000000";
    xxinput_modulexxbodyxxlptr_alloc_base_address <= "101001";
    xxinput_modulexxbodyxxnval_alloc_base_address <= "101101";
    array_obj_ref_486_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_14_482, dout => array_obj_ref_486_resized_base_address, req => array_obj_ref_486_base_resize_req_0, ack => array_obj_ref_486_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_486_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_486_root_address, dout => iNsTr_15_487, req => array_obj_ref_486_final_reg_req_0, ack => array_obj_ref_486_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_489_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_15_487, dout => ptr_deref_489_resized_base_address, req => ptr_deref_489_base_resize_req_0, ack => ptr_deref_489_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_434_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_433_wire, dout => iNsTr_4_435, req => type_cast_434_inst_req_0, ack => type_cast_434_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_438_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_4_435, dout => iNsTr_5_439, req => type_cast_438_inst_req_0, ack => type_cast_438_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_469_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_468_wire, dout => iNsTr_11_470, req => type_cast_469_inst_req_0, ack => type_cast_469_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_498_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_17_495, dout => iNsTr_18_499, req => type_cast_498_inst_req_0, ack => type_cast_498_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_507_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_18_499, dout => type_cast_507_wire, req => type_cast_507_inst_req_0, ack => type_cast_507_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_441_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_441_gather_scatter_ack_0 <= ptr_deref_441_gather_scatter_req_0;
      aggregated_sig <= iNsTr_5_439;
      ptr_deref_441_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_441_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_441_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_441_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_446_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_446_gather_scatter_ack_0 <= ptr_deref_446_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_446_data_0 & ptr_deref_446_data_1 & ptr_deref_446_data_2 & ptr_deref_446_data_3;
      iNsTr_7_447 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_472_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_472_gather_scatter_ack_0 <= ptr_deref_472_gather_scatter_req_0;
      aggregated_sig <= iNsTr_11_470;
      ptr_deref_472_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_472_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_472_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_472_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_477_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_477_gather_scatter_ack_0 <= ptr_deref_477_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_477_data_0 & ptr_deref_477_data_1 & ptr_deref_477_data_2 & ptr_deref_477_data_3;
      iNsTr_13_478 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_481_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_481_gather_scatter_ack_0 <= ptr_deref_481_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_481_data_0 & ptr_deref_481_data_1 & ptr_deref_481_data_2 & ptr_deref_481_data_3;
      iNsTr_14_482 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_489_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_489_gather_scatter_ack_0 <= ptr_deref_489_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_478;
      ptr_deref_489_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_489_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_489_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_489_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_489_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_489_root_address_inst_ack_0 <= ptr_deref_489_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_489_resized_base_address;
      ptr_deref_489_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_494_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_494_gather_scatter_ack_0 <= ptr_deref_494_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_494_data_0 & ptr_deref_494_data_1 & ptr_deref_494_data_2 & ptr_deref_494_data_3;
      iNsTr_17_495 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_455_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_8_454;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_455_branch_req_0,
          ack0 => if_stmt_455_branch_ack_0,
          ack1 => if_stmt_455_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_486_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_486_resized_base_address;
      array_obj_ref_486_root_address <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000100",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_486_root_address_inst_req_0,
          ackL => array_obj_ref_486_root_address_inst_ack_0,
          reqR => array_obj_ref_486_root_address_inst_req_1,
          ackR => array_obj_ref_486_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_453_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_450_wire;
      iNsTr_8_454 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_453_inst_req_0,
          ackL => binary_453_inst_ack_0,
          reqR => binary_453_inst_req_1,
          ackR => binary_453_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ptr_deref_489_addr_0 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_0 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_489_addr_0_req_0,
          ackL => ptr_deref_489_addr_0_ack_0,
          reqR => ptr_deref_489_addr_0_req_1,
          ackR => ptr_deref_489_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ptr_deref_489_addr_1 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_1 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_489_addr_1_req_0,
          ackL => ptr_deref_489_addr_1_ack_0,
          reqR => ptr_deref_489_addr_1_req_1,
          ackR => ptr_deref_489_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ptr_deref_489_addr_2 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_2 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_489_addr_2_req_0,
          ackL => ptr_deref_489_addr_2_ack_0,
          reqR => ptr_deref_489_addr_2_req_1,
          ackR => ptr_deref_489_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : ptr_deref_489_addr_3 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_3 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000011",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_489_addr_3_req_0,
          ackL => ptr_deref_489_addr_3_ack_0,
          reqR => ptr_deref_489_addr_3_req_1,
          ackR => ptr_deref_489_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : type_cast_450_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_7_447;
      type_cast_450_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => type_cast_450_inst_req_0,
          ackL => type_cast_450_inst_ack_0,
          reqR => type_cast_450_inst_req_1,
          ackR => type_cast_450_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared load operator group (0) : ptr_deref_446_load_0 ptr_deref_477_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_446_load_0_req_0;
      reqL(0) <= ptr_deref_477_load_0_req_0;
      ptr_deref_446_load_0_ack_0 <= ackL(1);
      ptr_deref_477_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_446_load_0_req_1;
      reqR(0) <= ptr_deref_477_load_0_req_1;
      ptr_deref_446_load_0_ack_1 <= ackR(1);
      ptr_deref_477_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_446_word_address_0 & ptr_deref_477_word_address_0;
      ptr_deref_446_data_0 <= data_out(15 downto 8);
      ptr_deref_477_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(11),
          mack => memory_space_1_lr_ack(11),
          maddr => memory_space_1_lr_addr(71 downto 66),
          mtag => memory_space_1_lr_tag(35 downto 33),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(11),
          mack => memory_space_1_lc_ack(11),
          mdata => memory_space_1_lc_data(95 downto 88),
          mtag => memory_space_1_lc_tag(35 downto 33),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_477_load_1 ptr_deref_446_load_1 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_477_load_1_req_0;
      reqL(0) <= ptr_deref_446_load_1_req_0;
      ptr_deref_477_load_1_ack_0 <= ackL(1);
      ptr_deref_446_load_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_477_load_1_req_1;
      reqR(0) <= ptr_deref_446_load_1_req_1;
      ptr_deref_477_load_1_ack_1 <= ackR(1);
      ptr_deref_446_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_477_word_address_1 & ptr_deref_446_word_address_1;
      ptr_deref_477_data_1 <= data_out(15 downto 8);
      ptr_deref_446_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(10),
          mack => memory_space_1_lr_ack(10),
          maddr => memory_space_1_lr_addr(65 downto 60),
          mtag => memory_space_1_lr_tag(32 downto 30),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(10),
          mack => memory_space_1_lc_ack(10),
          mdata => memory_space_1_lc_data(87 downto 80),
          mtag => memory_space_1_lc_tag(32 downto 30),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_477_load_2 ptr_deref_446_load_2 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_477_load_2_req_0;
      reqL(0) <= ptr_deref_446_load_2_req_0;
      ptr_deref_477_load_2_ack_0 <= ackL(1);
      ptr_deref_446_load_2_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_477_load_2_req_1;
      reqR(0) <= ptr_deref_446_load_2_req_1;
      ptr_deref_477_load_2_ack_1 <= ackR(1);
      ptr_deref_446_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_477_word_address_2 & ptr_deref_446_word_address_2;
      ptr_deref_477_data_2 <= data_out(15 downto 8);
      ptr_deref_446_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(9),
          mack => memory_space_1_lr_ack(9),
          maddr => memory_space_1_lr_addr(59 downto 54),
          mtag => memory_space_1_lr_tag(29 downto 27),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(9),
          mack => memory_space_1_lc_ack(9),
          mdata => memory_space_1_lc_data(79 downto 72),
          mtag => memory_space_1_lc_tag(29 downto 27),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_446_load_3 ptr_deref_477_load_3 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_446_load_3_req_0;
      reqL(0) <= ptr_deref_477_load_3_req_0;
      ptr_deref_446_load_3_ack_0 <= ackL(1);
      ptr_deref_477_load_3_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_446_load_3_req_1;
      reqR(0) <= ptr_deref_477_load_3_req_1;
      ptr_deref_446_load_3_ack_1 <= ackR(1);
      ptr_deref_477_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_446_word_address_3 & ptr_deref_477_word_address_3;
      ptr_deref_446_data_3 <= data_out(15 downto 8);
      ptr_deref_477_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(8),
          mack => memory_space_1_lr_ack(8),
          maddr => memory_space_1_lr_addr(53 downto 48),
          mtag => memory_space_1_lr_tag(26 downto 24),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(8),
          mack => memory_space_1_lc_ack(8),
          mdata => memory_space_1_lc_data(71 downto 64),
          mtag => memory_space_1_lc_tag(26 downto 24),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_481_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_481_load_0_req_0;
      ptr_deref_481_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_481_load_0_req_1;
      ptr_deref_481_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_481_word_address_0;
      ptr_deref_481_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(7),
          mack => memory_space_1_lr_ack(7),
          maddr => memory_space_1_lr_addr(47 downto 42),
          mtag => memory_space_1_lr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(7),
          mack => memory_space_1_lc_ack(7),
          mdata => memory_space_1_lc_data(63 downto 56),
          mtag => memory_space_1_lc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_481_load_1 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_481_load_1_req_0;
      ptr_deref_481_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_481_load_1_req_1;
      ptr_deref_481_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_481_word_address_1;
      ptr_deref_481_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(6),
          mack => memory_space_1_lr_ack(6),
          maddr => memory_space_1_lr_addr(41 downto 36),
          mtag => memory_space_1_lr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(6),
          mack => memory_space_1_lc_ack(6),
          mdata => memory_space_1_lc_data(55 downto 48),
          mtag => memory_space_1_lc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_481_load_2 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_481_load_2_req_0;
      ptr_deref_481_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_481_load_2_req_1;
      ptr_deref_481_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_481_word_address_2;
      ptr_deref_481_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(5),
          mack => memory_space_1_lr_ack(5),
          maddr => memory_space_1_lr_addr(35 downto 30),
          mtag => memory_space_1_lr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(5),
          mack => memory_space_1_lc_ack(5),
          mdata => memory_space_1_lc_data(47 downto 40),
          mtag => memory_space_1_lc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_481_load_3 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_481_load_3_req_0;
      ptr_deref_481_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_481_load_3_req_1;
      ptr_deref_481_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_481_word_address_3;
      ptr_deref_481_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(4),
          mack => memory_space_1_lr_ack(4),
          maddr => memory_space_1_lr_addr(29 downto 24),
          mtag => memory_space_1_lr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(4),
          mack => memory_space_1_lc_ack(4),
          mdata => memory_space_1_lc_data(39 downto 32),
          mtag => memory_space_1_lc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared load operator group (8) : ptr_deref_494_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_494_load_0_req_0;
      ptr_deref_494_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_494_load_0_req_1;
      ptr_deref_494_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_494_word_address_0;
      ptr_deref_494_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(3),
          mack => memory_space_1_lr_ack(3),
          maddr => memory_space_1_lr_addr(23 downto 18),
          mtag => memory_space_1_lr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(3),
          mack => memory_space_1_lc_ack(3),
          mdata => memory_space_1_lc_data(31 downto 24),
          mtag => memory_space_1_lc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- shared load operator group (9) : ptr_deref_494_load_1 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_494_load_1_req_0;
      ptr_deref_494_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_494_load_1_req_1;
      ptr_deref_494_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_494_word_address_1;
      ptr_deref_494_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(2),
          mack => memory_space_1_lr_ack(2),
          maddr => memory_space_1_lr_addr(17 downto 12),
          mtag => memory_space_1_lr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(2),
          mack => memory_space_1_lc_ack(2),
          mdata => memory_space_1_lc_data(23 downto 16),
          mtag => memory_space_1_lc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    -- shared load operator group (10) : ptr_deref_494_load_2 
    LoadGroup10: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_494_load_2_req_0;
      ptr_deref_494_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_494_load_2_req_1;
      ptr_deref_494_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_494_word_address_2;
      ptr_deref_494_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(1),
          mack => memory_space_1_lr_ack(1),
          maddr => memory_space_1_lr_addr(11 downto 6),
          mtag => memory_space_1_lr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(1),
          mack => memory_space_1_lc_ack(1),
          mdata => memory_space_1_lc_data(15 downto 8),
          mtag => memory_space_1_lc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 10
    -- shared load operator group (11) : ptr_deref_494_load_3 
    LoadGroup11: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_494_load_3_req_0;
      ptr_deref_494_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_494_load_3_req_1;
      ptr_deref_494_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_494_word_address_3;
      ptr_deref_494_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(5 downto 0),
          mtag => memory_space_1_lr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 11
    -- shared store operator group (0) : ptr_deref_441_store_0 ptr_deref_472_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_441_store_0_req_0;
      reqL(0) <= ptr_deref_472_store_0_req_0;
      ptr_deref_441_store_0_ack_0 <= ackL(1);
      ptr_deref_472_store_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_441_store_0_req_1;
      reqR(0) <= ptr_deref_472_store_0_req_1;
      ptr_deref_441_store_0_ack_1 <= ackR(1);
      ptr_deref_472_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_441_word_address_0 & ptr_deref_472_word_address_0;
      data_in <= ptr_deref_441_data_0 & ptr_deref_472_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(7),
          mack => memory_space_1_sr_ack(7),
          maddr => memory_space_1_sr_addr(47 downto 42),
          mdata => memory_space_1_sr_data(63 downto 56),
          mtag => memory_space_1_sr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(7),
          mack => memory_space_1_sc_ack(7),
          mtag => memory_space_1_sc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_472_store_1 ptr_deref_441_store_1 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_472_store_1_req_0;
      reqL(0) <= ptr_deref_441_store_1_req_0;
      ptr_deref_472_store_1_ack_0 <= ackL(1);
      ptr_deref_441_store_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_472_store_1_req_1;
      reqR(0) <= ptr_deref_441_store_1_req_1;
      ptr_deref_472_store_1_ack_1 <= ackR(1);
      ptr_deref_441_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_472_word_address_1 & ptr_deref_441_word_address_1;
      data_in <= ptr_deref_472_data_1 & ptr_deref_441_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(6),
          mack => memory_space_1_sr_ack(6),
          maddr => memory_space_1_sr_addr(41 downto 36),
          mdata => memory_space_1_sr_data(55 downto 48),
          mtag => memory_space_1_sr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(6),
          mack => memory_space_1_sc_ack(6),
          mtag => memory_space_1_sc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_441_store_2 ptr_deref_472_store_2 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_441_store_2_req_0;
      reqL(0) <= ptr_deref_472_store_2_req_0;
      ptr_deref_441_store_2_ack_0 <= ackL(1);
      ptr_deref_472_store_2_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_441_store_2_req_1;
      reqR(0) <= ptr_deref_472_store_2_req_1;
      ptr_deref_441_store_2_ack_1 <= ackR(1);
      ptr_deref_472_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_441_word_address_2 & ptr_deref_472_word_address_2;
      data_in <= ptr_deref_441_data_2 & ptr_deref_472_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(5),
          mack => memory_space_1_sr_ack(5),
          maddr => memory_space_1_sr_addr(35 downto 30),
          mdata => memory_space_1_sr_data(47 downto 40),
          mtag => memory_space_1_sr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(5),
          mack => memory_space_1_sc_ack(5),
          mtag => memory_space_1_sc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_472_store_3 ptr_deref_441_store_3 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_472_store_3_req_0;
      reqL(0) <= ptr_deref_441_store_3_req_0;
      ptr_deref_472_store_3_ack_0 <= ackL(1);
      ptr_deref_441_store_3_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_472_store_3_req_1;
      reqR(0) <= ptr_deref_441_store_3_req_1;
      ptr_deref_472_store_3_ack_1 <= ackR(1);
      ptr_deref_441_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_472_word_address_3 & ptr_deref_441_word_address_3;
      data_in <= ptr_deref_472_data_3 & ptr_deref_441_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(4),
          mack => memory_space_1_sr_ack(4),
          maddr => memory_space_1_sr_addr(29 downto 24),
          mdata => memory_space_1_sr_data(39 downto 32),
          mtag => memory_space_1_sr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(4),
          mack => memory_space_1_sc_ack(4),
          mtag => memory_space_1_sc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_489_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_489_store_0_req_0;
      ptr_deref_489_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_489_store_0_req_1;
      ptr_deref_489_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_489_word_address_0;
      data_in <= ptr_deref_489_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(3),
          mack => memory_space_1_sr_ack(3),
          maddr => memory_space_1_sr_addr(23 downto 18),
          mdata => memory_space_1_sr_data(31 downto 24),
          mtag => memory_space_1_sr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(3),
          mack => memory_space_1_sc_ack(3),
          mtag => memory_space_1_sc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_489_store_1 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_489_store_1_req_0;
      ptr_deref_489_store_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_489_store_1_req_1;
      ptr_deref_489_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_489_word_address_1;
      data_in <= ptr_deref_489_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(2),
          mack => memory_space_1_sr_ack(2),
          maddr => memory_space_1_sr_addr(17 downto 12),
          mdata => memory_space_1_sr_data(23 downto 16),
          mtag => memory_space_1_sr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(2),
          mack => memory_space_1_sc_ack(2),
          mtag => memory_space_1_sc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_489_store_2 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_489_store_2_req_0;
      ptr_deref_489_store_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_489_store_2_req_1;
      ptr_deref_489_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_489_word_address_2;
      data_in <= ptr_deref_489_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(1),
          mack => memory_space_1_sr_ack(1),
          maddr => memory_space_1_sr_addr(11 downto 6),
          mdata => memory_space_1_sr_data(15 downto 8),
          mtag => memory_space_1_sr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(1),
          mack => memory_space_1_sc_ack(1),
          mtag => memory_space_1_sc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_489_store_3 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_489_store_3_req_0;
      ptr_deref_489_store_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_489_store_3_req_1;
      ptr_deref_489_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_489_word_address_3;
      data_in <= ptr_deref_489_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(5 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : simple_obj_ref_433_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_433_inst_req_0;
      simple_obj_ref_433_inst_ack_0 <= ack(0);
      simple_obj_ref_433_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_get_pipe_read_req(0),
          oack => free_queue_get_pipe_read_ack(0),
          odata => free_queue_get_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_468_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_468_inst_req_0;
      simple_obj_ref_468_inst_ack_0 <= ack(0);
      simple_obj_ref_468_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => input_data_pipe_read_req(0),
          oack => input_data_pipe_read_ack(0),
          odata => input_data_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_423_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_423_inst_req_0;
      simple_obj_ref_423_inst_ack_0 <= ack(0);
      data_in <= type_cast_425_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_505_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_505_inst_req_0;
      simple_obj_ref_505_inst_ack_0 <= ack(0);
      data_in <= type_cast_507_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => foo_in_pipe_write_req(0),
          oack => foo_in_pipe_write_ack(0),
          odata => foo_in_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity mem_load_x_x is -- 
  port ( -- 
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(7 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity mem_load_x_x;
architecture Default of mem_load_x_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal binary_10_inst_ack_0 : boolean;
  signal binary_10_inst_ack_1 : boolean;
  signal binary_12_inst_ack_1 : boolean;
  signal array_obj_ref_13_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_13_offset_inst_ack_0 : boolean;
  signal binary_12_inst_req_1 : boolean;
  signal array_obj_ref_13_index_0_rename_req_0 : boolean;
  signal binary_10_inst_req_0 : boolean;
  signal array_obj_ref_13_index_0_resize_req_0 : boolean;
  signal binary_12_inst_ack_0 : boolean;
  signal array_obj_ref_13_root_address_inst_req_0 : boolean;
  signal array_obj_ref_13_addr_0_ack_0 : boolean;
  signal array_obj_ref_13_gather_scatter_ack_0 : boolean;
  signal binary_10_inst_req_1 : boolean;
  signal array_obj_ref_13_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_13_load_0_req_1 : boolean;
  signal array_obj_ref_13_index_0_rename_ack_0 : boolean;
  signal binary_12_inst_req_0 : boolean;
  signal array_obj_ref_13_load_0_ack_1 : boolean;
  signal array_obj_ref_13_gather_scatter_req_0 : boolean;
  signal array_obj_ref_13_addr_0_req_0 : boolean;
  signal array_obj_ref_13_load_0_req_0 : boolean;
  signal array_obj_ref_13_offset_inst_req_0 : boolean;
  signal array_obj_ref_13_load_0_ack_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  mem_load_x_xx_xCP_3277: Block -- control-path 
    signal mem_load_x_xx_xCP_3277_start: Boolean;
    signal Xentry_3278_symbol: Boolean;
    signal Xexit_3279_symbol: Boolean;
    signal assign_stmt_14_3280_symbol : Boolean;
    -- 
  begin -- 
    mem_load_x_xx_xCP_3277_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_3278_symbol  <= mem_load_x_xx_xCP_3277_start; -- transition $entry
    assign_stmt_14_3280: Block -- assign_stmt_14 
      signal assign_stmt_14_3280_start: Boolean;
      signal Xentry_3281_symbol: Boolean;
      signal Xexit_3282_symbol: Boolean;
      signal assign_stmt_14_active_x_x3283_symbol : Boolean;
      signal assign_stmt_14_completed_x_x3284_symbol : Boolean;
      signal array_obj_ref_13_trigger_x_x3285_symbol : Boolean;
      signal array_obj_ref_13_active_x_x3286_symbol : Boolean;
      signal array_obj_ref_13_root_address_calculated_3287_symbol : Boolean;
      signal array_obj_ref_13_word_address_calculated_3288_symbol : Boolean;
      signal array_obj_ref_13_indices_scaled_3289_symbol : Boolean;
      signal array_obj_ref_13_offset_calculated_3290_symbol : Boolean;
      signal array_obj_ref_13_index_computed_0_3291_symbol : Boolean;
      signal array_obj_ref_13_index_resized_0_3292_symbol : Boolean;
      signal binary_12_active_x_x3293_symbol : Boolean;
      signal binary_12_trigger_x_x3294_symbol : Boolean;
      signal binary_10_active_x_x3295_symbol : Boolean;
      signal binary_10_trigger_x_x3296_symbol : Boolean;
      signal simple_obj_ref_8_complete_3297_symbol : Boolean;
      signal binary_10_complete_3298_symbol : Boolean;
      signal binary_12_complete_3305_symbol : Boolean;
      signal array_obj_ref_13_index_resize_0_3312_symbol : Boolean;
      signal array_obj_ref_13_index_scale_0_3317_symbol : Boolean;
      signal array_obj_ref_13_add_indices_3322_symbol : Boolean;
      signal array_obj_ref_13_base_plus_offset_3327_symbol : Boolean;
      signal array_obj_ref_13_word_addrgen_3332_symbol : Boolean;
      signal array_obj_ref_13_request_3337_symbol : Boolean;
      signal array_obj_ref_13_complete_3348_symbol : Boolean;
      -- 
    begin -- 
      assign_stmt_14_3280_start <= Xentry_3278_symbol; -- control passed to block
      Xentry_3281_symbol  <= assign_stmt_14_3280_start; -- transition assign_stmt_14/$entry
      assign_stmt_14_active_x_x3283_symbol <= array_obj_ref_13_complete_3348_symbol; -- transition assign_stmt_14/assign_stmt_14_active_
      assign_stmt_14_completed_x_x3284_symbol <= assign_stmt_14_active_x_x3283_symbol; -- transition assign_stmt_14/assign_stmt_14_completed_
      array_obj_ref_13_trigger_x_x3285_symbol <= array_obj_ref_13_word_address_calculated_3288_symbol; -- transition assign_stmt_14/array_obj_ref_13_trigger_
      array_obj_ref_13_active_x_x3286_symbol <= array_obj_ref_13_request_3337_symbol; -- transition assign_stmt_14/array_obj_ref_13_active_
      array_obj_ref_13_root_address_calculated_3287_symbol <= array_obj_ref_13_base_plus_offset_3327_symbol; -- transition assign_stmt_14/array_obj_ref_13_root_address_calculated
      array_obj_ref_13_word_address_calculated_3288_symbol <= array_obj_ref_13_word_addrgen_3332_symbol; -- transition assign_stmt_14/array_obj_ref_13_word_address_calculated
      array_obj_ref_13_indices_scaled_3289_symbol <= array_obj_ref_13_index_scale_0_3317_symbol; -- transition assign_stmt_14/array_obj_ref_13_indices_scaled
      array_obj_ref_13_offset_calculated_3290_symbol <= array_obj_ref_13_add_indices_3322_symbol; -- transition assign_stmt_14/array_obj_ref_13_offset_calculated
      array_obj_ref_13_index_computed_0_3291_symbol <= binary_12_complete_3305_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_computed_0
      array_obj_ref_13_index_resized_0_3292_symbol <= array_obj_ref_13_index_resize_0_3312_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_resized_0
      binary_12_active_x_x3293_block : Block -- non-trivial join transition assign_stmt_14/binary_12_active_ 
        signal binary_12_active_x_x3293_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_12_active_x_x3293_predecessors(0) <= binary_12_trigger_x_x3294_symbol;
        binary_12_active_x_x3293_predecessors(1) <= binary_10_complete_3298_symbol;
        binary_12_active_x_x3293_join: join -- 
          port map( -- 
            preds => binary_12_active_x_x3293_predecessors,
            symbol_out => binary_12_active_x_x3293_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_14/binary_12_active_
      binary_12_trigger_x_x3294_symbol <= Xentry_3281_symbol; -- transition assign_stmt_14/binary_12_trigger_
      binary_10_active_x_x3295_block : Block -- non-trivial join transition assign_stmt_14/binary_10_active_ 
        signal binary_10_active_x_x3295_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_10_active_x_x3295_predecessors(0) <= binary_10_trigger_x_x3296_symbol;
        binary_10_active_x_x3295_predecessors(1) <= simple_obj_ref_8_complete_3297_symbol;
        binary_10_active_x_x3295_join: join -- 
          port map( -- 
            preds => binary_10_active_x_x3295_predecessors,
            symbol_out => binary_10_active_x_x3295_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_14/binary_10_active_
      binary_10_trigger_x_x3296_symbol <= Xentry_3281_symbol; -- transition assign_stmt_14/binary_10_trigger_
      simple_obj_ref_8_complete_3297_symbol <= Xentry_3281_symbol; -- transition assign_stmt_14/simple_obj_ref_8_complete
      binary_10_complete_3298: Block -- assign_stmt_14/binary_10_complete 
        signal binary_10_complete_3298_start: Boolean;
        signal Xentry_3299_symbol: Boolean;
        signal Xexit_3300_symbol: Boolean;
        signal rr_3301_symbol : Boolean;
        signal ra_3302_symbol : Boolean;
        signal cr_3303_symbol : Boolean;
        signal ca_3304_symbol : Boolean;
        -- 
      begin -- 
        binary_10_complete_3298_start <= binary_10_active_x_x3295_symbol; -- control passed to block
        Xentry_3299_symbol  <= binary_10_complete_3298_start; -- transition assign_stmt_14/binary_10_complete/$entry
        rr_3301_symbol <= Xentry_3299_symbol; -- transition assign_stmt_14/binary_10_complete/rr
        binary_10_inst_req_0 <= rr_3301_symbol; -- link to DP
        ra_3302_symbol <= binary_10_inst_ack_0; -- transition assign_stmt_14/binary_10_complete/ra
        cr_3303_symbol <= ra_3302_symbol; -- transition assign_stmt_14/binary_10_complete/cr
        binary_10_inst_req_1 <= cr_3303_symbol; -- link to DP
        ca_3304_symbol <= binary_10_inst_ack_1; -- transition assign_stmt_14/binary_10_complete/ca
        Xexit_3300_symbol <= ca_3304_symbol; -- transition assign_stmt_14/binary_10_complete/$exit
        binary_10_complete_3298_symbol <= Xexit_3300_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/binary_10_complete
      binary_12_complete_3305: Block -- assign_stmt_14/binary_12_complete 
        signal binary_12_complete_3305_start: Boolean;
        signal Xentry_3306_symbol: Boolean;
        signal Xexit_3307_symbol: Boolean;
        signal rr_3308_symbol : Boolean;
        signal ra_3309_symbol : Boolean;
        signal cr_3310_symbol : Boolean;
        signal ca_3311_symbol : Boolean;
        -- 
      begin -- 
        binary_12_complete_3305_start <= binary_12_active_x_x3293_symbol; -- control passed to block
        Xentry_3306_symbol  <= binary_12_complete_3305_start; -- transition assign_stmt_14/binary_12_complete/$entry
        rr_3308_symbol <= Xentry_3306_symbol; -- transition assign_stmt_14/binary_12_complete/rr
        binary_12_inst_req_0 <= rr_3308_symbol; -- link to DP
        ra_3309_symbol <= binary_12_inst_ack_0; -- transition assign_stmt_14/binary_12_complete/ra
        cr_3310_symbol <= ra_3309_symbol; -- transition assign_stmt_14/binary_12_complete/cr
        binary_12_inst_req_1 <= cr_3310_symbol; -- link to DP
        ca_3311_symbol <= binary_12_inst_ack_1; -- transition assign_stmt_14/binary_12_complete/ca
        Xexit_3307_symbol <= ca_3311_symbol; -- transition assign_stmt_14/binary_12_complete/$exit
        binary_12_complete_3305_symbol <= Xexit_3307_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/binary_12_complete
      array_obj_ref_13_index_resize_0_3312: Block -- assign_stmt_14/array_obj_ref_13_index_resize_0 
        signal array_obj_ref_13_index_resize_0_3312_start: Boolean;
        signal Xentry_3313_symbol: Boolean;
        signal Xexit_3314_symbol: Boolean;
        signal index_resize_req_3315_symbol : Boolean;
        signal index_resize_ack_3316_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_index_resize_0_3312_start <= array_obj_ref_13_index_computed_0_3291_symbol; -- control passed to block
        Xentry_3313_symbol  <= array_obj_ref_13_index_resize_0_3312_start; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/$entry
        index_resize_req_3315_symbol <= Xentry_3313_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/index_resize_req
        array_obj_ref_13_index_0_resize_req_0 <= index_resize_req_3315_symbol; -- link to DP
        index_resize_ack_3316_symbol <= array_obj_ref_13_index_0_resize_ack_0; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/index_resize_ack
        Xexit_3314_symbol <= index_resize_ack_3316_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/$exit
        array_obj_ref_13_index_resize_0_3312_symbol <= Xexit_3314_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_index_resize_0
      array_obj_ref_13_index_scale_0_3317: Block -- assign_stmt_14/array_obj_ref_13_index_scale_0 
        signal array_obj_ref_13_index_scale_0_3317_start: Boolean;
        signal Xentry_3318_symbol: Boolean;
        signal Xexit_3319_symbol: Boolean;
        signal scale_rename_req_3320_symbol : Boolean;
        signal scale_rename_ack_3321_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_index_scale_0_3317_start <= array_obj_ref_13_index_resized_0_3292_symbol; -- control passed to block
        Xentry_3318_symbol  <= array_obj_ref_13_index_scale_0_3317_start; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/$entry
        scale_rename_req_3320_symbol <= Xentry_3318_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/scale_rename_req
        array_obj_ref_13_index_0_rename_req_0 <= scale_rename_req_3320_symbol; -- link to DP
        scale_rename_ack_3321_symbol <= array_obj_ref_13_index_0_rename_ack_0; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/scale_rename_ack
        Xexit_3319_symbol <= scale_rename_ack_3321_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/$exit
        array_obj_ref_13_index_scale_0_3317_symbol <= Xexit_3319_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_index_scale_0
      array_obj_ref_13_add_indices_3322: Block -- assign_stmt_14/array_obj_ref_13_add_indices 
        signal array_obj_ref_13_add_indices_3322_start: Boolean;
        signal Xentry_3323_symbol: Boolean;
        signal Xexit_3324_symbol: Boolean;
        signal final_index_req_3325_symbol : Boolean;
        signal final_index_ack_3326_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_add_indices_3322_start <= array_obj_ref_13_indices_scaled_3289_symbol; -- control passed to block
        Xentry_3323_symbol  <= array_obj_ref_13_add_indices_3322_start; -- transition assign_stmt_14/array_obj_ref_13_add_indices/$entry
        final_index_req_3325_symbol <= Xentry_3323_symbol; -- transition assign_stmt_14/array_obj_ref_13_add_indices/final_index_req
        array_obj_ref_13_offset_inst_req_0 <= final_index_req_3325_symbol; -- link to DP
        final_index_ack_3326_symbol <= array_obj_ref_13_offset_inst_ack_0; -- transition assign_stmt_14/array_obj_ref_13_add_indices/final_index_ack
        Xexit_3324_symbol <= final_index_ack_3326_symbol; -- transition assign_stmt_14/array_obj_ref_13_add_indices/$exit
        array_obj_ref_13_add_indices_3322_symbol <= Xexit_3324_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_add_indices
      array_obj_ref_13_base_plus_offset_3327: Block -- assign_stmt_14/array_obj_ref_13_base_plus_offset 
        signal array_obj_ref_13_base_plus_offset_3327_start: Boolean;
        signal Xentry_3328_symbol: Boolean;
        signal Xexit_3329_symbol: Boolean;
        signal sum_rename_req_3330_symbol : Boolean;
        signal sum_rename_ack_3331_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_base_plus_offset_3327_start <= array_obj_ref_13_offset_calculated_3290_symbol; -- control passed to block
        Xentry_3328_symbol  <= array_obj_ref_13_base_plus_offset_3327_start; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/$entry
        sum_rename_req_3330_symbol <= Xentry_3328_symbol; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/sum_rename_req
        array_obj_ref_13_root_address_inst_req_0 <= sum_rename_req_3330_symbol; -- link to DP
        sum_rename_ack_3331_symbol <= array_obj_ref_13_root_address_inst_ack_0; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/sum_rename_ack
        Xexit_3329_symbol <= sum_rename_ack_3331_symbol; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/$exit
        array_obj_ref_13_base_plus_offset_3327_symbol <= Xexit_3329_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_base_plus_offset
      array_obj_ref_13_word_addrgen_3332: Block -- assign_stmt_14/array_obj_ref_13_word_addrgen 
        signal array_obj_ref_13_word_addrgen_3332_start: Boolean;
        signal Xentry_3333_symbol: Boolean;
        signal Xexit_3334_symbol: Boolean;
        signal root_rename_req_3335_symbol : Boolean;
        signal root_rename_ack_3336_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_word_addrgen_3332_start <= array_obj_ref_13_root_address_calculated_3287_symbol; -- control passed to block
        Xentry_3333_symbol  <= array_obj_ref_13_word_addrgen_3332_start; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/$entry
        root_rename_req_3335_symbol <= Xentry_3333_symbol; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/root_rename_req
        array_obj_ref_13_addr_0_req_0 <= root_rename_req_3335_symbol; -- link to DP
        root_rename_ack_3336_symbol <= array_obj_ref_13_addr_0_ack_0; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/root_rename_ack
        Xexit_3334_symbol <= root_rename_ack_3336_symbol; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/$exit
        array_obj_ref_13_word_addrgen_3332_symbol <= Xexit_3334_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_word_addrgen
      array_obj_ref_13_request_3337: Block -- assign_stmt_14/array_obj_ref_13_request 
        signal array_obj_ref_13_request_3337_start: Boolean;
        signal Xentry_3338_symbol: Boolean;
        signal Xexit_3339_symbol: Boolean;
        signal word_access_3340_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_request_3337_start <= array_obj_ref_13_trigger_x_x3285_symbol; -- control passed to block
        Xentry_3338_symbol  <= array_obj_ref_13_request_3337_start; -- transition assign_stmt_14/array_obj_ref_13_request/$entry
        word_access_3340: Block -- assign_stmt_14/array_obj_ref_13_request/word_access 
          signal word_access_3340_start: Boolean;
          signal Xentry_3341_symbol: Boolean;
          signal Xexit_3342_symbol: Boolean;
          signal word_access_0_3343_symbol : Boolean;
          -- 
        begin -- 
          word_access_3340_start <= Xentry_3338_symbol; -- control passed to block
          Xentry_3341_symbol  <= word_access_3340_start; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/$entry
          word_access_0_3343: Block -- assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0 
            signal word_access_0_3343_start: Boolean;
            signal Xentry_3344_symbol: Boolean;
            signal Xexit_3345_symbol: Boolean;
            signal rr_3346_symbol : Boolean;
            signal ra_3347_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_3343_start <= Xentry_3341_symbol; -- control passed to block
            Xentry_3344_symbol  <= word_access_0_3343_start; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/$entry
            rr_3346_symbol <= Xentry_3344_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/rr
            array_obj_ref_13_load_0_req_0 <= rr_3346_symbol; -- link to DP
            ra_3347_symbol <= array_obj_ref_13_load_0_ack_0; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/ra
            Xexit_3345_symbol <= ra_3347_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/$exit
            word_access_0_3343_symbol <= Xexit_3345_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0
          Xexit_3342_symbol <= word_access_0_3343_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/$exit
          word_access_3340_symbol <= Xexit_3342_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_14/array_obj_ref_13_request/word_access
        Xexit_3339_symbol <= word_access_3340_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/$exit
        array_obj_ref_13_request_3337_symbol <= Xexit_3339_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_request
      array_obj_ref_13_complete_3348: Block -- assign_stmt_14/array_obj_ref_13_complete 
        signal array_obj_ref_13_complete_3348_start: Boolean;
        signal Xentry_3349_symbol: Boolean;
        signal Xexit_3350_symbol: Boolean;
        signal word_access_3351_symbol : Boolean;
        signal merge_req_3359_symbol : Boolean;
        signal merge_ack_3360_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_complete_3348_start <= array_obj_ref_13_active_x_x3286_symbol; -- control passed to block
        Xentry_3349_symbol  <= array_obj_ref_13_complete_3348_start; -- transition assign_stmt_14/array_obj_ref_13_complete/$entry
        word_access_3351: Block -- assign_stmt_14/array_obj_ref_13_complete/word_access 
          signal word_access_3351_start: Boolean;
          signal Xentry_3352_symbol: Boolean;
          signal Xexit_3353_symbol: Boolean;
          signal word_access_0_3354_symbol : Boolean;
          -- 
        begin -- 
          word_access_3351_start <= Xentry_3349_symbol; -- control passed to block
          Xentry_3352_symbol  <= word_access_3351_start; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/$entry
          word_access_0_3354: Block -- assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0 
            signal word_access_0_3354_start: Boolean;
            signal Xentry_3355_symbol: Boolean;
            signal Xexit_3356_symbol: Boolean;
            signal cr_3357_symbol : Boolean;
            signal ca_3358_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_3354_start <= Xentry_3352_symbol; -- control passed to block
            Xentry_3355_symbol  <= word_access_0_3354_start; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/$entry
            cr_3357_symbol <= Xentry_3355_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/cr
            array_obj_ref_13_load_0_req_1 <= cr_3357_symbol; -- link to DP
            ca_3358_symbol <= array_obj_ref_13_load_0_ack_1; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/ca
            Xexit_3356_symbol <= ca_3358_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/$exit
            word_access_0_3354_symbol <= Xexit_3356_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0
          Xexit_3353_symbol <= word_access_0_3354_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/$exit
          word_access_3351_symbol <= Xexit_3353_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_14/array_obj_ref_13_complete/word_access
        merge_req_3359_symbol <= word_access_3351_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/merge_req
        array_obj_ref_13_gather_scatter_req_0 <= merge_req_3359_symbol; -- link to DP
        merge_ack_3360_symbol <= array_obj_ref_13_gather_scatter_ack_0; -- transition assign_stmt_14/array_obj_ref_13_complete/merge_ack
        Xexit_3350_symbol <= merge_ack_3360_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/$exit
        array_obj_ref_13_complete_3348_symbol <= Xexit_3350_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_complete
      Xexit_3282_symbol <= assign_stmt_14_completed_x_x3284_symbol; -- transition assign_stmt_14/$exit
      assign_stmt_14_3280_symbol <= Xexit_3282_symbol; -- control passed from block 
      -- 
    end Block; -- assign_stmt_14
    Xexit_3279_symbol <= assign_stmt_14_3280_symbol; -- transition $exit
    fin  <=  '1' when Xexit_3279_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_13_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_13_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_word_offset_0 : std_logic_vector(0 downto 0);
    signal binary_10_wire : std_logic_vector(31 downto 0);
    signal binary_12_resized : std_logic_vector(0 downto 0);
    signal binary_12_scaled : std_logic_vector(0 downto 0);
    signal binary_12_wire : std_logic_vector(31 downto 0);
    signal expr_11_wire_constant : std_logic_vector(31 downto 0);
    signal expr_9_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_13_offset_scale_factor_0 <= "1";
    array_obj_ref_13_resized_base_address <= "0";
    array_obj_ref_13_word_offset_0 <= "0";
    expr_11_wire_constant <= "00000000000000000000000000000000";
    expr_9_wire_constant <= "00000000000000000000000000000001";
    array_obj_ref_13_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 1) -- 
      port map( din => binary_12_wire, dout => binary_12_resized, req => array_obj_ref_13_index_0_resize_req_0, ack => array_obj_ref_13_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_13_offset_inst: RegisterBase generic map(in_data_width => 1,out_data_width => 1) -- 
      port map( din => binary_12_scaled, dout => array_obj_ref_13_final_offset, req => array_obj_ref_13_offset_inst_req_0, ack => array_obj_ref_13_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_13_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_13_addr_0_ack_0 <= array_obj_ref_13_addr_0_req_0;
      aggregated_sig <= array_obj_ref_13_root_address;
      array_obj_ref_13_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_13_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_13_gather_scatter_ack_0 <= array_obj_ref_13_gather_scatter_req_0;
      aggregated_sig <= array_obj_ref_13_data_0;
      data <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_13_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_13_index_0_rename_ack_0 <= array_obj_ref_13_index_0_rename_req_0;
      aggregated_sig <= binary_12_resized;
      binary_12_scaled <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_13_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_13_root_address_inst_ack_0 <= array_obj_ref_13_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_13_final_offset;
      array_obj_ref_13_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    -- shared split operator group (0) : binary_10_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= address;
      binary_10_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_10_inst_req_0,
          ackL => binary_10_inst_ack_0,
          reqR => binary_10_inst_req_1,
          ackR => binary_10_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_12_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_10_wire;
      binary_12_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_12_inst_req_0,
          ackL => binary_12_inst_ack_0,
          reqR => binary_12_inst_req_1,
          ackR => binary_12_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared load operator group (0) : array_obj_ref_13_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_13_load_0_req_0;
      array_obj_ref_13_load_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_13_load_0_req_1;
      array_obj_ref_13_load_0_ack_1 <= ackR(0);
      data_in <= array_obj_ref_13_word_address_0;
      array_obj_ref_13_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(7 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity mem_store_x_x is -- 
  port ( -- 
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(7 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity mem_store_x_x;
architecture Default of mem_store_x_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_24_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_24_gather_scatter_req_0 : boolean;
  signal binary_21_inst_req_1 : boolean;
  signal binary_21_inst_ack_1 : boolean;
  signal array_obj_ref_24_gather_scatter_ack_0 : boolean;
  signal binary_21_inst_req_0 : boolean;
  signal binary_21_inst_ack_0 : boolean;
  signal binary_23_inst_req_0 : boolean;
  signal array_obj_ref_24_store_0_req_1 : boolean;
  signal binary_23_inst_req_1 : boolean;
  signal binary_23_inst_ack_0 : boolean;
  signal array_obj_ref_24_store_0_ack_1 : boolean;
  signal array_obj_ref_24_root_address_inst_req_0 : boolean;
  signal array_obj_ref_24_addr_0_req_0 : boolean;
  signal array_obj_ref_24_addr_0_ack_0 : boolean;
  signal array_obj_ref_24_store_0_ack_0 : boolean;
  signal array_obj_ref_24_store_0_req_0 : boolean;
  signal binary_23_inst_ack_1 : boolean;
  signal array_obj_ref_24_index_0_resize_req_0 : boolean;
  signal array_obj_ref_24_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_24_index_0_rename_req_0 : boolean;
  signal array_obj_ref_24_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_24_offset_inst_req_0 : boolean;
  signal array_obj_ref_24_offset_inst_ack_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  mem_store_x_xx_xCP_3361: Block -- control-path 
    signal mem_store_x_xx_xCP_3361_start: Boolean;
    signal Xentry_3362_symbol: Boolean;
    signal Xexit_3363_symbol: Boolean;
    signal assign_stmt_26_3364_symbol : Boolean;
    -- 
  begin -- 
    mem_store_x_xx_xCP_3361_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_3362_symbol  <= mem_store_x_xx_xCP_3361_start; -- transition $entry
    assign_stmt_26_3364: Block -- assign_stmt_26 
      signal assign_stmt_26_3364_start: Boolean;
      signal Xentry_3365_symbol: Boolean;
      signal Xexit_3366_symbol: Boolean;
      signal assign_stmt_26_active_x_x3367_symbol : Boolean;
      signal assign_stmt_26_completed_x_x3368_symbol : Boolean;
      signal simple_obj_ref_25_complete_3369_symbol : Boolean;
      signal array_obj_ref_24_trigger_x_x3370_symbol : Boolean;
      signal array_obj_ref_24_active_x_x3371_symbol : Boolean;
      signal array_obj_ref_24_root_address_calculated_3372_symbol : Boolean;
      signal array_obj_ref_24_word_address_calculated_3373_symbol : Boolean;
      signal array_obj_ref_24_indices_scaled_3374_symbol : Boolean;
      signal array_obj_ref_24_offset_calculated_3375_symbol : Boolean;
      signal array_obj_ref_24_index_computed_0_3376_symbol : Boolean;
      signal array_obj_ref_24_index_resized_0_3377_symbol : Boolean;
      signal binary_23_active_x_x3378_symbol : Boolean;
      signal binary_23_trigger_x_x3379_symbol : Boolean;
      signal binary_21_active_x_x3380_symbol : Boolean;
      signal binary_21_trigger_x_x3381_symbol : Boolean;
      signal simple_obj_ref_19_complete_3382_symbol : Boolean;
      signal binary_21_complete_3383_symbol : Boolean;
      signal binary_23_complete_3390_symbol : Boolean;
      signal array_obj_ref_24_index_resize_0_3397_symbol : Boolean;
      signal array_obj_ref_24_index_scale_0_3402_symbol : Boolean;
      signal array_obj_ref_24_add_indices_3407_symbol : Boolean;
      signal array_obj_ref_24_base_plus_offset_3412_symbol : Boolean;
      signal array_obj_ref_24_word_addrgen_3417_symbol : Boolean;
      signal array_obj_ref_24_request_3422_symbol : Boolean;
      signal array_obj_ref_24_complete_3435_symbol : Boolean;
      -- 
    begin -- 
      assign_stmt_26_3364_start <= Xentry_3362_symbol; -- control passed to block
      Xentry_3365_symbol  <= assign_stmt_26_3364_start; -- transition assign_stmt_26/$entry
      assign_stmt_26_active_x_x3367_symbol <= simple_obj_ref_25_complete_3369_symbol; -- transition assign_stmt_26/assign_stmt_26_active_
      assign_stmt_26_completed_x_x3368_symbol <= array_obj_ref_24_complete_3435_symbol; -- transition assign_stmt_26/assign_stmt_26_completed_
      simple_obj_ref_25_complete_3369_symbol <= Xentry_3365_symbol; -- transition assign_stmt_26/simple_obj_ref_25_complete
      array_obj_ref_24_trigger_x_x3370_block : Block -- non-trivial join transition assign_stmt_26/array_obj_ref_24_trigger_ 
        signal array_obj_ref_24_trigger_x_x3370_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        array_obj_ref_24_trigger_x_x3370_predecessors(0) <= array_obj_ref_24_word_address_calculated_3373_symbol;
        array_obj_ref_24_trigger_x_x3370_predecessors(1) <= assign_stmt_26_active_x_x3367_symbol;
        array_obj_ref_24_trigger_x_x3370_join: join -- 
          port map( -- 
            preds => array_obj_ref_24_trigger_x_x3370_predecessors,
            symbol_out => array_obj_ref_24_trigger_x_x3370_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_26/array_obj_ref_24_trigger_
      array_obj_ref_24_active_x_x3371_symbol <= array_obj_ref_24_request_3422_symbol; -- transition assign_stmt_26/array_obj_ref_24_active_
      array_obj_ref_24_root_address_calculated_3372_symbol <= array_obj_ref_24_base_plus_offset_3412_symbol; -- transition assign_stmt_26/array_obj_ref_24_root_address_calculated
      array_obj_ref_24_word_address_calculated_3373_symbol <= array_obj_ref_24_word_addrgen_3417_symbol; -- transition assign_stmt_26/array_obj_ref_24_word_address_calculated
      array_obj_ref_24_indices_scaled_3374_symbol <= array_obj_ref_24_index_scale_0_3402_symbol; -- transition assign_stmt_26/array_obj_ref_24_indices_scaled
      array_obj_ref_24_offset_calculated_3375_symbol <= array_obj_ref_24_add_indices_3407_symbol; -- transition assign_stmt_26/array_obj_ref_24_offset_calculated
      array_obj_ref_24_index_computed_0_3376_symbol <= binary_23_complete_3390_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_computed_0
      array_obj_ref_24_index_resized_0_3377_symbol <= array_obj_ref_24_index_resize_0_3397_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_resized_0
      binary_23_active_x_x3378_block : Block -- non-trivial join transition assign_stmt_26/binary_23_active_ 
        signal binary_23_active_x_x3378_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_23_active_x_x3378_predecessors(0) <= binary_23_trigger_x_x3379_symbol;
        binary_23_active_x_x3378_predecessors(1) <= binary_21_complete_3383_symbol;
        binary_23_active_x_x3378_join: join -- 
          port map( -- 
            preds => binary_23_active_x_x3378_predecessors,
            symbol_out => binary_23_active_x_x3378_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_26/binary_23_active_
      binary_23_trigger_x_x3379_symbol <= Xentry_3365_symbol; -- transition assign_stmt_26/binary_23_trigger_
      binary_21_active_x_x3380_block : Block -- non-trivial join transition assign_stmt_26/binary_21_active_ 
        signal binary_21_active_x_x3380_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_21_active_x_x3380_predecessors(0) <= binary_21_trigger_x_x3381_symbol;
        binary_21_active_x_x3380_predecessors(1) <= simple_obj_ref_19_complete_3382_symbol;
        binary_21_active_x_x3380_join: join -- 
          port map( -- 
            preds => binary_21_active_x_x3380_predecessors,
            symbol_out => binary_21_active_x_x3380_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_26/binary_21_active_
      binary_21_trigger_x_x3381_symbol <= Xentry_3365_symbol; -- transition assign_stmt_26/binary_21_trigger_
      simple_obj_ref_19_complete_3382_symbol <= Xentry_3365_symbol; -- transition assign_stmt_26/simple_obj_ref_19_complete
      binary_21_complete_3383: Block -- assign_stmt_26/binary_21_complete 
        signal binary_21_complete_3383_start: Boolean;
        signal Xentry_3384_symbol: Boolean;
        signal Xexit_3385_symbol: Boolean;
        signal rr_3386_symbol : Boolean;
        signal ra_3387_symbol : Boolean;
        signal cr_3388_symbol : Boolean;
        signal ca_3389_symbol : Boolean;
        -- 
      begin -- 
        binary_21_complete_3383_start <= binary_21_active_x_x3380_symbol; -- control passed to block
        Xentry_3384_symbol  <= binary_21_complete_3383_start; -- transition assign_stmt_26/binary_21_complete/$entry
        rr_3386_symbol <= Xentry_3384_symbol; -- transition assign_stmt_26/binary_21_complete/rr
        binary_21_inst_req_0 <= rr_3386_symbol; -- link to DP
        ra_3387_symbol <= binary_21_inst_ack_0; -- transition assign_stmt_26/binary_21_complete/ra
        cr_3388_symbol <= ra_3387_symbol; -- transition assign_stmt_26/binary_21_complete/cr
        binary_21_inst_req_1 <= cr_3388_symbol; -- link to DP
        ca_3389_symbol <= binary_21_inst_ack_1; -- transition assign_stmt_26/binary_21_complete/ca
        Xexit_3385_symbol <= ca_3389_symbol; -- transition assign_stmt_26/binary_21_complete/$exit
        binary_21_complete_3383_symbol <= Xexit_3385_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/binary_21_complete
      binary_23_complete_3390: Block -- assign_stmt_26/binary_23_complete 
        signal binary_23_complete_3390_start: Boolean;
        signal Xentry_3391_symbol: Boolean;
        signal Xexit_3392_symbol: Boolean;
        signal rr_3393_symbol : Boolean;
        signal ra_3394_symbol : Boolean;
        signal cr_3395_symbol : Boolean;
        signal ca_3396_symbol : Boolean;
        -- 
      begin -- 
        binary_23_complete_3390_start <= binary_23_active_x_x3378_symbol; -- control passed to block
        Xentry_3391_symbol  <= binary_23_complete_3390_start; -- transition assign_stmt_26/binary_23_complete/$entry
        rr_3393_symbol <= Xentry_3391_symbol; -- transition assign_stmt_26/binary_23_complete/rr
        binary_23_inst_req_0 <= rr_3393_symbol; -- link to DP
        ra_3394_symbol <= binary_23_inst_ack_0; -- transition assign_stmt_26/binary_23_complete/ra
        cr_3395_symbol <= ra_3394_symbol; -- transition assign_stmt_26/binary_23_complete/cr
        binary_23_inst_req_1 <= cr_3395_symbol; -- link to DP
        ca_3396_symbol <= binary_23_inst_ack_1; -- transition assign_stmt_26/binary_23_complete/ca
        Xexit_3392_symbol <= ca_3396_symbol; -- transition assign_stmt_26/binary_23_complete/$exit
        binary_23_complete_3390_symbol <= Xexit_3392_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/binary_23_complete
      array_obj_ref_24_index_resize_0_3397: Block -- assign_stmt_26/array_obj_ref_24_index_resize_0 
        signal array_obj_ref_24_index_resize_0_3397_start: Boolean;
        signal Xentry_3398_symbol: Boolean;
        signal Xexit_3399_symbol: Boolean;
        signal index_resize_req_3400_symbol : Boolean;
        signal index_resize_ack_3401_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_index_resize_0_3397_start <= array_obj_ref_24_index_computed_0_3376_symbol; -- control passed to block
        Xentry_3398_symbol  <= array_obj_ref_24_index_resize_0_3397_start; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/$entry
        index_resize_req_3400_symbol <= Xentry_3398_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/index_resize_req
        array_obj_ref_24_index_0_resize_req_0 <= index_resize_req_3400_symbol; -- link to DP
        index_resize_ack_3401_symbol <= array_obj_ref_24_index_0_resize_ack_0; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/index_resize_ack
        Xexit_3399_symbol <= index_resize_ack_3401_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/$exit
        array_obj_ref_24_index_resize_0_3397_symbol <= Xexit_3399_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_index_resize_0
      array_obj_ref_24_index_scale_0_3402: Block -- assign_stmt_26/array_obj_ref_24_index_scale_0 
        signal array_obj_ref_24_index_scale_0_3402_start: Boolean;
        signal Xentry_3403_symbol: Boolean;
        signal Xexit_3404_symbol: Boolean;
        signal scale_rename_req_3405_symbol : Boolean;
        signal scale_rename_ack_3406_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_index_scale_0_3402_start <= array_obj_ref_24_index_resized_0_3377_symbol; -- control passed to block
        Xentry_3403_symbol  <= array_obj_ref_24_index_scale_0_3402_start; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/$entry
        scale_rename_req_3405_symbol <= Xentry_3403_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/scale_rename_req
        array_obj_ref_24_index_0_rename_req_0 <= scale_rename_req_3405_symbol; -- link to DP
        scale_rename_ack_3406_symbol <= array_obj_ref_24_index_0_rename_ack_0; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/scale_rename_ack
        Xexit_3404_symbol <= scale_rename_ack_3406_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/$exit
        array_obj_ref_24_index_scale_0_3402_symbol <= Xexit_3404_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_index_scale_0
      array_obj_ref_24_add_indices_3407: Block -- assign_stmt_26/array_obj_ref_24_add_indices 
        signal array_obj_ref_24_add_indices_3407_start: Boolean;
        signal Xentry_3408_symbol: Boolean;
        signal Xexit_3409_symbol: Boolean;
        signal final_index_req_3410_symbol : Boolean;
        signal final_index_ack_3411_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_add_indices_3407_start <= array_obj_ref_24_indices_scaled_3374_symbol; -- control passed to block
        Xentry_3408_symbol  <= array_obj_ref_24_add_indices_3407_start; -- transition assign_stmt_26/array_obj_ref_24_add_indices/$entry
        final_index_req_3410_symbol <= Xentry_3408_symbol; -- transition assign_stmt_26/array_obj_ref_24_add_indices/final_index_req
        array_obj_ref_24_offset_inst_req_0 <= final_index_req_3410_symbol; -- link to DP
        final_index_ack_3411_symbol <= array_obj_ref_24_offset_inst_ack_0; -- transition assign_stmt_26/array_obj_ref_24_add_indices/final_index_ack
        Xexit_3409_symbol <= final_index_ack_3411_symbol; -- transition assign_stmt_26/array_obj_ref_24_add_indices/$exit
        array_obj_ref_24_add_indices_3407_symbol <= Xexit_3409_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_add_indices
      array_obj_ref_24_base_plus_offset_3412: Block -- assign_stmt_26/array_obj_ref_24_base_plus_offset 
        signal array_obj_ref_24_base_plus_offset_3412_start: Boolean;
        signal Xentry_3413_symbol: Boolean;
        signal Xexit_3414_symbol: Boolean;
        signal sum_rename_req_3415_symbol : Boolean;
        signal sum_rename_ack_3416_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_base_plus_offset_3412_start <= array_obj_ref_24_offset_calculated_3375_symbol; -- control passed to block
        Xentry_3413_symbol  <= array_obj_ref_24_base_plus_offset_3412_start; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/$entry
        sum_rename_req_3415_symbol <= Xentry_3413_symbol; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/sum_rename_req
        array_obj_ref_24_root_address_inst_req_0 <= sum_rename_req_3415_symbol; -- link to DP
        sum_rename_ack_3416_symbol <= array_obj_ref_24_root_address_inst_ack_0; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/sum_rename_ack
        Xexit_3414_symbol <= sum_rename_ack_3416_symbol; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/$exit
        array_obj_ref_24_base_plus_offset_3412_symbol <= Xexit_3414_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_base_plus_offset
      array_obj_ref_24_word_addrgen_3417: Block -- assign_stmt_26/array_obj_ref_24_word_addrgen 
        signal array_obj_ref_24_word_addrgen_3417_start: Boolean;
        signal Xentry_3418_symbol: Boolean;
        signal Xexit_3419_symbol: Boolean;
        signal root_rename_req_3420_symbol : Boolean;
        signal root_rename_ack_3421_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_word_addrgen_3417_start <= array_obj_ref_24_root_address_calculated_3372_symbol; -- control passed to block
        Xentry_3418_symbol  <= array_obj_ref_24_word_addrgen_3417_start; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/$entry
        root_rename_req_3420_symbol <= Xentry_3418_symbol; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/root_rename_req
        array_obj_ref_24_addr_0_req_0 <= root_rename_req_3420_symbol; -- link to DP
        root_rename_ack_3421_symbol <= array_obj_ref_24_addr_0_ack_0; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/root_rename_ack
        Xexit_3419_symbol <= root_rename_ack_3421_symbol; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/$exit
        array_obj_ref_24_word_addrgen_3417_symbol <= Xexit_3419_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_word_addrgen
      array_obj_ref_24_request_3422: Block -- assign_stmt_26/array_obj_ref_24_request 
        signal array_obj_ref_24_request_3422_start: Boolean;
        signal Xentry_3423_symbol: Boolean;
        signal Xexit_3424_symbol: Boolean;
        signal split_req_3425_symbol : Boolean;
        signal split_ack_3426_symbol : Boolean;
        signal word_access_3427_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_request_3422_start <= array_obj_ref_24_trigger_x_x3370_symbol; -- control passed to block
        Xentry_3423_symbol  <= array_obj_ref_24_request_3422_start; -- transition assign_stmt_26/array_obj_ref_24_request/$entry
        split_req_3425_symbol <= Xentry_3423_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/split_req
        array_obj_ref_24_gather_scatter_req_0 <= split_req_3425_symbol; -- link to DP
        split_ack_3426_symbol <= array_obj_ref_24_gather_scatter_ack_0; -- transition assign_stmt_26/array_obj_ref_24_request/split_ack
        word_access_3427: Block -- assign_stmt_26/array_obj_ref_24_request/word_access 
          signal word_access_3427_start: Boolean;
          signal Xentry_3428_symbol: Boolean;
          signal Xexit_3429_symbol: Boolean;
          signal word_access_0_3430_symbol : Boolean;
          -- 
        begin -- 
          word_access_3427_start <= split_ack_3426_symbol; -- control passed to block
          Xentry_3428_symbol  <= word_access_3427_start; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/$entry
          word_access_0_3430: Block -- assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0 
            signal word_access_0_3430_start: Boolean;
            signal Xentry_3431_symbol: Boolean;
            signal Xexit_3432_symbol: Boolean;
            signal rr_3433_symbol : Boolean;
            signal ra_3434_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_3430_start <= Xentry_3428_symbol; -- control passed to block
            Xentry_3431_symbol  <= word_access_0_3430_start; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/$entry
            rr_3433_symbol <= Xentry_3431_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/rr
            array_obj_ref_24_store_0_req_0 <= rr_3433_symbol; -- link to DP
            ra_3434_symbol <= array_obj_ref_24_store_0_ack_0; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/ra
            Xexit_3432_symbol <= ra_3434_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/$exit
            word_access_0_3430_symbol <= Xexit_3432_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0
          Xexit_3429_symbol <= word_access_0_3430_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/$exit
          word_access_3427_symbol <= Xexit_3429_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_26/array_obj_ref_24_request/word_access
        Xexit_3424_symbol <= word_access_3427_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/$exit
        array_obj_ref_24_request_3422_symbol <= Xexit_3424_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_request
      array_obj_ref_24_complete_3435: Block -- assign_stmt_26/array_obj_ref_24_complete 
        signal array_obj_ref_24_complete_3435_start: Boolean;
        signal Xentry_3436_symbol: Boolean;
        signal Xexit_3437_symbol: Boolean;
        signal word_access_3438_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_complete_3435_start <= array_obj_ref_24_active_x_x3371_symbol; -- control passed to block
        Xentry_3436_symbol  <= array_obj_ref_24_complete_3435_start; -- transition assign_stmt_26/array_obj_ref_24_complete/$entry
        word_access_3438: Block -- assign_stmt_26/array_obj_ref_24_complete/word_access 
          signal word_access_3438_start: Boolean;
          signal Xentry_3439_symbol: Boolean;
          signal Xexit_3440_symbol: Boolean;
          signal word_access_0_3441_symbol : Boolean;
          -- 
        begin -- 
          word_access_3438_start <= Xentry_3436_symbol; -- control passed to block
          Xentry_3439_symbol  <= word_access_3438_start; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/$entry
          word_access_0_3441: Block -- assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0 
            signal word_access_0_3441_start: Boolean;
            signal Xentry_3442_symbol: Boolean;
            signal Xexit_3443_symbol: Boolean;
            signal cr_3444_symbol : Boolean;
            signal ca_3445_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_3441_start <= Xentry_3439_symbol; -- control passed to block
            Xentry_3442_symbol  <= word_access_0_3441_start; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/$entry
            cr_3444_symbol <= Xentry_3442_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/cr
            array_obj_ref_24_store_0_req_1 <= cr_3444_symbol; -- link to DP
            ca_3445_symbol <= array_obj_ref_24_store_0_ack_1; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/ca
            Xexit_3443_symbol <= ca_3445_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/$exit
            word_access_0_3441_symbol <= Xexit_3443_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0
          Xexit_3440_symbol <= word_access_0_3441_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/$exit
          word_access_3438_symbol <= Xexit_3440_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_26/array_obj_ref_24_complete/word_access
        Xexit_3437_symbol <= word_access_3438_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/$exit
        array_obj_ref_24_complete_3435_symbol <= Xexit_3437_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_complete
      Xexit_3366_symbol <= assign_stmt_26_completed_x_x3368_symbol; -- transition assign_stmt_26/$exit
      assign_stmt_26_3364_symbol <= Xexit_3366_symbol; -- control passed from block 
      -- 
    end Block; -- assign_stmt_26
    Xexit_3363_symbol <= assign_stmt_26_3364_symbol; -- transition $exit
    fin  <=  '1' when Xexit_3363_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_24_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_24_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_word_offset_0 : std_logic_vector(0 downto 0);
    signal binary_21_wire : std_logic_vector(31 downto 0);
    signal binary_23_resized : std_logic_vector(0 downto 0);
    signal binary_23_scaled : std_logic_vector(0 downto 0);
    signal binary_23_wire : std_logic_vector(31 downto 0);
    signal expr_20_wire_constant : std_logic_vector(31 downto 0);
    signal expr_22_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_24_offset_scale_factor_0 <= "1";
    array_obj_ref_24_resized_base_address <= "0";
    array_obj_ref_24_word_offset_0 <= "0";
    expr_20_wire_constant <= "00000000000000000000000000000001";
    expr_22_wire_constant <= "00000000000000000000000000000000";
    array_obj_ref_24_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 1) -- 
      port map( din => binary_23_wire, dout => binary_23_resized, req => array_obj_ref_24_index_0_resize_req_0, ack => array_obj_ref_24_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_24_offset_inst: RegisterBase generic map(in_data_width => 1,out_data_width => 1) -- 
      port map( din => binary_23_scaled, dout => array_obj_ref_24_final_offset, req => array_obj_ref_24_offset_inst_req_0, ack => array_obj_ref_24_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_24_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_24_addr_0_ack_0 <= array_obj_ref_24_addr_0_req_0;
      aggregated_sig <= array_obj_ref_24_root_address;
      array_obj_ref_24_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_24_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_24_gather_scatter_ack_0 <= array_obj_ref_24_gather_scatter_req_0;
      aggregated_sig <= data;
      array_obj_ref_24_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_24_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_24_index_0_rename_ack_0 <= array_obj_ref_24_index_0_rename_req_0;
      aggregated_sig <= binary_23_resized;
      binary_23_scaled <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_24_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_24_root_address_inst_ack_0 <= array_obj_ref_24_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_24_final_offset;
      array_obj_ref_24_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    -- shared split operator group (0) : binary_21_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= address;
      binary_21_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_21_inst_req_0,
          ackL => binary_21_inst_ack_0,
          reqR => binary_21_inst_req_1,
          ackR => binary_21_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_23_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_21_wire;
      binary_23_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_23_inst_req_0,
          ackL => binary_23_inst_ack_0,
          reqR => binary_23_inst_req_1,
          ackR => binary_23_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_24_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_24_store_0_req_0;
      array_obj_ref_24_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_24_store_0_req_1;
      array_obj_ref_24_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_24_word_address_0;
      data_in <= array_obj_ref_24_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(7 downto 0),
          mtag => memory_space_0_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity output_module is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(47 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(23 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(7 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(7 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(23 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(3 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(23 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(11 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(3 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(3 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(11 downto 0);
    foo_out_pipe_read_req : out  std_logic_vector(0 downto 0);
    foo_out_pipe_read_ack : in   std_logic_vector(0 downto 0);
    foo_out_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_data_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity output_module;
architecture Default of output_module is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_535_store_0_req_1 : boolean;
  signal ptr_deref_540_load_1_ack_1 : boolean;
  signal ptr_deref_535_store_0_ack_1 : boolean;
  signal ptr_deref_535_store_1_ack_0 : boolean;
  signal array_obj_ref_545_base_resize_req_0 : boolean;
  signal type_cast_532_inst_ack_0 : boolean;
  signal ptr_deref_540_load_0_ack_1 : boolean;
  signal type_cast_532_inst_req_0 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal ptr_deref_540_load_3_req_1 : boolean;
  signal ptr_deref_540_load_2_req_1 : boolean;
  signal simple_obj_ref_527_inst_ack_0 : boolean;
  signal simple_obj_ref_527_inst_req_0 : boolean;
  signal ptr_deref_540_load_0_req_0 : boolean;
  signal ptr_deref_535_gather_scatter_req_0 : boolean;
  signal ptr_deref_540_load_3_ack_1 : boolean;
  signal ptr_deref_535_store_2_req_0 : boolean;
  signal ptr_deref_540_load_2_req_0 : boolean;
  signal ptr_deref_535_store_2_ack_0 : boolean;
  signal ptr_deref_540_load_0_ack_0 : boolean;
  signal ptr_deref_535_store_1_req_0 : boolean;
  signal ptr_deref_540_load_3_ack_0 : boolean;
  signal ptr_deref_535_gather_scatter_ack_0 : boolean;
  signal ptr_deref_540_load_3_req_0 : boolean;
  signal ptr_deref_535_store_2_ack_1 : boolean;
  signal ptr_deref_540_gather_scatter_ack_0 : boolean;
  signal ptr_deref_540_load_1_req_0 : boolean;
  signal ptr_deref_535_store_0_req_0 : boolean;
  signal array_obj_ref_545_base_resize_ack_0 : boolean;
  signal ptr_deref_540_load_1_req_1 : boolean;
  signal ptr_deref_535_store_3_ack_1 : boolean;
  signal ptr_deref_535_store_3_req_0 : boolean;
  signal ptr_deref_535_store_2_req_1 : boolean;
  signal ptr_deref_540_load_0_req_1 : boolean;
  signal ptr_deref_535_store_0_ack_0 : boolean;
  signal ptr_deref_540_gather_scatter_req_0 : boolean;
  signal ptr_deref_535_store_1_ack_1 : boolean;
  signal ptr_deref_540_load_2_ack_1 : boolean;
  signal ptr_deref_540_load_1_ack_0 : boolean;
  signal ptr_deref_540_load_2_ack_0 : boolean;
  signal ptr_deref_535_store_3_req_1 : boolean;
  signal ptr_deref_535_store_3_ack_0 : boolean;
  signal ptr_deref_535_store_1_req_1 : boolean;
  signal array_obj_ref_545_root_address_inst_req_0 : boolean;
  signal array_obj_ref_545_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_545_root_address_inst_req_1 : boolean;
  signal array_obj_ref_545_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_545_final_reg_req_0 : boolean;
  signal array_obj_ref_545_final_reg_ack_0 : boolean;
  signal ptr_deref_549_base_resize_req_0 : boolean;
  signal ptr_deref_549_base_resize_ack_0 : boolean;
  signal ptr_deref_549_root_address_inst_req_0 : boolean;
  signal ptr_deref_549_root_address_inst_ack_0 : boolean;
  signal ptr_deref_549_addr_0_req_0 : boolean;
  signal ptr_deref_549_addr_0_ack_0 : boolean;
  signal ptr_deref_549_addr_0_req_1 : boolean;
  signal ptr_deref_549_addr_0_ack_1 : boolean;
  signal ptr_deref_549_addr_1_req_0 : boolean;
  signal ptr_deref_549_addr_1_ack_0 : boolean;
  signal ptr_deref_549_addr_1_req_1 : boolean;
  signal ptr_deref_549_addr_1_ack_1 : boolean;
  signal ptr_deref_549_addr_2_req_0 : boolean;
  signal ptr_deref_549_addr_2_ack_0 : boolean;
  signal ptr_deref_549_addr_2_req_1 : boolean;
  signal ptr_deref_549_addr_2_ack_1 : boolean;
  signal ptr_deref_549_addr_3_req_0 : boolean;
  signal ptr_deref_549_addr_3_ack_0 : boolean;
  signal ptr_deref_549_addr_3_req_1 : boolean;
  signal ptr_deref_549_addr_3_ack_1 : boolean;
  signal ptr_deref_549_load_0_req_0 : boolean;
  signal ptr_deref_549_load_0_ack_0 : boolean;
  signal ptr_deref_549_load_1_req_0 : boolean;
  signal ptr_deref_549_load_1_ack_0 : boolean;
  signal ptr_deref_549_load_2_req_0 : boolean;
  signal ptr_deref_549_load_2_ack_0 : boolean;
  signal ptr_deref_549_load_3_req_0 : boolean;
  signal ptr_deref_549_load_3_ack_0 : boolean;
  signal ptr_deref_549_load_0_req_1 : boolean;
  signal ptr_deref_549_load_0_ack_1 : boolean;
  signal ptr_deref_549_load_1_req_1 : boolean;
  signal ptr_deref_549_load_1_ack_1 : boolean;
  signal ptr_deref_549_load_2_req_1 : boolean;
  signal ptr_deref_549_load_2_ack_1 : boolean;
  signal ptr_deref_549_load_3_req_1 : boolean;
  signal ptr_deref_549_load_3_ack_1 : boolean;
  signal ptr_deref_549_gather_scatter_req_0 : boolean;
  signal ptr_deref_549_gather_scatter_ack_0 : boolean;
  signal type_cast_558_inst_req_0 : boolean;
  signal type_cast_558_inst_ack_0 : boolean;
  signal simple_obj_ref_556_inst_req_0 : boolean;
  signal simple_obj_ref_556_inst_ack_0 : boolean;
  signal simple_obj_ref_565_inst_req_0 : boolean;
  signal simple_obj_ref_565_inst_ack_0 : boolean;
  signal ptr_deref_571_load_0_req_0 : boolean;
  signal ptr_deref_571_load_0_ack_0 : boolean;
  signal ptr_deref_571_load_1_req_0 : boolean;
  signal ptr_deref_571_load_1_ack_0 : boolean;
  signal ptr_deref_571_load_2_req_0 : boolean;
  signal ptr_deref_571_load_2_ack_0 : boolean;
  signal ptr_deref_571_load_3_req_0 : boolean;
  signal ptr_deref_571_load_3_ack_0 : boolean;
  signal ptr_deref_571_load_0_req_1 : boolean;
  signal ptr_deref_571_load_0_ack_1 : boolean;
  signal ptr_deref_571_load_1_req_1 : boolean;
  signal ptr_deref_571_load_1_ack_1 : boolean;
  signal ptr_deref_571_load_2_req_1 : boolean;
  signal ptr_deref_571_load_2_ack_1 : boolean;
  signal ptr_deref_571_load_3_req_1 : boolean;
  signal ptr_deref_571_load_3_ack_1 : boolean;
  signal ptr_deref_571_gather_scatter_req_0 : boolean;
  signal ptr_deref_571_gather_scatter_ack_0 : boolean;
  signal type_cast_575_inst_req_0 : boolean;
  signal type_cast_575_inst_ack_0 : boolean;
  signal type_cast_584_inst_req_0 : boolean;
  signal type_cast_584_inst_ack_0 : boolean;
  signal simple_obj_ref_582_inst_req_0 : boolean;
  signal simple_obj_ref_582_inst_ack_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  output_module_CP_3446: Block -- control-path 
    signal output_module_CP_3446_start: Boolean;
    signal Xentry_3447_symbol: Boolean;
    signal Xexit_3448_symbol: Boolean;
    signal branch_block_stmt_513_3449_symbol : Boolean;
    -- 
  begin -- 
    output_module_CP_3446_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_3447_symbol  <= output_module_CP_3446_start; -- transition $entry
    branch_block_stmt_513_3449: Block -- branch_block_stmt_513 
      signal branch_block_stmt_513_3449_start: Boolean;
      signal Xentry_3450_symbol: Boolean;
      signal Xexit_3451_symbol: Boolean;
      signal branch_block_stmt_513_x_xentry_x_xx_x3452_symbol : Boolean;
      signal branch_block_stmt_513_x_xexit_x_xx_x3453_symbol : Boolean;
      signal assign_stmt_518_x_xentry_x_xx_x3454_symbol : Boolean;
      signal assign_stmt_518_x_xexit_x_xx_x3455_symbol : Boolean;
      signal bb_0_bb_1_3456_symbol : Boolean;
      signal merge_stmt_520_x_xexit_x_xx_x3457_symbol : Boolean;
      signal assign_stmt_525_x_xentry_x_xx_x3458_symbol : Boolean;
      signal assign_stmt_525_x_xexit_x_xx_x3459_symbol : Boolean;
      signal assign_stmt_529_x_xentry_x_xx_x3460_symbol : Boolean;
      signal assign_stmt_529_x_xexit_x_xx_x3461_symbol : Boolean;
      signal assign_stmt_533_to_assign_stmt_555_x_xentry_x_xx_x3462_symbol : Boolean;
      signal assign_stmt_533_to_assign_stmt_555_x_xexit_x_xx_x3463_symbol : Boolean;
      signal assign_stmt_559_x_xentry_x_xx_x3464_symbol : Boolean;
      signal assign_stmt_559_x_xexit_x_xx_x3465_symbol : Boolean;
      signal assign_stmt_564_x_xentry_x_xx_x3466_symbol : Boolean;
      signal assign_stmt_564_x_xexit_x_xx_x3467_symbol : Boolean;
      signal assign_stmt_568_x_xentry_x_xx_x3468_symbol : Boolean;
      signal assign_stmt_568_x_xexit_x_xx_x3469_symbol : Boolean;
      signal assign_stmt_572_to_assign_stmt_581_x_xentry_x_xx_x3470_symbol : Boolean;
      signal assign_stmt_572_to_assign_stmt_581_x_xexit_x_xx_x3471_symbol : Boolean;
      signal assign_stmt_585_x_xentry_x_xx_x3472_symbol : Boolean;
      signal assign_stmt_585_x_xexit_x_xx_x3473_symbol : Boolean;
      signal bb_1_bb_1_3474_symbol : Boolean;
      signal assign_stmt_518_3475_symbol : Boolean;
      signal assign_stmt_525_3478_symbol : Boolean;
      signal assign_stmt_529_3481_symbol : Boolean;
      signal assign_stmt_533_to_assign_stmt_555_3499_symbol : Boolean;
      signal assign_stmt_559_3764_symbol : Boolean;
      signal assign_stmt_564_3783_symbol : Boolean;
      signal assign_stmt_568_3786_symbol : Boolean;
      signal assign_stmt_572_to_assign_stmt_581_3797_symbol : Boolean;
      signal assign_stmt_585_3871_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_3890_symbol : Boolean;
      signal bb_1_bb_1_PhiReq_3893_symbol : Boolean;
      signal merge_stmt_520_PhiReqMerge_3896_symbol : Boolean;
      signal merge_stmt_520_PhiAck_3897_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_513_3449_start <= Xentry_3447_symbol; -- control passed to block
      Xentry_3450_symbol  <= branch_block_stmt_513_3449_start; -- transition branch_block_stmt_513/$entry
      branch_block_stmt_513_x_xentry_x_xx_x3452_symbol  <=  Xentry_3450_symbol; -- place branch_block_stmt_513/branch_block_stmt_513__entry__ (optimized away) 
      branch_block_stmt_513_x_xexit_x_xx_x3453_symbol  <=   false ; -- place branch_block_stmt_513/branch_block_stmt_513__exit__ (optimized away) 
      assign_stmt_518_x_xentry_x_xx_x3454_symbol  <=  branch_block_stmt_513_x_xentry_x_xx_x3452_symbol; -- place branch_block_stmt_513/assign_stmt_518__entry__ (optimized away) 
      assign_stmt_518_x_xexit_x_xx_x3455_symbol  <=  assign_stmt_518_3475_symbol; -- place branch_block_stmt_513/assign_stmt_518__exit__ (optimized away) 
      bb_0_bb_1_3456_symbol  <=  assign_stmt_518_x_xexit_x_xx_x3455_symbol; -- place branch_block_stmt_513/bb_0_bb_1 (optimized away) 
      merge_stmt_520_x_xexit_x_xx_x3457_symbol  <=  merge_stmt_520_PhiAck_3897_symbol; -- place branch_block_stmt_513/merge_stmt_520__exit__ (optimized away) 
      assign_stmt_525_x_xentry_x_xx_x3458_symbol  <=  merge_stmt_520_x_xexit_x_xx_x3457_symbol; -- place branch_block_stmt_513/assign_stmt_525__entry__ (optimized away) 
      assign_stmt_525_x_xexit_x_xx_x3459_symbol  <=  assign_stmt_525_3478_symbol; -- place branch_block_stmt_513/assign_stmt_525__exit__ (optimized away) 
      assign_stmt_529_x_xentry_x_xx_x3460_symbol  <=  assign_stmt_525_x_xexit_x_xx_x3459_symbol; -- place branch_block_stmt_513/assign_stmt_529__entry__ (optimized away) 
      assign_stmt_529_x_xexit_x_xx_x3461_symbol  <=  assign_stmt_529_3481_symbol; -- place branch_block_stmt_513/assign_stmt_529__exit__ (optimized away) 
      assign_stmt_533_to_assign_stmt_555_x_xentry_x_xx_x3462_symbol  <=  assign_stmt_529_x_xexit_x_xx_x3461_symbol; -- place branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555__entry__ (optimized away) 
      assign_stmt_533_to_assign_stmt_555_x_xexit_x_xx_x3463_symbol  <=  assign_stmt_533_to_assign_stmt_555_3499_symbol; -- place branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555__exit__ (optimized away) 
      assign_stmt_559_x_xentry_x_xx_x3464_symbol  <=  assign_stmt_533_to_assign_stmt_555_x_xexit_x_xx_x3463_symbol; -- place branch_block_stmt_513/assign_stmt_559__entry__ (optimized away) 
      assign_stmt_559_x_xexit_x_xx_x3465_symbol  <=  assign_stmt_559_3764_symbol; -- place branch_block_stmt_513/assign_stmt_559__exit__ (optimized away) 
      assign_stmt_564_x_xentry_x_xx_x3466_symbol  <=  assign_stmt_559_x_xexit_x_xx_x3465_symbol; -- place branch_block_stmt_513/assign_stmt_564__entry__ (optimized away) 
      assign_stmt_564_x_xexit_x_xx_x3467_symbol  <=  assign_stmt_564_3783_symbol; -- place branch_block_stmt_513/assign_stmt_564__exit__ (optimized away) 
      assign_stmt_568_x_xentry_x_xx_x3468_symbol  <=  assign_stmt_564_x_xexit_x_xx_x3467_symbol; -- place branch_block_stmt_513/assign_stmt_568__entry__ (optimized away) 
      assign_stmt_568_x_xexit_x_xx_x3469_symbol  <=  assign_stmt_568_3786_symbol; -- place branch_block_stmt_513/assign_stmt_568__exit__ (optimized away) 
      assign_stmt_572_to_assign_stmt_581_x_xentry_x_xx_x3470_symbol  <=  assign_stmt_568_x_xexit_x_xx_x3469_symbol; -- place branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581__entry__ (optimized away) 
      assign_stmt_572_to_assign_stmt_581_x_xexit_x_xx_x3471_symbol  <=  assign_stmt_572_to_assign_stmt_581_3797_symbol; -- place branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581__exit__ (optimized away) 
      assign_stmt_585_x_xentry_x_xx_x3472_symbol  <=  assign_stmt_572_to_assign_stmt_581_x_xexit_x_xx_x3471_symbol; -- place branch_block_stmt_513/assign_stmt_585__entry__ (optimized away) 
      assign_stmt_585_x_xexit_x_xx_x3473_symbol  <=  assign_stmt_585_3871_symbol; -- place branch_block_stmt_513/assign_stmt_585__exit__ (optimized away) 
      bb_1_bb_1_3474_symbol  <=  assign_stmt_585_x_xexit_x_xx_x3473_symbol; -- place branch_block_stmt_513/bb_1_bb_1 (optimized away) 
      assign_stmt_518_3475: Block -- branch_block_stmt_513/assign_stmt_518 
        signal assign_stmt_518_3475_start: Boolean;
        signal Xentry_3476_symbol: Boolean;
        signal Xexit_3477_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_518_3475_start <= assign_stmt_518_x_xentry_x_xx_x3454_symbol; -- control passed to block
        Xentry_3476_symbol  <= assign_stmt_518_3475_start; -- transition branch_block_stmt_513/assign_stmt_518/$entry
        Xexit_3477_symbol <= Xentry_3476_symbol; -- transition branch_block_stmt_513/assign_stmt_518/$exit
        assign_stmt_518_3475_symbol <= Xexit_3477_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_518
      assign_stmt_525_3478: Block -- branch_block_stmt_513/assign_stmt_525 
        signal assign_stmt_525_3478_start: Boolean;
        signal Xentry_3479_symbol: Boolean;
        signal Xexit_3480_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_525_3478_start <= assign_stmt_525_x_xentry_x_xx_x3458_symbol; -- control passed to block
        Xentry_3479_symbol  <= assign_stmt_525_3478_start; -- transition branch_block_stmt_513/assign_stmt_525/$entry
        Xexit_3480_symbol <= Xentry_3479_symbol; -- transition branch_block_stmt_513/assign_stmt_525/$exit
        assign_stmt_525_3478_symbol <= Xexit_3480_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_525
      assign_stmt_529_3481: Block -- branch_block_stmt_513/assign_stmt_529 
        signal assign_stmt_529_3481_start: Boolean;
        signal Xentry_3482_symbol: Boolean;
        signal Xexit_3483_symbol: Boolean;
        signal assign_stmt_529_active_x_x3484_symbol : Boolean;
        signal assign_stmt_529_completed_x_x3485_symbol : Boolean;
        signal type_cast_528_active_x_x3486_symbol : Boolean;
        signal type_cast_528_trigger_x_x3487_symbol : Boolean;
        signal simple_obj_ref_527_trigger_x_x3488_symbol : Boolean;
        signal simple_obj_ref_527_complete_3489_symbol : Boolean;
        signal type_cast_528_complete_3494_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_529_3481_start <= assign_stmt_529_x_xentry_x_xx_x3460_symbol; -- control passed to block
        Xentry_3482_symbol  <= assign_stmt_529_3481_start; -- transition branch_block_stmt_513/assign_stmt_529/$entry
        assign_stmt_529_active_x_x3484_symbol <= type_cast_528_complete_3494_symbol; -- transition branch_block_stmt_513/assign_stmt_529/assign_stmt_529_active_
        assign_stmt_529_completed_x_x3485_symbol <= assign_stmt_529_active_x_x3484_symbol; -- transition branch_block_stmt_513/assign_stmt_529/assign_stmt_529_completed_
        type_cast_528_active_x_x3486_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_529/type_cast_528_active_ 
          signal type_cast_528_active_x_x3486_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_528_active_x_x3486_predecessors(0) <= type_cast_528_trigger_x_x3487_symbol;
          type_cast_528_active_x_x3486_predecessors(1) <= simple_obj_ref_527_complete_3489_symbol;
          type_cast_528_active_x_x3486_join: join -- 
            port map( -- 
              preds => type_cast_528_active_x_x3486_predecessors,
              symbol_out => type_cast_528_active_x_x3486_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_529/type_cast_528_active_
        type_cast_528_trigger_x_x3487_symbol <= Xentry_3482_symbol; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_trigger_
        simple_obj_ref_527_trigger_x_x3488_symbol <= Xentry_3482_symbol; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_trigger_
        simple_obj_ref_527_complete_3489: Block -- branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete 
          signal simple_obj_ref_527_complete_3489_start: Boolean;
          signal Xentry_3490_symbol: Boolean;
          signal Xexit_3491_symbol: Boolean;
          signal req_3492_symbol : Boolean;
          signal ack_3493_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_527_complete_3489_start <= simple_obj_ref_527_trigger_x_x3488_symbol; -- control passed to block
          Xentry_3490_symbol  <= simple_obj_ref_527_complete_3489_start; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/$entry
          req_3492_symbol <= Xentry_3490_symbol; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/req
          simple_obj_ref_527_inst_req_0 <= req_3492_symbol; -- link to DP
          ack_3493_symbol <= simple_obj_ref_527_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/ack
          Xexit_3491_symbol <= ack_3493_symbol; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/$exit
          simple_obj_ref_527_complete_3489_symbol <= Xexit_3491_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete
        type_cast_528_complete_3494: Block -- branch_block_stmt_513/assign_stmt_529/type_cast_528_complete 
          signal type_cast_528_complete_3494_start: Boolean;
          signal Xentry_3495_symbol: Boolean;
          signal Xexit_3496_symbol: Boolean;
          signal req_3497_symbol : Boolean;
          signal ack_3498_symbol : Boolean;
          -- 
        begin -- 
          type_cast_528_complete_3494_start <= type_cast_528_active_x_x3486_symbol; -- control passed to block
          Xentry_3495_symbol  <= type_cast_528_complete_3494_start; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/$entry
          req_3497_symbol <= Xentry_3495_symbol; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/req
          type_cast_528_inst_req_0 <= req_3497_symbol; -- link to DP
          ack_3498_symbol <= type_cast_528_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/ack
          Xexit_3496_symbol <= ack_3498_symbol; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/$exit
          type_cast_528_complete_3494_symbol <= Xexit_3496_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_529/type_cast_528_complete
        Xexit_3483_symbol <= assign_stmt_529_completed_x_x3485_symbol; -- transition branch_block_stmt_513/assign_stmt_529/$exit
        assign_stmt_529_3481_symbol <= Xexit_3483_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_529
      assign_stmt_533_to_assign_stmt_555_3499: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555 
        signal assign_stmt_533_to_assign_stmt_555_3499_start: Boolean;
        signal Xentry_3500_symbol: Boolean;
        signal Xexit_3501_symbol: Boolean;
        signal assign_stmt_533_active_x_x3502_symbol : Boolean;
        signal assign_stmt_533_completed_x_x3503_symbol : Boolean;
        signal type_cast_532_active_x_x3504_symbol : Boolean;
        signal type_cast_532_trigger_x_x3505_symbol : Boolean;
        signal simple_obj_ref_531_complete_3506_symbol : Boolean;
        signal type_cast_532_complete_3507_symbol : Boolean;
        signal assign_stmt_537_active_x_x3512_symbol : Boolean;
        signal assign_stmt_537_completed_x_x3513_symbol : Boolean;
        signal simple_obj_ref_536_complete_3514_symbol : Boolean;
        signal ptr_deref_535_trigger_x_x3515_symbol : Boolean;
        signal ptr_deref_535_active_x_x3516_symbol : Boolean;
        signal ptr_deref_535_base_address_calculated_3517_symbol : Boolean;
        signal ptr_deref_535_root_address_calculated_3518_symbol : Boolean;
        signal ptr_deref_535_word_address_calculated_3519_symbol : Boolean;
        signal ptr_deref_535_request_3520_symbol : Boolean;
        signal ptr_deref_535_complete_3548_symbol : Boolean;
        signal assign_stmt_541_active_x_x3574_symbol : Boolean;
        signal assign_stmt_541_completed_x_x3575_symbol : Boolean;
        signal ptr_deref_540_trigger_x_x3576_symbol : Boolean;
        signal ptr_deref_540_active_x_x3577_symbol : Boolean;
        signal ptr_deref_540_base_address_calculated_3578_symbol : Boolean;
        signal ptr_deref_540_root_address_calculated_3579_symbol : Boolean;
        signal ptr_deref_540_word_address_calculated_3580_symbol : Boolean;
        signal ptr_deref_540_request_3581_symbol : Boolean;
        signal ptr_deref_540_complete_3607_symbol : Boolean;
        signal assign_stmt_546_active_x_x3635_symbol : Boolean;
        signal assign_stmt_546_completed_x_x3636_symbol : Boolean;
        signal array_obj_ref_545_trigger_x_x3637_symbol : Boolean;
        signal array_obj_ref_545_active_x_x3638_symbol : Boolean;
        signal array_obj_ref_545_base_address_calculated_3639_symbol : Boolean;
        signal array_obj_ref_545_root_address_calculated_3640_symbol : Boolean;
        signal array_obj_ref_545_base_address_resized_3641_symbol : Boolean;
        signal array_obj_ref_545_base_addr_resize_3642_symbol : Boolean;
        signal array_obj_ref_545_base_plus_offset_trigger_3647_symbol : Boolean;
        signal array_obj_ref_545_base_plus_offset_3648_symbol : Boolean;
        signal array_obj_ref_545_complete_3655_symbol : Boolean;
        signal assign_stmt_550_active_x_x3660_symbol : Boolean;
        signal assign_stmt_550_completed_x_x3661_symbol : Boolean;
        signal ptr_deref_549_trigger_x_x3662_symbol : Boolean;
        signal ptr_deref_549_active_x_x3663_symbol : Boolean;
        signal ptr_deref_549_base_address_calculated_3664_symbol : Boolean;
        signal simple_obj_ref_548_complete_3665_symbol : Boolean;
        signal ptr_deref_549_root_address_calculated_3666_symbol : Boolean;
        signal ptr_deref_549_word_address_calculated_3667_symbol : Boolean;
        signal ptr_deref_549_base_address_resized_3668_symbol : Boolean;
        signal ptr_deref_549_base_addr_resize_3669_symbol : Boolean;
        signal ptr_deref_549_base_plus_offset_3674_symbol : Boolean;
        signal ptr_deref_549_word_addrgen_3679_symbol : Boolean;
        signal ptr_deref_549_request_3710_symbol : Boolean;
        signal ptr_deref_549_complete_3736_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_533_to_assign_stmt_555_3499_start <= assign_stmt_533_to_assign_stmt_555_x_xentry_x_xx_x3462_symbol; -- control passed to block
        Xentry_3500_symbol  <= assign_stmt_533_to_assign_stmt_555_3499_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/$entry
        assign_stmt_533_active_x_x3502_symbol <= type_cast_532_complete_3507_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_533_active_
        assign_stmt_533_completed_x_x3503_symbol <= assign_stmt_533_active_x_x3502_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_533_completed_
        type_cast_532_active_x_x3504_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_active_ 
          signal type_cast_532_active_x_x3504_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_532_active_x_x3504_predecessors(0) <= type_cast_532_trigger_x_x3505_symbol;
          type_cast_532_active_x_x3504_predecessors(1) <= simple_obj_ref_531_complete_3506_symbol;
          type_cast_532_active_x_x3504_join: join -- 
            port map( -- 
              preds => type_cast_532_active_x_x3504_predecessors,
              symbol_out => type_cast_532_active_x_x3504_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_active_
        type_cast_532_trigger_x_x3505_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_trigger_
        simple_obj_ref_531_complete_3506_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/simple_obj_ref_531_complete
        type_cast_532_complete_3507: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete 
          signal type_cast_532_complete_3507_start: Boolean;
          signal Xentry_3508_symbol: Boolean;
          signal Xexit_3509_symbol: Boolean;
          signal req_3510_symbol : Boolean;
          signal ack_3511_symbol : Boolean;
          -- 
        begin -- 
          type_cast_532_complete_3507_start <= type_cast_532_active_x_x3504_symbol; -- control passed to block
          Xentry_3508_symbol  <= type_cast_532_complete_3507_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/$entry
          req_3510_symbol <= Xentry_3508_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/req
          type_cast_532_inst_req_0 <= req_3510_symbol; -- link to DP
          ack_3511_symbol <= type_cast_532_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/ack
          Xexit_3509_symbol <= ack_3511_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/$exit
          type_cast_532_complete_3507_symbol <= Xexit_3509_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete
        assign_stmt_537_active_x_x3512_symbol <= simple_obj_ref_536_complete_3514_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_537_active_
        assign_stmt_537_completed_x_x3513_symbol <= ptr_deref_535_complete_3548_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_537_completed_
        simple_obj_ref_536_complete_3514_symbol <= assign_stmt_533_completed_x_x3503_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/simple_obj_ref_536_complete
        ptr_deref_535_trigger_x_x3515_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_trigger_ 
          signal ptr_deref_535_trigger_x_x3515_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_535_trigger_x_x3515_predecessors(0) <= ptr_deref_535_word_address_calculated_3519_symbol;
          ptr_deref_535_trigger_x_x3515_predecessors(1) <= assign_stmt_537_active_x_x3512_symbol;
          ptr_deref_535_trigger_x_x3515_join: join -- 
            port map( -- 
              preds => ptr_deref_535_trigger_x_x3515_predecessors,
              symbol_out => ptr_deref_535_trigger_x_x3515_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_trigger_
        ptr_deref_535_active_x_x3516_symbol <= ptr_deref_535_request_3520_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_active_
        ptr_deref_535_base_address_calculated_3517_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_base_address_calculated
        ptr_deref_535_root_address_calculated_3518_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_root_address_calculated
        ptr_deref_535_word_address_calculated_3519_symbol <= ptr_deref_535_root_address_calculated_3518_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_word_address_calculated
        ptr_deref_535_request_3520: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request 
          signal ptr_deref_535_request_3520_start: Boolean;
          signal Xentry_3521_symbol: Boolean;
          signal Xexit_3522_symbol: Boolean;
          signal split_req_3523_symbol : Boolean;
          signal split_ack_3524_symbol : Boolean;
          signal word_access_3525_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_535_request_3520_start <= ptr_deref_535_trigger_x_x3515_symbol; -- control passed to block
          Xentry_3521_symbol  <= ptr_deref_535_request_3520_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/$entry
          split_req_3523_symbol <= Xentry_3521_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/split_req
          ptr_deref_535_gather_scatter_req_0 <= split_req_3523_symbol; -- link to DP
          split_ack_3524_symbol <= ptr_deref_535_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/split_ack
          word_access_3525: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access 
            signal word_access_3525_start: Boolean;
            signal Xentry_3526_symbol: Boolean;
            signal Xexit_3527_symbol: Boolean;
            signal word_access_0_3528_symbol : Boolean;
            signal word_access_1_3533_symbol : Boolean;
            signal word_access_2_3538_symbol : Boolean;
            signal word_access_3_3543_symbol : Boolean;
            -- 
          begin -- 
            word_access_3525_start <= split_ack_3524_symbol; -- control passed to block
            Xentry_3526_symbol  <= word_access_3525_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/$entry
            word_access_0_3528: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0 
              signal word_access_0_3528_start: Boolean;
              signal Xentry_3529_symbol: Boolean;
              signal Xexit_3530_symbol: Boolean;
              signal rr_3531_symbol : Boolean;
              signal ra_3532_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3528_start <= Xentry_3526_symbol; -- control passed to block
              Xentry_3529_symbol  <= word_access_0_3528_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/$entry
              rr_3531_symbol <= Xentry_3529_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/rr
              ptr_deref_535_store_0_req_0 <= rr_3531_symbol; -- link to DP
              ra_3532_symbol <= ptr_deref_535_store_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/ra
              Xexit_3530_symbol <= ra_3532_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/$exit
              word_access_0_3528_symbol <= Xexit_3530_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0
            word_access_1_3533: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_1 
              signal word_access_1_3533_start: Boolean;
              signal Xentry_3534_symbol: Boolean;
              signal Xexit_3535_symbol: Boolean;
              signal rr_3536_symbol : Boolean;
              signal ra_3537_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3533_start <= Xentry_3526_symbol; -- control passed to block
              Xentry_3534_symbol  <= word_access_1_3533_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_1/$entry
              rr_3536_symbol <= Xentry_3534_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_1/rr
              ptr_deref_535_store_1_req_0 <= rr_3536_symbol; -- link to DP
              ra_3537_symbol <= ptr_deref_535_store_1_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_1/ra
              Xexit_3535_symbol <= ra_3537_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_1/$exit
              word_access_1_3533_symbol <= Xexit_3535_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_1
            word_access_2_3538: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_2 
              signal word_access_2_3538_start: Boolean;
              signal Xentry_3539_symbol: Boolean;
              signal Xexit_3540_symbol: Boolean;
              signal rr_3541_symbol : Boolean;
              signal ra_3542_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3538_start <= Xentry_3526_symbol; -- control passed to block
              Xentry_3539_symbol  <= word_access_2_3538_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_2/$entry
              rr_3541_symbol <= Xentry_3539_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_2/rr
              ptr_deref_535_store_2_req_0 <= rr_3541_symbol; -- link to DP
              ra_3542_symbol <= ptr_deref_535_store_2_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_2/ra
              Xexit_3540_symbol <= ra_3542_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_2/$exit
              word_access_2_3538_symbol <= Xexit_3540_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_2
            word_access_3_3543: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_3 
              signal word_access_3_3543_start: Boolean;
              signal Xentry_3544_symbol: Boolean;
              signal Xexit_3545_symbol: Boolean;
              signal rr_3546_symbol : Boolean;
              signal ra_3547_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3543_start <= Xentry_3526_symbol; -- control passed to block
              Xentry_3544_symbol  <= word_access_3_3543_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_3/$entry
              rr_3546_symbol <= Xentry_3544_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_3/rr
              ptr_deref_535_store_3_req_0 <= rr_3546_symbol; -- link to DP
              ra_3547_symbol <= ptr_deref_535_store_3_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_3/ra
              Xexit_3545_symbol <= ra_3547_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_3/$exit
              word_access_3_3543_symbol <= Xexit_3545_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_3
            Xexit_3527_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/$exit 
              signal Xexit_3527_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3527_predecessors(0) <= word_access_0_3528_symbol;
              Xexit_3527_predecessors(1) <= word_access_1_3533_symbol;
              Xexit_3527_predecessors(2) <= word_access_2_3538_symbol;
              Xexit_3527_predecessors(3) <= word_access_3_3543_symbol;
              Xexit_3527_join: join -- 
                port map( -- 
                  preds => Xexit_3527_predecessors,
                  symbol_out => Xexit_3527_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/$exit
            word_access_3525_symbol <= Xexit_3527_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access
          Xexit_3522_symbol <= word_access_3525_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/$exit
          ptr_deref_535_request_3520_symbol <= Xexit_3522_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request
        ptr_deref_535_complete_3548: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete 
          signal ptr_deref_535_complete_3548_start: Boolean;
          signal Xentry_3549_symbol: Boolean;
          signal Xexit_3550_symbol: Boolean;
          signal word_access_3551_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_535_complete_3548_start <= ptr_deref_535_active_x_x3516_symbol; -- control passed to block
          Xentry_3549_symbol  <= ptr_deref_535_complete_3548_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/$entry
          word_access_3551: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access 
            signal word_access_3551_start: Boolean;
            signal Xentry_3552_symbol: Boolean;
            signal Xexit_3553_symbol: Boolean;
            signal word_access_0_3554_symbol : Boolean;
            signal word_access_1_3559_symbol : Boolean;
            signal word_access_2_3564_symbol : Boolean;
            signal word_access_3_3569_symbol : Boolean;
            -- 
          begin -- 
            word_access_3551_start <= Xentry_3549_symbol; -- control passed to block
            Xentry_3552_symbol  <= word_access_3551_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/$entry
            word_access_0_3554: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0 
              signal word_access_0_3554_start: Boolean;
              signal Xentry_3555_symbol: Boolean;
              signal Xexit_3556_symbol: Boolean;
              signal cr_3557_symbol : Boolean;
              signal ca_3558_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3554_start <= Xentry_3552_symbol; -- control passed to block
              Xentry_3555_symbol  <= word_access_0_3554_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/$entry
              cr_3557_symbol <= Xentry_3555_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/cr
              ptr_deref_535_store_0_req_1 <= cr_3557_symbol; -- link to DP
              ca_3558_symbol <= ptr_deref_535_store_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/ca
              Xexit_3556_symbol <= ca_3558_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/$exit
              word_access_0_3554_symbol <= Xexit_3556_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0
            word_access_1_3559: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_1 
              signal word_access_1_3559_start: Boolean;
              signal Xentry_3560_symbol: Boolean;
              signal Xexit_3561_symbol: Boolean;
              signal cr_3562_symbol : Boolean;
              signal ca_3563_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3559_start <= Xentry_3552_symbol; -- control passed to block
              Xentry_3560_symbol  <= word_access_1_3559_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_1/$entry
              cr_3562_symbol <= Xentry_3560_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_1/cr
              ptr_deref_535_store_1_req_1 <= cr_3562_symbol; -- link to DP
              ca_3563_symbol <= ptr_deref_535_store_1_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_1/ca
              Xexit_3561_symbol <= ca_3563_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_1/$exit
              word_access_1_3559_symbol <= Xexit_3561_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_1
            word_access_2_3564: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_2 
              signal word_access_2_3564_start: Boolean;
              signal Xentry_3565_symbol: Boolean;
              signal Xexit_3566_symbol: Boolean;
              signal cr_3567_symbol : Boolean;
              signal ca_3568_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3564_start <= Xentry_3552_symbol; -- control passed to block
              Xentry_3565_symbol  <= word_access_2_3564_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_2/$entry
              cr_3567_symbol <= Xentry_3565_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_2/cr
              ptr_deref_535_store_2_req_1 <= cr_3567_symbol; -- link to DP
              ca_3568_symbol <= ptr_deref_535_store_2_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_2/ca
              Xexit_3566_symbol <= ca_3568_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_2/$exit
              word_access_2_3564_symbol <= Xexit_3566_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_2
            word_access_3_3569: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_3 
              signal word_access_3_3569_start: Boolean;
              signal Xentry_3570_symbol: Boolean;
              signal Xexit_3571_symbol: Boolean;
              signal cr_3572_symbol : Boolean;
              signal ca_3573_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3569_start <= Xentry_3552_symbol; -- control passed to block
              Xentry_3570_symbol  <= word_access_3_3569_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_3/$entry
              cr_3572_symbol <= Xentry_3570_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_3/cr
              ptr_deref_535_store_3_req_1 <= cr_3572_symbol; -- link to DP
              ca_3573_symbol <= ptr_deref_535_store_3_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_3/ca
              Xexit_3571_symbol <= ca_3573_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_3/$exit
              word_access_3_3569_symbol <= Xexit_3571_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_3
            Xexit_3553_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/$exit 
              signal Xexit_3553_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3553_predecessors(0) <= word_access_0_3554_symbol;
              Xexit_3553_predecessors(1) <= word_access_1_3559_symbol;
              Xexit_3553_predecessors(2) <= word_access_2_3564_symbol;
              Xexit_3553_predecessors(3) <= word_access_3_3569_symbol;
              Xexit_3553_join: join -- 
                port map( -- 
                  preds => Xexit_3553_predecessors,
                  symbol_out => Xexit_3553_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/$exit
            word_access_3551_symbol <= Xexit_3553_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access
          Xexit_3550_symbol <= word_access_3551_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/$exit
          ptr_deref_535_complete_3548_symbol <= Xexit_3550_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete
        assign_stmt_541_active_x_x3574_symbol <= ptr_deref_540_complete_3607_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_541_active_
        assign_stmt_541_completed_x_x3575_symbol <= assign_stmt_541_active_x_x3574_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_541_completed_
        ptr_deref_540_trigger_x_x3576_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_trigger_ 
          signal ptr_deref_540_trigger_x_x3576_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_540_trigger_x_x3576_predecessors(0) <= ptr_deref_540_word_address_calculated_3580_symbol;
          ptr_deref_540_trigger_x_x3576_predecessors(1) <= ptr_deref_535_active_x_x3516_symbol;
          ptr_deref_540_trigger_x_x3576_join: join -- 
            port map( -- 
              preds => ptr_deref_540_trigger_x_x3576_predecessors,
              symbol_out => ptr_deref_540_trigger_x_x3576_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_trigger_
        ptr_deref_540_active_x_x3577_symbol <= ptr_deref_540_request_3581_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_active_
        ptr_deref_540_base_address_calculated_3578_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_base_address_calculated
        ptr_deref_540_root_address_calculated_3579_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_root_address_calculated
        ptr_deref_540_word_address_calculated_3580_symbol <= ptr_deref_540_root_address_calculated_3579_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_word_address_calculated
        ptr_deref_540_request_3581: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request 
          signal ptr_deref_540_request_3581_start: Boolean;
          signal Xentry_3582_symbol: Boolean;
          signal Xexit_3583_symbol: Boolean;
          signal word_access_3584_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_540_request_3581_start <= ptr_deref_540_trigger_x_x3576_symbol; -- control passed to block
          Xentry_3582_symbol  <= ptr_deref_540_request_3581_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/$entry
          word_access_3584: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access 
            signal word_access_3584_start: Boolean;
            signal Xentry_3585_symbol: Boolean;
            signal Xexit_3586_symbol: Boolean;
            signal word_access_0_3587_symbol : Boolean;
            signal word_access_1_3592_symbol : Boolean;
            signal word_access_2_3597_symbol : Boolean;
            signal word_access_3_3602_symbol : Boolean;
            -- 
          begin -- 
            word_access_3584_start <= Xentry_3582_symbol; -- control passed to block
            Xentry_3585_symbol  <= word_access_3584_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/$entry
            word_access_0_3587: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0 
              signal word_access_0_3587_start: Boolean;
              signal Xentry_3588_symbol: Boolean;
              signal Xexit_3589_symbol: Boolean;
              signal rr_3590_symbol : Boolean;
              signal ra_3591_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3587_start <= Xentry_3585_symbol; -- control passed to block
              Xentry_3588_symbol  <= word_access_0_3587_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/$entry
              rr_3590_symbol <= Xentry_3588_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/rr
              ptr_deref_540_load_0_req_0 <= rr_3590_symbol; -- link to DP
              ra_3591_symbol <= ptr_deref_540_load_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/ra
              Xexit_3589_symbol <= ra_3591_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/$exit
              word_access_0_3587_symbol <= Xexit_3589_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0
            word_access_1_3592: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_1 
              signal word_access_1_3592_start: Boolean;
              signal Xentry_3593_symbol: Boolean;
              signal Xexit_3594_symbol: Boolean;
              signal rr_3595_symbol : Boolean;
              signal ra_3596_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3592_start <= Xentry_3585_symbol; -- control passed to block
              Xentry_3593_symbol  <= word_access_1_3592_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_1/$entry
              rr_3595_symbol <= Xentry_3593_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_1/rr
              ptr_deref_540_load_1_req_0 <= rr_3595_symbol; -- link to DP
              ra_3596_symbol <= ptr_deref_540_load_1_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_1/ra
              Xexit_3594_symbol <= ra_3596_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_1/$exit
              word_access_1_3592_symbol <= Xexit_3594_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_1
            word_access_2_3597: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_2 
              signal word_access_2_3597_start: Boolean;
              signal Xentry_3598_symbol: Boolean;
              signal Xexit_3599_symbol: Boolean;
              signal rr_3600_symbol : Boolean;
              signal ra_3601_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3597_start <= Xentry_3585_symbol; -- control passed to block
              Xentry_3598_symbol  <= word_access_2_3597_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_2/$entry
              rr_3600_symbol <= Xentry_3598_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_2/rr
              ptr_deref_540_load_2_req_0 <= rr_3600_symbol; -- link to DP
              ra_3601_symbol <= ptr_deref_540_load_2_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_2/ra
              Xexit_3599_symbol <= ra_3601_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_2/$exit
              word_access_2_3597_symbol <= Xexit_3599_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_2
            word_access_3_3602: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_3 
              signal word_access_3_3602_start: Boolean;
              signal Xentry_3603_symbol: Boolean;
              signal Xexit_3604_symbol: Boolean;
              signal rr_3605_symbol : Boolean;
              signal ra_3606_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3602_start <= Xentry_3585_symbol; -- control passed to block
              Xentry_3603_symbol  <= word_access_3_3602_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_3/$entry
              rr_3605_symbol <= Xentry_3603_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_3/rr
              ptr_deref_540_load_3_req_0 <= rr_3605_symbol; -- link to DP
              ra_3606_symbol <= ptr_deref_540_load_3_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_3/ra
              Xexit_3604_symbol <= ra_3606_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_3/$exit
              word_access_3_3602_symbol <= Xexit_3604_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_3
            Xexit_3586_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/$exit 
              signal Xexit_3586_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3586_predecessors(0) <= word_access_0_3587_symbol;
              Xexit_3586_predecessors(1) <= word_access_1_3592_symbol;
              Xexit_3586_predecessors(2) <= word_access_2_3597_symbol;
              Xexit_3586_predecessors(3) <= word_access_3_3602_symbol;
              Xexit_3586_join: join -- 
                port map( -- 
                  preds => Xexit_3586_predecessors,
                  symbol_out => Xexit_3586_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/$exit
            word_access_3584_symbol <= Xexit_3586_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access
          Xexit_3583_symbol <= word_access_3584_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/$exit
          ptr_deref_540_request_3581_symbol <= Xexit_3583_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request
        ptr_deref_540_complete_3607: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete 
          signal ptr_deref_540_complete_3607_start: Boolean;
          signal Xentry_3608_symbol: Boolean;
          signal Xexit_3609_symbol: Boolean;
          signal word_access_3610_symbol : Boolean;
          signal merge_req_3633_symbol : Boolean;
          signal merge_ack_3634_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_540_complete_3607_start <= ptr_deref_540_active_x_x3577_symbol; -- control passed to block
          Xentry_3608_symbol  <= ptr_deref_540_complete_3607_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/$entry
          word_access_3610: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access 
            signal word_access_3610_start: Boolean;
            signal Xentry_3611_symbol: Boolean;
            signal Xexit_3612_symbol: Boolean;
            signal word_access_0_3613_symbol : Boolean;
            signal word_access_1_3618_symbol : Boolean;
            signal word_access_2_3623_symbol : Boolean;
            signal word_access_3_3628_symbol : Boolean;
            -- 
          begin -- 
            word_access_3610_start <= Xentry_3608_symbol; -- control passed to block
            Xentry_3611_symbol  <= word_access_3610_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/$entry
            word_access_0_3613: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0 
              signal word_access_0_3613_start: Boolean;
              signal Xentry_3614_symbol: Boolean;
              signal Xexit_3615_symbol: Boolean;
              signal cr_3616_symbol : Boolean;
              signal ca_3617_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3613_start <= Xentry_3611_symbol; -- control passed to block
              Xentry_3614_symbol  <= word_access_0_3613_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/$entry
              cr_3616_symbol <= Xentry_3614_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/cr
              ptr_deref_540_load_0_req_1 <= cr_3616_symbol; -- link to DP
              ca_3617_symbol <= ptr_deref_540_load_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/ca
              Xexit_3615_symbol <= ca_3617_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/$exit
              word_access_0_3613_symbol <= Xexit_3615_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0
            word_access_1_3618: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_1 
              signal word_access_1_3618_start: Boolean;
              signal Xentry_3619_symbol: Boolean;
              signal Xexit_3620_symbol: Boolean;
              signal cr_3621_symbol : Boolean;
              signal ca_3622_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3618_start <= Xentry_3611_symbol; -- control passed to block
              Xentry_3619_symbol  <= word_access_1_3618_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_1/$entry
              cr_3621_symbol <= Xentry_3619_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_1/cr
              ptr_deref_540_load_1_req_1 <= cr_3621_symbol; -- link to DP
              ca_3622_symbol <= ptr_deref_540_load_1_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_1/ca
              Xexit_3620_symbol <= ca_3622_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_1/$exit
              word_access_1_3618_symbol <= Xexit_3620_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_1
            word_access_2_3623: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_2 
              signal word_access_2_3623_start: Boolean;
              signal Xentry_3624_symbol: Boolean;
              signal Xexit_3625_symbol: Boolean;
              signal cr_3626_symbol : Boolean;
              signal ca_3627_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3623_start <= Xentry_3611_symbol; -- control passed to block
              Xentry_3624_symbol  <= word_access_2_3623_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_2/$entry
              cr_3626_symbol <= Xentry_3624_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_2/cr
              ptr_deref_540_load_2_req_1 <= cr_3626_symbol; -- link to DP
              ca_3627_symbol <= ptr_deref_540_load_2_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_2/ca
              Xexit_3625_symbol <= ca_3627_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_2/$exit
              word_access_2_3623_symbol <= Xexit_3625_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_2
            word_access_3_3628: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_3 
              signal word_access_3_3628_start: Boolean;
              signal Xentry_3629_symbol: Boolean;
              signal Xexit_3630_symbol: Boolean;
              signal cr_3631_symbol : Boolean;
              signal ca_3632_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3628_start <= Xentry_3611_symbol; -- control passed to block
              Xentry_3629_symbol  <= word_access_3_3628_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_3/$entry
              cr_3631_symbol <= Xentry_3629_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_3/cr
              ptr_deref_540_load_3_req_1 <= cr_3631_symbol; -- link to DP
              ca_3632_symbol <= ptr_deref_540_load_3_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_3/ca
              Xexit_3630_symbol <= ca_3632_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_3/$exit
              word_access_3_3628_symbol <= Xexit_3630_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_3
            Xexit_3612_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/$exit 
              signal Xexit_3612_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3612_predecessors(0) <= word_access_0_3613_symbol;
              Xexit_3612_predecessors(1) <= word_access_1_3618_symbol;
              Xexit_3612_predecessors(2) <= word_access_2_3623_symbol;
              Xexit_3612_predecessors(3) <= word_access_3_3628_symbol;
              Xexit_3612_join: join -- 
                port map( -- 
                  preds => Xexit_3612_predecessors,
                  symbol_out => Xexit_3612_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/$exit
            word_access_3610_symbol <= Xexit_3612_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access
          merge_req_3633_symbol <= word_access_3610_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/merge_req
          ptr_deref_540_gather_scatter_req_0 <= merge_req_3633_symbol; -- link to DP
          merge_ack_3634_symbol <= ptr_deref_540_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/merge_ack
          Xexit_3609_symbol <= merge_ack_3634_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/$exit
          ptr_deref_540_complete_3607_symbol <= Xexit_3609_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete
        assign_stmt_546_active_x_x3635_symbol <= array_obj_ref_545_complete_3655_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_546_active_
        assign_stmt_546_completed_x_x3636_symbol <= assign_stmt_546_active_x_x3635_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_546_completed_
        array_obj_ref_545_trigger_x_x3637_symbol <= Xentry_3500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_trigger_
        array_obj_ref_545_active_x_x3638_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_active_ 
          signal array_obj_ref_545_active_x_x3638_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_545_active_x_x3638_predecessors(0) <= array_obj_ref_545_trigger_x_x3637_symbol;
          array_obj_ref_545_active_x_x3638_predecessors(1) <= array_obj_ref_545_root_address_calculated_3640_symbol;
          array_obj_ref_545_active_x_x3638_join: join -- 
            port map( -- 
              preds => array_obj_ref_545_active_x_x3638_predecessors,
              symbol_out => array_obj_ref_545_active_x_x3638_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_active_
        array_obj_ref_545_base_address_calculated_3639_symbol <= assign_stmt_541_completed_x_x3575_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_address_calculated
        array_obj_ref_545_root_address_calculated_3640_symbol <= array_obj_ref_545_base_plus_offset_3648_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_root_address_calculated
        array_obj_ref_545_base_address_resized_3641_symbol <= array_obj_ref_545_base_addr_resize_3642_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_address_resized
        array_obj_ref_545_base_addr_resize_3642: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize 
          signal array_obj_ref_545_base_addr_resize_3642_start: Boolean;
          signal Xentry_3643_symbol: Boolean;
          signal Xexit_3644_symbol: Boolean;
          signal base_resize_req_3645_symbol : Boolean;
          signal base_resize_ack_3646_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_545_base_addr_resize_3642_start <= array_obj_ref_545_base_address_calculated_3639_symbol; -- control passed to block
          Xentry_3643_symbol  <= array_obj_ref_545_base_addr_resize_3642_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/$entry
          base_resize_req_3645_symbol <= Xentry_3643_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/base_resize_req
          array_obj_ref_545_base_resize_req_0 <= base_resize_req_3645_symbol; -- link to DP
          base_resize_ack_3646_symbol <= array_obj_ref_545_base_resize_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/base_resize_ack
          Xexit_3644_symbol <= base_resize_ack_3646_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/$exit
          array_obj_ref_545_base_addr_resize_3642_symbol <= Xexit_3644_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize
        array_obj_ref_545_base_plus_offset_trigger_3647_symbol <= array_obj_ref_545_base_address_resized_3641_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset_trigger
        array_obj_ref_545_base_plus_offset_3648: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset 
          signal array_obj_ref_545_base_plus_offset_3648_start: Boolean;
          signal Xentry_3649_symbol: Boolean;
          signal Xexit_3650_symbol: Boolean;
          signal plus_base_rr_3651_symbol : Boolean;
          signal plus_base_ra_3652_symbol : Boolean;
          signal plus_base_cr_3653_symbol : Boolean;
          signal plus_base_ca_3654_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_545_base_plus_offset_3648_start <= array_obj_ref_545_base_plus_offset_trigger_3647_symbol; -- control passed to block
          Xentry_3649_symbol  <= array_obj_ref_545_base_plus_offset_3648_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/$entry
          plus_base_rr_3651_symbol <= Xentry_3649_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_rr
          array_obj_ref_545_root_address_inst_req_0 <= plus_base_rr_3651_symbol; -- link to DP
          plus_base_ra_3652_symbol <= array_obj_ref_545_root_address_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_ra
          plus_base_cr_3653_symbol <= plus_base_ra_3652_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_cr
          array_obj_ref_545_root_address_inst_req_1 <= plus_base_cr_3653_symbol; -- link to DP
          plus_base_ca_3654_symbol <= array_obj_ref_545_root_address_inst_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_ca
          Xexit_3650_symbol <= plus_base_ca_3654_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/$exit
          array_obj_ref_545_base_plus_offset_3648_symbol <= Xexit_3650_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset
        array_obj_ref_545_complete_3655: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete 
          signal array_obj_ref_545_complete_3655_start: Boolean;
          signal Xentry_3656_symbol: Boolean;
          signal Xexit_3657_symbol: Boolean;
          signal final_reg_req_3658_symbol : Boolean;
          signal final_reg_ack_3659_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_545_complete_3655_start <= array_obj_ref_545_active_x_x3638_symbol; -- control passed to block
          Xentry_3656_symbol  <= array_obj_ref_545_complete_3655_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/$entry
          final_reg_req_3658_symbol <= Xentry_3656_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/final_reg_req
          array_obj_ref_545_final_reg_req_0 <= final_reg_req_3658_symbol; -- link to DP
          final_reg_ack_3659_symbol <= array_obj_ref_545_final_reg_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/final_reg_ack
          Xexit_3657_symbol <= final_reg_ack_3659_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/$exit
          array_obj_ref_545_complete_3655_symbol <= Xexit_3657_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete
        assign_stmt_550_active_x_x3660_symbol <= ptr_deref_549_complete_3736_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_550_active_
        assign_stmt_550_completed_x_x3661_symbol <= assign_stmt_550_active_x_x3660_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_550_completed_
        ptr_deref_549_trigger_x_x3662_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_trigger_ 
          signal ptr_deref_549_trigger_x_x3662_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          ptr_deref_549_trigger_x_x3662_predecessors(0) <= ptr_deref_549_word_address_calculated_3667_symbol;
          ptr_deref_549_trigger_x_x3662_predecessors(1) <= ptr_deref_549_base_address_calculated_3664_symbol;
          ptr_deref_549_trigger_x_x3662_predecessors(2) <= ptr_deref_535_active_x_x3516_symbol;
          ptr_deref_549_trigger_x_x3662_join: join -- 
            port map( -- 
              preds => ptr_deref_549_trigger_x_x3662_predecessors,
              symbol_out => ptr_deref_549_trigger_x_x3662_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_trigger_
        ptr_deref_549_active_x_x3663_symbol <= ptr_deref_549_request_3710_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_active_
        ptr_deref_549_base_address_calculated_3664_symbol <= simple_obj_ref_548_complete_3665_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_address_calculated
        simple_obj_ref_548_complete_3665_symbol <= assign_stmt_546_completed_x_x3636_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/simple_obj_ref_548_complete
        ptr_deref_549_root_address_calculated_3666_symbol <= ptr_deref_549_base_plus_offset_3674_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_root_address_calculated
        ptr_deref_549_word_address_calculated_3667_symbol <= ptr_deref_549_word_addrgen_3679_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_address_calculated
        ptr_deref_549_base_address_resized_3668_symbol <= ptr_deref_549_base_addr_resize_3669_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_address_resized
        ptr_deref_549_base_addr_resize_3669: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize 
          signal ptr_deref_549_base_addr_resize_3669_start: Boolean;
          signal Xentry_3670_symbol: Boolean;
          signal Xexit_3671_symbol: Boolean;
          signal base_resize_req_3672_symbol : Boolean;
          signal base_resize_ack_3673_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_base_addr_resize_3669_start <= ptr_deref_549_base_address_calculated_3664_symbol; -- control passed to block
          Xentry_3670_symbol  <= ptr_deref_549_base_addr_resize_3669_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/$entry
          base_resize_req_3672_symbol <= Xentry_3670_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/base_resize_req
          ptr_deref_549_base_resize_req_0 <= base_resize_req_3672_symbol; -- link to DP
          base_resize_ack_3673_symbol <= ptr_deref_549_base_resize_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/base_resize_ack
          Xexit_3671_symbol <= base_resize_ack_3673_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/$exit
          ptr_deref_549_base_addr_resize_3669_symbol <= Xexit_3671_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize
        ptr_deref_549_base_plus_offset_3674: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset 
          signal ptr_deref_549_base_plus_offset_3674_start: Boolean;
          signal Xentry_3675_symbol: Boolean;
          signal Xexit_3676_symbol: Boolean;
          signal sum_rename_req_3677_symbol : Boolean;
          signal sum_rename_ack_3678_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_base_plus_offset_3674_start <= ptr_deref_549_base_address_resized_3668_symbol; -- control passed to block
          Xentry_3675_symbol  <= ptr_deref_549_base_plus_offset_3674_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/$entry
          sum_rename_req_3677_symbol <= Xentry_3675_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/sum_rename_req
          ptr_deref_549_root_address_inst_req_0 <= sum_rename_req_3677_symbol; -- link to DP
          sum_rename_ack_3678_symbol <= ptr_deref_549_root_address_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/sum_rename_ack
          Xexit_3676_symbol <= sum_rename_ack_3678_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/$exit
          ptr_deref_549_base_plus_offset_3674_symbol <= Xexit_3676_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset
        ptr_deref_549_word_addrgen_3679: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen 
          signal ptr_deref_549_word_addrgen_3679_start: Boolean;
          signal Xentry_3680_symbol: Boolean;
          signal Xexit_3681_symbol: Boolean;
          signal word_0_3682_symbol : Boolean;
          signal word_1_3689_symbol : Boolean;
          signal word_2_3696_symbol : Boolean;
          signal word_3_3703_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_word_addrgen_3679_start <= ptr_deref_549_root_address_calculated_3666_symbol; -- control passed to block
          Xentry_3680_symbol  <= ptr_deref_549_word_addrgen_3679_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/$entry
          word_0_3682: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0 
            signal word_0_3682_start: Boolean;
            signal Xentry_3683_symbol: Boolean;
            signal Xexit_3684_symbol: Boolean;
            signal rr_3685_symbol : Boolean;
            signal ra_3686_symbol : Boolean;
            signal cr_3687_symbol : Boolean;
            signal ca_3688_symbol : Boolean;
            -- 
          begin -- 
            word_0_3682_start <= Xentry_3680_symbol; -- control passed to block
            Xentry_3683_symbol  <= word_0_3682_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0/$entry
            rr_3685_symbol <= Xentry_3683_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0/rr
            ptr_deref_549_addr_0_req_0 <= rr_3685_symbol; -- link to DP
            ra_3686_symbol <= ptr_deref_549_addr_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0/ra
            cr_3687_symbol <= ra_3686_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0/cr
            ptr_deref_549_addr_0_req_1 <= cr_3687_symbol; -- link to DP
            ca_3688_symbol <= ptr_deref_549_addr_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0/ca
            Xexit_3684_symbol <= ca_3688_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0/$exit
            word_0_3682_symbol <= Xexit_3684_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_0
          word_1_3689: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1 
            signal word_1_3689_start: Boolean;
            signal Xentry_3690_symbol: Boolean;
            signal Xexit_3691_symbol: Boolean;
            signal rr_3692_symbol : Boolean;
            signal ra_3693_symbol : Boolean;
            signal cr_3694_symbol : Boolean;
            signal ca_3695_symbol : Boolean;
            -- 
          begin -- 
            word_1_3689_start <= Xentry_3680_symbol; -- control passed to block
            Xentry_3690_symbol  <= word_1_3689_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1/$entry
            rr_3692_symbol <= Xentry_3690_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1/rr
            ptr_deref_549_addr_1_req_0 <= rr_3692_symbol; -- link to DP
            ra_3693_symbol <= ptr_deref_549_addr_1_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1/ra
            cr_3694_symbol <= ra_3693_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1/cr
            ptr_deref_549_addr_1_req_1 <= cr_3694_symbol; -- link to DP
            ca_3695_symbol <= ptr_deref_549_addr_1_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1/ca
            Xexit_3691_symbol <= ca_3695_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1/$exit
            word_1_3689_symbol <= Xexit_3691_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_1
          word_2_3696: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2 
            signal word_2_3696_start: Boolean;
            signal Xentry_3697_symbol: Boolean;
            signal Xexit_3698_symbol: Boolean;
            signal rr_3699_symbol : Boolean;
            signal ra_3700_symbol : Boolean;
            signal cr_3701_symbol : Boolean;
            signal ca_3702_symbol : Boolean;
            -- 
          begin -- 
            word_2_3696_start <= Xentry_3680_symbol; -- control passed to block
            Xentry_3697_symbol  <= word_2_3696_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2/$entry
            rr_3699_symbol <= Xentry_3697_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2/rr
            ptr_deref_549_addr_2_req_0 <= rr_3699_symbol; -- link to DP
            ra_3700_symbol <= ptr_deref_549_addr_2_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2/ra
            cr_3701_symbol <= ra_3700_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2/cr
            ptr_deref_549_addr_2_req_1 <= cr_3701_symbol; -- link to DP
            ca_3702_symbol <= ptr_deref_549_addr_2_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2/ca
            Xexit_3698_symbol <= ca_3702_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2/$exit
            word_2_3696_symbol <= Xexit_3698_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_2
          word_3_3703: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3 
            signal word_3_3703_start: Boolean;
            signal Xentry_3704_symbol: Boolean;
            signal Xexit_3705_symbol: Boolean;
            signal rr_3706_symbol : Boolean;
            signal ra_3707_symbol : Boolean;
            signal cr_3708_symbol : Boolean;
            signal ca_3709_symbol : Boolean;
            -- 
          begin -- 
            word_3_3703_start <= Xentry_3680_symbol; -- control passed to block
            Xentry_3704_symbol  <= word_3_3703_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3/$entry
            rr_3706_symbol <= Xentry_3704_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3/rr
            ptr_deref_549_addr_3_req_0 <= rr_3706_symbol; -- link to DP
            ra_3707_symbol <= ptr_deref_549_addr_3_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3/ra
            cr_3708_symbol <= ra_3707_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3/cr
            ptr_deref_549_addr_3_req_1 <= cr_3708_symbol; -- link to DP
            ca_3709_symbol <= ptr_deref_549_addr_3_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3/ca
            Xexit_3705_symbol <= ca_3709_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3/$exit
            word_3_3703_symbol <= Xexit_3705_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/word_3
          Xexit_3681_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/$exit 
            signal Xexit_3681_predecessors: BooleanArray(3 downto 0);
            -- 
          begin -- 
            Xexit_3681_predecessors(0) <= word_0_3682_symbol;
            Xexit_3681_predecessors(1) <= word_1_3689_symbol;
            Xexit_3681_predecessors(2) <= word_2_3696_symbol;
            Xexit_3681_predecessors(3) <= word_3_3703_symbol;
            Xexit_3681_join: join -- 
              port map( -- 
                preds => Xexit_3681_predecessors,
                symbol_out => Xexit_3681_symbol,
                clk => clk,
                reset => reset); -- 
            -- 
          end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/$exit
          ptr_deref_549_word_addrgen_3679_symbol <= Xexit_3681_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen
        ptr_deref_549_request_3710: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request 
          signal ptr_deref_549_request_3710_start: Boolean;
          signal Xentry_3711_symbol: Boolean;
          signal Xexit_3712_symbol: Boolean;
          signal word_access_3713_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_request_3710_start <= ptr_deref_549_trigger_x_x3662_symbol; -- control passed to block
          Xentry_3711_symbol  <= ptr_deref_549_request_3710_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/$entry
          word_access_3713: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access 
            signal word_access_3713_start: Boolean;
            signal Xentry_3714_symbol: Boolean;
            signal Xexit_3715_symbol: Boolean;
            signal word_access_0_3716_symbol : Boolean;
            signal word_access_1_3721_symbol : Boolean;
            signal word_access_2_3726_symbol : Boolean;
            signal word_access_3_3731_symbol : Boolean;
            -- 
          begin -- 
            word_access_3713_start <= Xentry_3711_symbol; -- control passed to block
            Xentry_3714_symbol  <= word_access_3713_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/$entry
            word_access_0_3716: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0 
              signal word_access_0_3716_start: Boolean;
              signal Xentry_3717_symbol: Boolean;
              signal Xexit_3718_symbol: Boolean;
              signal rr_3719_symbol : Boolean;
              signal ra_3720_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3716_start <= Xentry_3714_symbol; -- control passed to block
              Xentry_3717_symbol  <= word_access_0_3716_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/$entry
              rr_3719_symbol <= Xentry_3717_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/rr
              ptr_deref_549_load_0_req_0 <= rr_3719_symbol; -- link to DP
              ra_3720_symbol <= ptr_deref_549_load_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/ra
              Xexit_3718_symbol <= ra_3720_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/$exit
              word_access_0_3716_symbol <= Xexit_3718_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0
            word_access_1_3721: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_1 
              signal word_access_1_3721_start: Boolean;
              signal Xentry_3722_symbol: Boolean;
              signal Xexit_3723_symbol: Boolean;
              signal rr_3724_symbol : Boolean;
              signal ra_3725_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3721_start <= Xentry_3714_symbol; -- control passed to block
              Xentry_3722_symbol  <= word_access_1_3721_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_1/$entry
              rr_3724_symbol <= Xentry_3722_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_1/rr
              ptr_deref_549_load_1_req_0 <= rr_3724_symbol; -- link to DP
              ra_3725_symbol <= ptr_deref_549_load_1_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_1/ra
              Xexit_3723_symbol <= ra_3725_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_1/$exit
              word_access_1_3721_symbol <= Xexit_3723_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_1
            word_access_2_3726: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_2 
              signal word_access_2_3726_start: Boolean;
              signal Xentry_3727_symbol: Boolean;
              signal Xexit_3728_symbol: Boolean;
              signal rr_3729_symbol : Boolean;
              signal ra_3730_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3726_start <= Xentry_3714_symbol; -- control passed to block
              Xentry_3727_symbol  <= word_access_2_3726_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_2/$entry
              rr_3729_symbol <= Xentry_3727_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_2/rr
              ptr_deref_549_load_2_req_0 <= rr_3729_symbol; -- link to DP
              ra_3730_symbol <= ptr_deref_549_load_2_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_2/ra
              Xexit_3728_symbol <= ra_3730_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_2/$exit
              word_access_2_3726_symbol <= Xexit_3728_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_2
            word_access_3_3731: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_3 
              signal word_access_3_3731_start: Boolean;
              signal Xentry_3732_symbol: Boolean;
              signal Xexit_3733_symbol: Boolean;
              signal rr_3734_symbol : Boolean;
              signal ra_3735_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3731_start <= Xentry_3714_symbol; -- control passed to block
              Xentry_3732_symbol  <= word_access_3_3731_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_3/$entry
              rr_3734_symbol <= Xentry_3732_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_3/rr
              ptr_deref_549_load_3_req_0 <= rr_3734_symbol; -- link to DP
              ra_3735_symbol <= ptr_deref_549_load_3_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_3/ra
              Xexit_3733_symbol <= ra_3735_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_3/$exit
              word_access_3_3731_symbol <= Xexit_3733_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_3
            Xexit_3715_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/$exit 
              signal Xexit_3715_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3715_predecessors(0) <= word_access_0_3716_symbol;
              Xexit_3715_predecessors(1) <= word_access_1_3721_symbol;
              Xexit_3715_predecessors(2) <= word_access_2_3726_symbol;
              Xexit_3715_predecessors(3) <= word_access_3_3731_symbol;
              Xexit_3715_join: join -- 
                port map( -- 
                  preds => Xexit_3715_predecessors,
                  symbol_out => Xexit_3715_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/$exit
            word_access_3713_symbol <= Xexit_3715_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access
          Xexit_3712_symbol <= word_access_3713_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/$exit
          ptr_deref_549_request_3710_symbol <= Xexit_3712_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request
        ptr_deref_549_complete_3736: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete 
          signal ptr_deref_549_complete_3736_start: Boolean;
          signal Xentry_3737_symbol: Boolean;
          signal Xexit_3738_symbol: Boolean;
          signal word_access_3739_symbol : Boolean;
          signal merge_req_3762_symbol : Boolean;
          signal merge_ack_3763_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_complete_3736_start <= ptr_deref_549_active_x_x3663_symbol; -- control passed to block
          Xentry_3737_symbol  <= ptr_deref_549_complete_3736_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/$entry
          word_access_3739: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access 
            signal word_access_3739_start: Boolean;
            signal Xentry_3740_symbol: Boolean;
            signal Xexit_3741_symbol: Boolean;
            signal word_access_0_3742_symbol : Boolean;
            signal word_access_1_3747_symbol : Boolean;
            signal word_access_2_3752_symbol : Boolean;
            signal word_access_3_3757_symbol : Boolean;
            -- 
          begin -- 
            word_access_3739_start <= Xentry_3737_symbol; -- control passed to block
            Xentry_3740_symbol  <= word_access_3739_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/$entry
            word_access_0_3742: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0 
              signal word_access_0_3742_start: Boolean;
              signal Xentry_3743_symbol: Boolean;
              signal Xexit_3744_symbol: Boolean;
              signal cr_3745_symbol : Boolean;
              signal ca_3746_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3742_start <= Xentry_3740_symbol; -- control passed to block
              Xentry_3743_symbol  <= word_access_0_3742_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/$entry
              cr_3745_symbol <= Xentry_3743_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/cr
              ptr_deref_549_load_0_req_1 <= cr_3745_symbol; -- link to DP
              ca_3746_symbol <= ptr_deref_549_load_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/ca
              Xexit_3744_symbol <= ca_3746_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/$exit
              word_access_0_3742_symbol <= Xexit_3744_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0
            word_access_1_3747: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_1 
              signal word_access_1_3747_start: Boolean;
              signal Xentry_3748_symbol: Boolean;
              signal Xexit_3749_symbol: Boolean;
              signal cr_3750_symbol : Boolean;
              signal ca_3751_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3747_start <= Xentry_3740_symbol; -- control passed to block
              Xentry_3748_symbol  <= word_access_1_3747_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_1/$entry
              cr_3750_symbol <= Xentry_3748_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_1/cr
              ptr_deref_549_load_1_req_1 <= cr_3750_symbol; -- link to DP
              ca_3751_symbol <= ptr_deref_549_load_1_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_1/ca
              Xexit_3749_symbol <= ca_3751_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_1/$exit
              word_access_1_3747_symbol <= Xexit_3749_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_1
            word_access_2_3752: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_2 
              signal word_access_2_3752_start: Boolean;
              signal Xentry_3753_symbol: Boolean;
              signal Xexit_3754_symbol: Boolean;
              signal cr_3755_symbol : Boolean;
              signal ca_3756_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3752_start <= Xentry_3740_symbol; -- control passed to block
              Xentry_3753_symbol  <= word_access_2_3752_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_2/$entry
              cr_3755_symbol <= Xentry_3753_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_2/cr
              ptr_deref_549_load_2_req_1 <= cr_3755_symbol; -- link to DP
              ca_3756_symbol <= ptr_deref_549_load_2_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_2/ca
              Xexit_3754_symbol <= ca_3756_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_2/$exit
              word_access_2_3752_symbol <= Xexit_3754_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_2
            word_access_3_3757: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_3 
              signal word_access_3_3757_start: Boolean;
              signal Xentry_3758_symbol: Boolean;
              signal Xexit_3759_symbol: Boolean;
              signal cr_3760_symbol : Boolean;
              signal ca_3761_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3757_start <= Xentry_3740_symbol; -- control passed to block
              Xentry_3758_symbol  <= word_access_3_3757_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_3/$entry
              cr_3760_symbol <= Xentry_3758_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_3/cr
              ptr_deref_549_load_3_req_1 <= cr_3760_symbol; -- link to DP
              ca_3761_symbol <= ptr_deref_549_load_3_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_3/ca
              Xexit_3759_symbol <= ca_3761_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_3/$exit
              word_access_3_3757_symbol <= Xexit_3759_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_3
            Xexit_3741_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/$exit 
              signal Xexit_3741_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3741_predecessors(0) <= word_access_0_3742_symbol;
              Xexit_3741_predecessors(1) <= word_access_1_3747_symbol;
              Xexit_3741_predecessors(2) <= word_access_2_3752_symbol;
              Xexit_3741_predecessors(3) <= word_access_3_3757_symbol;
              Xexit_3741_join: join -- 
                port map( -- 
                  preds => Xexit_3741_predecessors,
                  symbol_out => Xexit_3741_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/$exit
            word_access_3739_symbol <= Xexit_3741_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access
          merge_req_3762_symbol <= word_access_3739_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/merge_req
          ptr_deref_549_gather_scatter_req_0 <= merge_req_3762_symbol; -- link to DP
          merge_ack_3763_symbol <= ptr_deref_549_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/merge_ack
          Xexit_3738_symbol <= merge_ack_3763_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/$exit
          ptr_deref_549_complete_3736_symbol <= Xexit_3738_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete
        Xexit_3501_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/$exit 
          signal Xexit_3501_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          Xexit_3501_predecessors(0) <= assign_stmt_537_completed_x_x3513_symbol;
          Xexit_3501_predecessors(1) <= ptr_deref_535_base_address_calculated_3517_symbol;
          Xexit_3501_predecessors(2) <= ptr_deref_540_base_address_calculated_3578_symbol;
          Xexit_3501_predecessors(3) <= assign_stmt_550_completed_x_x3661_symbol;
          Xexit_3501_join: join -- 
            port map( -- 
              preds => Xexit_3501_predecessors,
              symbol_out => Xexit_3501_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/$exit
        assign_stmt_533_to_assign_stmt_555_3499_symbol <= Xexit_3501_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555
      assign_stmt_559_3764: Block -- branch_block_stmt_513/assign_stmt_559 
        signal assign_stmt_559_3764_start: Boolean;
        signal Xentry_3765_symbol: Boolean;
        signal Xexit_3766_symbol: Boolean;
        signal assign_stmt_559_active_x_x3767_symbol : Boolean;
        signal assign_stmt_559_completed_x_x3768_symbol : Boolean;
        signal type_cast_558_active_x_x3769_symbol : Boolean;
        signal type_cast_558_trigger_x_x3770_symbol : Boolean;
        signal simple_obj_ref_557_complete_3771_symbol : Boolean;
        signal type_cast_558_complete_3772_symbol : Boolean;
        signal simple_obj_ref_556_trigger_x_x3777_symbol : Boolean;
        signal simple_obj_ref_556_complete_3778_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_559_3764_start <= assign_stmt_559_x_xentry_x_xx_x3464_symbol; -- control passed to block
        Xentry_3765_symbol  <= assign_stmt_559_3764_start; -- transition branch_block_stmt_513/assign_stmt_559/$entry
        assign_stmt_559_active_x_x3767_symbol <= type_cast_558_complete_3772_symbol; -- transition branch_block_stmt_513/assign_stmt_559/assign_stmt_559_active_
        assign_stmt_559_completed_x_x3768_symbol <= simple_obj_ref_556_complete_3778_symbol; -- transition branch_block_stmt_513/assign_stmt_559/assign_stmt_559_completed_
        type_cast_558_active_x_x3769_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_559/type_cast_558_active_ 
          signal type_cast_558_active_x_x3769_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_558_active_x_x3769_predecessors(0) <= type_cast_558_trigger_x_x3770_symbol;
          type_cast_558_active_x_x3769_predecessors(1) <= simple_obj_ref_557_complete_3771_symbol;
          type_cast_558_active_x_x3769_join: join -- 
            port map( -- 
              preds => type_cast_558_active_x_x3769_predecessors,
              symbol_out => type_cast_558_active_x_x3769_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_559/type_cast_558_active_
        type_cast_558_trigger_x_x3770_symbol <= Xentry_3765_symbol; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_trigger_
        simple_obj_ref_557_complete_3771_symbol <= Xentry_3765_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_557_complete
        type_cast_558_complete_3772: Block -- branch_block_stmt_513/assign_stmt_559/type_cast_558_complete 
          signal type_cast_558_complete_3772_start: Boolean;
          signal Xentry_3773_symbol: Boolean;
          signal Xexit_3774_symbol: Boolean;
          signal req_3775_symbol : Boolean;
          signal ack_3776_symbol : Boolean;
          -- 
        begin -- 
          type_cast_558_complete_3772_start <= type_cast_558_active_x_x3769_symbol; -- control passed to block
          Xentry_3773_symbol  <= type_cast_558_complete_3772_start; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/$entry
          req_3775_symbol <= Xentry_3773_symbol; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/req
          type_cast_558_inst_req_0 <= req_3775_symbol; -- link to DP
          ack_3776_symbol <= type_cast_558_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/ack
          Xexit_3774_symbol <= ack_3776_symbol; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/$exit
          type_cast_558_complete_3772_symbol <= Xexit_3774_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_559/type_cast_558_complete
        simple_obj_ref_556_trigger_x_x3777_symbol <= assign_stmt_559_active_x_x3767_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_trigger_
        simple_obj_ref_556_complete_3778: Block -- branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete 
          signal simple_obj_ref_556_complete_3778_start: Boolean;
          signal Xentry_3779_symbol: Boolean;
          signal Xexit_3780_symbol: Boolean;
          signal pipe_wreq_3781_symbol : Boolean;
          signal pipe_wack_3782_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_556_complete_3778_start <= simple_obj_ref_556_trigger_x_x3777_symbol; -- control passed to block
          Xentry_3779_symbol  <= simple_obj_ref_556_complete_3778_start; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/$entry
          pipe_wreq_3781_symbol <= Xentry_3779_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/pipe_wreq
          simple_obj_ref_556_inst_req_0 <= pipe_wreq_3781_symbol; -- link to DP
          pipe_wack_3782_symbol <= simple_obj_ref_556_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/pipe_wack
          Xexit_3780_symbol <= pipe_wack_3782_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/$exit
          simple_obj_ref_556_complete_3778_symbol <= Xexit_3780_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete
        Xexit_3766_symbol <= assign_stmt_559_completed_x_x3768_symbol; -- transition branch_block_stmt_513/assign_stmt_559/$exit
        assign_stmt_559_3764_symbol <= Xexit_3766_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_559
      assign_stmt_564_3783: Block -- branch_block_stmt_513/assign_stmt_564 
        signal assign_stmt_564_3783_start: Boolean;
        signal Xentry_3784_symbol: Boolean;
        signal Xexit_3785_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_564_3783_start <= assign_stmt_564_x_xentry_x_xx_x3466_symbol; -- control passed to block
        Xentry_3784_symbol  <= assign_stmt_564_3783_start; -- transition branch_block_stmt_513/assign_stmt_564/$entry
        Xexit_3785_symbol <= Xentry_3784_symbol; -- transition branch_block_stmt_513/assign_stmt_564/$exit
        assign_stmt_564_3783_symbol <= Xexit_3785_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_564
      assign_stmt_568_3786: Block -- branch_block_stmt_513/assign_stmt_568 
        signal assign_stmt_568_3786_start: Boolean;
        signal Xentry_3787_symbol: Boolean;
        signal Xexit_3788_symbol: Boolean;
        signal assign_stmt_568_active_x_x3789_symbol : Boolean;
        signal assign_stmt_568_completed_x_x3790_symbol : Boolean;
        signal simple_obj_ref_565_trigger_x_x3791_symbol : Boolean;
        signal simple_obj_ref_565_complete_3792_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_568_3786_start <= assign_stmt_568_x_xentry_x_xx_x3468_symbol; -- control passed to block
        Xentry_3787_symbol  <= assign_stmt_568_3786_start; -- transition branch_block_stmt_513/assign_stmt_568/$entry
        assign_stmt_568_active_x_x3789_symbol <= Xentry_3787_symbol; -- transition branch_block_stmt_513/assign_stmt_568/assign_stmt_568_active_
        assign_stmt_568_completed_x_x3790_symbol <= simple_obj_ref_565_complete_3792_symbol; -- transition branch_block_stmt_513/assign_stmt_568/assign_stmt_568_completed_
        simple_obj_ref_565_trigger_x_x3791_symbol <= assign_stmt_568_active_x_x3789_symbol; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_trigger_
        simple_obj_ref_565_complete_3792: Block -- branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete 
          signal simple_obj_ref_565_complete_3792_start: Boolean;
          signal Xentry_3793_symbol: Boolean;
          signal Xexit_3794_symbol: Boolean;
          signal pipe_wreq_3795_symbol : Boolean;
          signal pipe_wack_3796_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_565_complete_3792_start <= simple_obj_ref_565_trigger_x_x3791_symbol; -- control passed to block
          Xentry_3793_symbol  <= simple_obj_ref_565_complete_3792_start; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/$entry
          pipe_wreq_3795_symbol <= Xentry_3793_symbol; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/pipe_wreq
          simple_obj_ref_565_inst_req_0 <= pipe_wreq_3795_symbol; -- link to DP
          pipe_wack_3796_symbol <= simple_obj_ref_565_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/pipe_wack
          Xexit_3794_symbol <= pipe_wack_3796_symbol; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/$exit
          simple_obj_ref_565_complete_3792_symbol <= Xexit_3794_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete
        Xexit_3788_symbol <= assign_stmt_568_completed_x_x3790_symbol; -- transition branch_block_stmt_513/assign_stmt_568/$exit
        assign_stmt_568_3786_symbol <= Xexit_3788_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_568
      assign_stmt_572_to_assign_stmt_581_3797: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581 
        signal assign_stmt_572_to_assign_stmt_581_3797_start: Boolean;
        signal Xentry_3798_symbol: Boolean;
        signal Xexit_3799_symbol: Boolean;
        signal assign_stmt_572_active_x_x3800_symbol : Boolean;
        signal assign_stmt_572_completed_x_x3801_symbol : Boolean;
        signal ptr_deref_571_trigger_x_x3802_symbol : Boolean;
        signal ptr_deref_571_active_x_x3803_symbol : Boolean;
        signal ptr_deref_571_base_address_calculated_3804_symbol : Boolean;
        signal ptr_deref_571_root_address_calculated_3805_symbol : Boolean;
        signal ptr_deref_571_word_address_calculated_3806_symbol : Boolean;
        signal ptr_deref_571_request_3807_symbol : Boolean;
        signal ptr_deref_571_complete_3833_symbol : Boolean;
        signal assign_stmt_576_active_x_x3861_symbol : Boolean;
        signal assign_stmt_576_completed_x_x3862_symbol : Boolean;
        signal type_cast_575_active_x_x3863_symbol : Boolean;
        signal type_cast_575_trigger_x_x3864_symbol : Boolean;
        signal simple_obj_ref_574_complete_3865_symbol : Boolean;
        signal type_cast_575_complete_3866_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_572_to_assign_stmt_581_3797_start <= assign_stmt_572_to_assign_stmt_581_x_xentry_x_xx_x3470_symbol; -- control passed to block
        Xentry_3798_symbol  <= assign_stmt_572_to_assign_stmt_581_3797_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/$entry
        assign_stmt_572_active_x_x3800_symbol <= ptr_deref_571_complete_3833_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_572_active_
        assign_stmt_572_completed_x_x3801_symbol <= assign_stmt_572_active_x_x3800_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_572_completed_
        ptr_deref_571_trigger_x_x3802_symbol <= ptr_deref_571_word_address_calculated_3806_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_trigger_
        ptr_deref_571_active_x_x3803_symbol <= ptr_deref_571_request_3807_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_active_
        ptr_deref_571_base_address_calculated_3804_symbol <= Xentry_3798_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_base_address_calculated
        ptr_deref_571_root_address_calculated_3805_symbol <= Xentry_3798_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_root_address_calculated
        ptr_deref_571_word_address_calculated_3806_symbol <= ptr_deref_571_root_address_calculated_3805_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_word_address_calculated
        ptr_deref_571_request_3807: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request 
          signal ptr_deref_571_request_3807_start: Boolean;
          signal Xentry_3808_symbol: Boolean;
          signal Xexit_3809_symbol: Boolean;
          signal word_access_3810_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_571_request_3807_start <= ptr_deref_571_trigger_x_x3802_symbol; -- control passed to block
          Xentry_3808_symbol  <= ptr_deref_571_request_3807_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/$entry
          word_access_3810: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access 
            signal word_access_3810_start: Boolean;
            signal Xentry_3811_symbol: Boolean;
            signal Xexit_3812_symbol: Boolean;
            signal word_access_0_3813_symbol : Boolean;
            signal word_access_1_3818_symbol : Boolean;
            signal word_access_2_3823_symbol : Boolean;
            signal word_access_3_3828_symbol : Boolean;
            -- 
          begin -- 
            word_access_3810_start <= Xentry_3808_symbol; -- control passed to block
            Xentry_3811_symbol  <= word_access_3810_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/$entry
            word_access_0_3813: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0 
              signal word_access_0_3813_start: Boolean;
              signal Xentry_3814_symbol: Boolean;
              signal Xexit_3815_symbol: Boolean;
              signal rr_3816_symbol : Boolean;
              signal ra_3817_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3813_start <= Xentry_3811_symbol; -- control passed to block
              Xentry_3814_symbol  <= word_access_0_3813_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/$entry
              rr_3816_symbol <= Xentry_3814_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/rr
              ptr_deref_571_load_0_req_0 <= rr_3816_symbol; -- link to DP
              ra_3817_symbol <= ptr_deref_571_load_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/ra
              Xexit_3815_symbol <= ra_3817_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/$exit
              word_access_0_3813_symbol <= Xexit_3815_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0
            word_access_1_3818: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_1 
              signal word_access_1_3818_start: Boolean;
              signal Xentry_3819_symbol: Boolean;
              signal Xexit_3820_symbol: Boolean;
              signal rr_3821_symbol : Boolean;
              signal ra_3822_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3818_start <= Xentry_3811_symbol; -- control passed to block
              Xentry_3819_symbol  <= word_access_1_3818_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_1/$entry
              rr_3821_symbol <= Xentry_3819_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_1/rr
              ptr_deref_571_load_1_req_0 <= rr_3821_symbol; -- link to DP
              ra_3822_symbol <= ptr_deref_571_load_1_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_1/ra
              Xexit_3820_symbol <= ra_3822_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_1/$exit
              word_access_1_3818_symbol <= Xexit_3820_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_1
            word_access_2_3823: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_2 
              signal word_access_2_3823_start: Boolean;
              signal Xentry_3824_symbol: Boolean;
              signal Xexit_3825_symbol: Boolean;
              signal rr_3826_symbol : Boolean;
              signal ra_3827_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3823_start <= Xentry_3811_symbol; -- control passed to block
              Xentry_3824_symbol  <= word_access_2_3823_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_2/$entry
              rr_3826_symbol <= Xentry_3824_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_2/rr
              ptr_deref_571_load_2_req_0 <= rr_3826_symbol; -- link to DP
              ra_3827_symbol <= ptr_deref_571_load_2_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_2/ra
              Xexit_3825_symbol <= ra_3827_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_2/$exit
              word_access_2_3823_symbol <= Xexit_3825_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_2
            word_access_3_3828: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_3 
              signal word_access_3_3828_start: Boolean;
              signal Xentry_3829_symbol: Boolean;
              signal Xexit_3830_symbol: Boolean;
              signal rr_3831_symbol : Boolean;
              signal ra_3832_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3828_start <= Xentry_3811_symbol; -- control passed to block
              Xentry_3829_symbol  <= word_access_3_3828_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_3/$entry
              rr_3831_symbol <= Xentry_3829_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_3/rr
              ptr_deref_571_load_3_req_0 <= rr_3831_symbol; -- link to DP
              ra_3832_symbol <= ptr_deref_571_load_3_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_3/ra
              Xexit_3830_symbol <= ra_3832_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_3/$exit
              word_access_3_3828_symbol <= Xexit_3830_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_3
            Xexit_3812_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/$exit 
              signal Xexit_3812_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3812_predecessors(0) <= word_access_0_3813_symbol;
              Xexit_3812_predecessors(1) <= word_access_1_3818_symbol;
              Xexit_3812_predecessors(2) <= word_access_2_3823_symbol;
              Xexit_3812_predecessors(3) <= word_access_3_3828_symbol;
              Xexit_3812_join: join -- 
                port map( -- 
                  preds => Xexit_3812_predecessors,
                  symbol_out => Xexit_3812_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/$exit
            word_access_3810_symbol <= Xexit_3812_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access
          Xexit_3809_symbol <= word_access_3810_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/$exit
          ptr_deref_571_request_3807_symbol <= Xexit_3809_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request
        ptr_deref_571_complete_3833: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete 
          signal ptr_deref_571_complete_3833_start: Boolean;
          signal Xentry_3834_symbol: Boolean;
          signal Xexit_3835_symbol: Boolean;
          signal word_access_3836_symbol : Boolean;
          signal merge_req_3859_symbol : Boolean;
          signal merge_ack_3860_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_571_complete_3833_start <= ptr_deref_571_active_x_x3803_symbol; -- control passed to block
          Xentry_3834_symbol  <= ptr_deref_571_complete_3833_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/$entry
          word_access_3836: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access 
            signal word_access_3836_start: Boolean;
            signal Xentry_3837_symbol: Boolean;
            signal Xexit_3838_symbol: Boolean;
            signal word_access_0_3839_symbol : Boolean;
            signal word_access_1_3844_symbol : Boolean;
            signal word_access_2_3849_symbol : Boolean;
            signal word_access_3_3854_symbol : Boolean;
            -- 
          begin -- 
            word_access_3836_start <= Xentry_3834_symbol; -- control passed to block
            Xentry_3837_symbol  <= word_access_3836_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/$entry
            word_access_0_3839: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0 
              signal word_access_0_3839_start: Boolean;
              signal Xentry_3840_symbol: Boolean;
              signal Xexit_3841_symbol: Boolean;
              signal cr_3842_symbol : Boolean;
              signal ca_3843_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_3839_start <= Xentry_3837_symbol; -- control passed to block
              Xentry_3840_symbol  <= word_access_0_3839_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/$entry
              cr_3842_symbol <= Xentry_3840_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/cr
              ptr_deref_571_load_0_req_1 <= cr_3842_symbol; -- link to DP
              ca_3843_symbol <= ptr_deref_571_load_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/ca
              Xexit_3841_symbol <= ca_3843_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/$exit
              word_access_0_3839_symbol <= Xexit_3841_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0
            word_access_1_3844: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_1 
              signal word_access_1_3844_start: Boolean;
              signal Xentry_3845_symbol: Boolean;
              signal Xexit_3846_symbol: Boolean;
              signal cr_3847_symbol : Boolean;
              signal ca_3848_symbol : Boolean;
              -- 
            begin -- 
              word_access_1_3844_start <= Xentry_3837_symbol; -- control passed to block
              Xentry_3845_symbol  <= word_access_1_3844_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_1/$entry
              cr_3847_symbol <= Xentry_3845_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_1/cr
              ptr_deref_571_load_1_req_1 <= cr_3847_symbol; -- link to DP
              ca_3848_symbol <= ptr_deref_571_load_1_ack_1; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_1/ca
              Xexit_3846_symbol <= ca_3848_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_1/$exit
              word_access_1_3844_symbol <= Xexit_3846_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_1
            word_access_2_3849: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_2 
              signal word_access_2_3849_start: Boolean;
              signal Xentry_3850_symbol: Boolean;
              signal Xexit_3851_symbol: Boolean;
              signal cr_3852_symbol : Boolean;
              signal ca_3853_symbol : Boolean;
              -- 
            begin -- 
              word_access_2_3849_start <= Xentry_3837_symbol; -- control passed to block
              Xentry_3850_symbol  <= word_access_2_3849_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_2/$entry
              cr_3852_symbol <= Xentry_3850_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_2/cr
              ptr_deref_571_load_2_req_1 <= cr_3852_symbol; -- link to DP
              ca_3853_symbol <= ptr_deref_571_load_2_ack_1; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_2/ca
              Xexit_3851_symbol <= ca_3853_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_2/$exit
              word_access_2_3849_symbol <= Xexit_3851_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_2
            word_access_3_3854: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_3 
              signal word_access_3_3854_start: Boolean;
              signal Xentry_3855_symbol: Boolean;
              signal Xexit_3856_symbol: Boolean;
              signal cr_3857_symbol : Boolean;
              signal ca_3858_symbol : Boolean;
              -- 
            begin -- 
              word_access_3_3854_start <= Xentry_3837_symbol; -- control passed to block
              Xentry_3855_symbol  <= word_access_3_3854_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_3/$entry
              cr_3857_symbol <= Xentry_3855_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_3/cr
              ptr_deref_571_load_3_req_1 <= cr_3857_symbol; -- link to DP
              ca_3858_symbol <= ptr_deref_571_load_3_ack_1; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_3/ca
              Xexit_3856_symbol <= ca_3858_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_3/$exit
              word_access_3_3854_symbol <= Xexit_3856_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_3
            Xexit_3838_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/$exit 
              signal Xexit_3838_predecessors: BooleanArray(3 downto 0);
              -- 
            begin -- 
              Xexit_3838_predecessors(0) <= word_access_0_3839_symbol;
              Xexit_3838_predecessors(1) <= word_access_1_3844_symbol;
              Xexit_3838_predecessors(2) <= word_access_2_3849_symbol;
              Xexit_3838_predecessors(3) <= word_access_3_3854_symbol;
              Xexit_3838_join: join -- 
                port map( -- 
                  preds => Xexit_3838_predecessors,
                  symbol_out => Xexit_3838_symbol,
                  clk => clk,
                  reset => reset); -- 
              -- 
            end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/$exit
            word_access_3836_symbol <= Xexit_3838_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access
          merge_req_3859_symbol <= word_access_3836_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/merge_req
          ptr_deref_571_gather_scatter_req_0 <= merge_req_3859_symbol; -- link to DP
          merge_ack_3860_symbol <= ptr_deref_571_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/merge_ack
          Xexit_3835_symbol <= merge_ack_3860_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/$exit
          ptr_deref_571_complete_3833_symbol <= Xexit_3835_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete
        assign_stmt_576_active_x_x3861_symbol <= type_cast_575_complete_3866_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_576_active_
        assign_stmt_576_completed_x_x3862_symbol <= assign_stmt_576_active_x_x3861_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_576_completed_
        type_cast_575_active_x_x3863_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_active_ 
          signal type_cast_575_active_x_x3863_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_575_active_x_x3863_predecessors(0) <= type_cast_575_trigger_x_x3864_symbol;
          type_cast_575_active_x_x3863_predecessors(1) <= simple_obj_ref_574_complete_3865_symbol;
          type_cast_575_active_x_x3863_join: join -- 
            port map( -- 
              preds => type_cast_575_active_x_x3863_predecessors,
              symbol_out => type_cast_575_active_x_x3863_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_active_
        type_cast_575_trigger_x_x3864_symbol <= Xentry_3798_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_trigger_
        simple_obj_ref_574_complete_3865_symbol <= assign_stmt_572_completed_x_x3801_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/simple_obj_ref_574_complete
        type_cast_575_complete_3866: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete 
          signal type_cast_575_complete_3866_start: Boolean;
          signal Xentry_3867_symbol: Boolean;
          signal Xexit_3868_symbol: Boolean;
          signal req_3869_symbol : Boolean;
          signal ack_3870_symbol : Boolean;
          -- 
        begin -- 
          type_cast_575_complete_3866_start <= type_cast_575_active_x_x3863_symbol; -- control passed to block
          Xentry_3867_symbol  <= type_cast_575_complete_3866_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/$entry
          req_3869_symbol <= Xentry_3867_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/req
          type_cast_575_inst_req_0 <= req_3869_symbol; -- link to DP
          ack_3870_symbol <= type_cast_575_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/ack
          Xexit_3868_symbol <= ack_3870_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/$exit
          type_cast_575_complete_3866_symbol <= Xexit_3868_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete
        Xexit_3799_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/$exit 
          signal Xexit_3799_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_3799_predecessors(0) <= ptr_deref_571_base_address_calculated_3804_symbol;
          Xexit_3799_predecessors(1) <= assign_stmt_576_completed_x_x3862_symbol;
          Xexit_3799_join: join -- 
            port map( -- 
              preds => Xexit_3799_predecessors,
              symbol_out => Xexit_3799_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/$exit
        assign_stmt_572_to_assign_stmt_581_3797_symbol <= Xexit_3799_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581
      assign_stmt_585_3871: Block -- branch_block_stmt_513/assign_stmt_585 
        signal assign_stmt_585_3871_start: Boolean;
        signal Xentry_3872_symbol: Boolean;
        signal Xexit_3873_symbol: Boolean;
        signal assign_stmt_585_active_x_x3874_symbol : Boolean;
        signal assign_stmt_585_completed_x_x3875_symbol : Boolean;
        signal type_cast_584_active_x_x3876_symbol : Boolean;
        signal type_cast_584_trigger_x_x3877_symbol : Boolean;
        signal simple_obj_ref_583_complete_3878_symbol : Boolean;
        signal type_cast_584_complete_3879_symbol : Boolean;
        signal simple_obj_ref_582_trigger_x_x3884_symbol : Boolean;
        signal simple_obj_ref_582_complete_3885_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_585_3871_start <= assign_stmt_585_x_xentry_x_xx_x3472_symbol; -- control passed to block
        Xentry_3872_symbol  <= assign_stmt_585_3871_start; -- transition branch_block_stmt_513/assign_stmt_585/$entry
        assign_stmt_585_active_x_x3874_symbol <= type_cast_584_complete_3879_symbol; -- transition branch_block_stmt_513/assign_stmt_585/assign_stmt_585_active_
        assign_stmt_585_completed_x_x3875_symbol <= simple_obj_ref_582_complete_3885_symbol; -- transition branch_block_stmt_513/assign_stmt_585/assign_stmt_585_completed_
        type_cast_584_active_x_x3876_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_585/type_cast_584_active_ 
          signal type_cast_584_active_x_x3876_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_584_active_x_x3876_predecessors(0) <= type_cast_584_trigger_x_x3877_symbol;
          type_cast_584_active_x_x3876_predecessors(1) <= simple_obj_ref_583_complete_3878_symbol;
          type_cast_584_active_x_x3876_join: join -- 
            port map( -- 
              preds => type_cast_584_active_x_x3876_predecessors,
              symbol_out => type_cast_584_active_x_x3876_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_585/type_cast_584_active_
        type_cast_584_trigger_x_x3877_symbol <= Xentry_3872_symbol; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_trigger_
        simple_obj_ref_583_complete_3878_symbol <= Xentry_3872_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_583_complete
        type_cast_584_complete_3879: Block -- branch_block_stmt_513/assign_stmt_585/type_cast_584_complete 
          signal type_cast_584_complete_3879_start: Boolean;
          signal Xentry_3880_symbol: Boolean;
          signal Xexit_3881_symbol: Boolean;
          signal req_3882_symbol : Boolean;
          signal ack_3883_symbol : Boolean;
          -- 
        begin -- 
          type_cast_584_complete_3879_start <= type_cast_584_active_x_x3876_symbol; -- control passed to block
          Xentry_3880_symbol  <= type_cast_584_complete_3879_start; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/$entry
          req_3882_symbol <= Xentry_3880_symbol; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/req
          type_cast_584_inst_req_0 <= req_3882_symbol; -- link to DP
          ack_3883_symbol <= type_cast_584_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/ack
          Xexit_3881_symbol <= ack_3883_symbol; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/$exit
          type_cast_584_complete_3879_symbol <= Xexit_3881_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_585/type_cast_584_complete
        simple_obj_ref_582_trigger_x_x3884_symbol <= assign_stmt_585_active_x_x3874_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_trigger_
        simple_obj_ref_582_complete_3885: Block -- branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete 
          signal simple_obj_ref_582_complete_3885_start: Boolean;
          signal Xentry_3886_symbol: Boolean;
          signal Xexit_3887_symbol: Boolean;
          signal pipe_wreq_3888_symbol : Boolean;
          signal pipe_wack_3889_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_582_complete_3885_start <= simple_obj_ref_582_trigger_x_x3884_symbol; -- control passed to block
          Xentry_3886_symbol  <= simple_obj_ref_582_complete_3885_start; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/$entry
          pipe_wreq_3888_symbol <= Xentry_3886_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/pipe_wreq
          simple_obj_ref_582_inst_req_0 <= pipe_wreq_3888_symbol; -- link to DP
          pipe_wack_3889_symbol <= simple_obj_ref_582_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/pipe_wack
          Xexit_3887_symbol <= pipe_wack_3889_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/$exit
          simple_obj_ref_582_complete_3885_symbol <= Xexit_3887_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete
        Xexit_3873_symbol <= assign_stmt_585_completed_x_x3875_symbol; -- transition branch_block_stmt_513/assign_stmt_585/$exit
        assign_stmt_585_3871_symbol <= Xexit_3873_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_585
      bb_0_bb_1_PhiReq_3890: Block -- branch_block_stmt_513/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_3890_start: Boolean;
        signal Xentry_3891_symbol: Boolean;
        signal Xexit_3892_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_3890_start <= bb_0_bb_1_3456_symbol; -- control passed to block
        Xentry_3891_symbol  <= bb_0_bb_1_PhiReq_3890_start; -- transition branch_block_stmt_513/bb_0_bb_1_PhiReq/$entry
        Xexit_3892_symbol <= Xentry_3891_symbol; -- transition branch_block_stmt_513/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_3890_symbol <= Xexit_3892_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/bb_0_bb_1_PhiReq
      bb_1_bb_1_PhiReq_3893: Block -- branch_block_stmt_513/bb_1_bb_1_PhiReq 
        signal bb_1_bb_1_PhiReq_3893_start: Boolean;
        signal Xentry_3894_symbol: Boolean;
        signal Xexit_3895_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_1_PhiReq_3893_start <= bb_1_bb_1_3474_symbol; -- control passed to block
        Xentry_3894_symbol  <= bb_1_bb_1_PhiReq_3893_start; -- transition branch_block_stmt_513/bb_1_bb_1_PhiReq/$entry
        Xexit_3895_symbol <= Xentry_3894_symbol; -- transition branch_block_stmt_513/bb_1_bb_1_PhiReq/$exit
        bb_1_bb_1_PhiReq_3893_symbol <= Xexit_3895_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/bb_1_bb_1_PhiReq
      merge_stmt_520_PhiReqMerge_3896_symbol  <=  bb_0_bb_1_PhiReq_3890_symbol or bb_1_bb_1_PhiReq_3893_symbol; -- place branch_block_stmt_513/merge_stmt_520_PhiReqMerge (optimized away) 
      merge_stmt_520_PhiAck_3897: Block -- branch_block_stmt_513/merge_stmt_520_PhiAck 
        signal merge_stmt_520_PhiAck_3897_start: Boolean;
        signal Xentry_3898_symbol: Boolean;
        signal Xexit_3899_symbol: Boolean;
        signal dummy_3900_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_520_PhiAck_3897_start <= merge_stmt_520_PhiReqMerge_3896_symbol; -- control passed to block
        Xentry_3898_symbol  <= merge_stmt_520_PhiAck_3897_start; -- transition branch_block_stmt_513/merge_stmt_520_PhiAck/$entry
        dummy_3900_symbol <= Xentry_3898_symbol; -- transition branch_block_stmt_513/merge_stmt_520_PhiAck/dummy
        Xexit_3899_symbol <= dummy_3900_symbol; -- transition branch_block_stmt_513/merge_stmt_520_PhiAck/$exit
        merge_stmt_520_PhiAck_3897_symbol <= Xexit_3899_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/merge_stmt_520_PhiAck
      Xexit_3451_symbol <= branch_block_stmt_513_x_xexit_x_xx_x3453_symbol; -- transition branch_block_stmt_513/$exit
      branch_block_stmt_513_3449_symbol <= Xexit_3451_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_513
    Xexit_3448_symbol <= branch_block_stmt_513_3449_symbol; -- transition $exit
    fin  <=  '1' when Xexit_3448_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_545_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_545_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_545_root_address : std_logic_vector(5 downto 0);
    signal iNsTr_10_564 : std_logic_vector(31 downto 0);
    signal iNsTr_12_572 : std_logic_vector(31 downto 0);
    signal iNsTr_13_576 : std_logic_vector(31 downto 0);
    signal iNsTr_14_581 : std_logic_vector(31 downto 0);
    signal iNsTr_1_525 : std_logic_vector(31 downto 0);
    signal iNsTr_2_529 : std_logic_vector(31 downto 0);
    signal iNsTr_3_533 : std_logic_vector(31 downto 0);
    signal iNsTr_5_541 : std_logic_vector(31 downto 0);
    signal iNsTr_6_546 : std_logic_vector(31 downto 0);
    signal iNsTr_7_550 : std_logic_vector(31 downto 0);
    signal iNsTr_8_555 : std_logic_vector(31 downto 0);
    signal lptr_518 : std_logic_vector(31 downto 0);
    signal ptr_deref_535_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_535_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_535_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_535_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_535_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_535_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_535_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_535_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_535_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_540_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_540_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_540_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_540_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_540_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_540_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_540_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_540_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_549_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_549_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_549_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_549_resized_base_address : std_logic_vector(5 downto 0);
    signal ptr_deref_549_root_address : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_address_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_offset_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_offset_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_offset_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_549_word_offset_3 : std_logic_vector(5 downto 0);
    signal ptr_deref_571_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_571_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_571_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_571_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_571_word_address_0 : std_logic_vector(5 downto 0);
    signal ptr_deref_571_word_address_1 : std_logic_vector(5 downto 0);
    signal ptr_deref_571_word_address_2 : std_logic_vector(5 downto 0);
    signal ptr_deref_571_word_address_3 : std_logic_vector(5 downto 0);
    signal simple_obj_ref_527_wire : std_logic_vector(31 downto 0);
    signal type_cast_558_wire : std_logic_vector(31 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_584_wire : std_logic_vector(31 downto 0);
    signal xxoutput_modulexxbodyxxlptr_alloc_base_address : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    array_obj_ref_545_final_offset <= "000100";
    iNsTr_10_564 <= "00000000000000000000000000000000";
    iNsTr_14_581 <= "00000000000000000000000000000000";
    iNsTr_1_525 <= "00000000000000000000000000000000";
    iNsTr_8_555 <= "00000000000000000000000000000000";
    lptr_518 <= "00000000000000000000000000110001";
    ptr_deref_535_word_address_0 <= "110001";
    ptr_deref_535_word_address_1 <= "110010";
    ptr_deref_535_word_address_2 <= "110011";
    ptr_deref_535_word_address_3 <= "110100";
    ptr_deref_540_word_address_0 <= "110001";
    ptr_deref_540_word_address_1 <= "110010";
    ptr_deref_540_word_address_2 <= "110011";
    ptr_deref_540_word_address_3 <= "110100";
    ptr_deref_549_word_offset_0 <= "000000";
    ptr_deref_549_word_offset_1 <= "000001";
    ptr_deref_549_word_offset_2 <= "000010";
    ptr_deref_549_word_offset_3 <= "000011";
    ptr_deref_571_word_address_0 <= "110001";
    ptr_deref_571_word_address_1 <= "110010";
    ptr_deref_571_word_address_2 <= "110011";
    ptr_deref_571_word_address_3 <= "110100";
    type_cast_567_wire_constant <= "00000001";
    xxoutput_modulexxbodyxxlptr_alloc_base_address <= "110001";
    array_obj_ref_545_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_5_541, dout => array_obj_ref_545_resized_base_address, req => array_obj_ref_545_base_resize_req_0, ack => array_obj_ref_545_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_545_final_reg: RegisterBase generic map(in_data_width => 6,out_data_width => 32) -- 
      port map( din => array_obj_ref_545_root_address, dout => iNsTr_6_546, req => array_obj_ref_545_final_reg_req_0, ack => array_obj_ref_545_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_549_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 6) -- 
      port map( din => iNsTr_6_546, dout => ptr_deref_549_resized_base_address, req => ptr_deref_549_base_resize_req_0, ack => ptr_deref_549_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_528_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_527_wire, dout => iNsTr_2_529, req => type_cast_528_inst_req_0, ack => type_cast_528_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_532_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_2_529, dout => iNsTr_3_533, req => type_cast_532_inst_req_0, ack => type_cast_532_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_558_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_7_550, dout => type_cast_558_wire, req => type_cast_558_inst_req_0, ack => type_cast_558_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_575_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_12_572, dout => iNsTr_13_576, req => type_cast_575_inst_req_0, ack => type_cast_575_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_584_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_13_576, dout => type_cast_584_wire, req => type_cast_584_inst_req_0, ack => type_cast_584_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_535_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_535_gather_scatter_ack_0 <= ptr_deref_535_gather_scatter_req_0;
      aggregated_sig <= iNsTr_3_533;
      ptr_deref_535_data_0 <= aggregated_sig(31 downto 24);
      ptr_deref_535_data_1 <= aggregated_sig(23 downto 16);
      ptr_deref_535_data_2 <= aggregated_sig(15 downto 8);
      ptr_deref_535_data_3 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_540_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_540_gather_scatter_ack_0 <= ptr_deref_540_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_540_data_0 & ptr_deref_540_data_1 & ptr_deref_540_data_2 & ptr_deref_540_data_3;
      iNsTr_5_541 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_549_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_549_gather_scatter_ack_0 <= ptr_deref_549_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_549_data_0 & ptr_deref_549_data_1 & ptr_deref_549_data_2 & ptr_deref_549_data_3;
      iNsTr_7_550 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_549_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(5 downto 0); --
    begin -- 
      ptr_deref_549_root_address_inst_ack_0 <= ptr_deref_549_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_549_resized_base_address;
      ptr_deref_549_root_address <= aggregated_sig(5 downto 0);
      --
    end Block;
    ptr_deref_571_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_571_gather_scatter_ack_0 <= ptr_deref_571_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_571_data_0 & ptr_deref_571_data_1 & ptr_deref_571_data_2 & ptr_deref_571_data_3;
      iNsTr_12_572 <= aggregated_sig(31 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_545_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_545_resized_base_address;
      array_obj_ref_545_root_address <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000100",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_545_root_address_inst_req_0,
          ackL => array_obj_ref_545_root_address_inst_ack_0,
          reqR => array_obj_ref_545_root_address_inst_req_1,
          ackR => array_obj_ref_545_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ptr_deref_549_addr_0 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_549_root_address;
      ptr_deref_549_word_address_0 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_549_addr_0_req_0,
          ackL => ptr_deref_549_addr_0_ack_0,
          reqR => ptr_deref_549_addr_0_req_1,
          ackR => ptr_deref_549_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ptr_deref_549_addr_1 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_549_root_address;
      ptr_deref_549_word_address_1 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_549_addr_1_req_0,
          ackL => ptr_deref_549_addr_1_ack_0,
          reqR => ptr_deref_549_addr_1_req_1,
          ackR => ptr_deref_549_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ptr_deref_549_addr_2 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_549_root_address;
      ptr_deref_549_word_address_2 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_549_addr_2_req_0,
          ackL => ptr_deref_549_addr_2_ack_0,
          reqR => ptr_deref_549_addr_2_req_1,
          ackR => ptr_deref_549_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ptr_deref_549_addr_3 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_549_root_address;
      ptr_deref_549_word_address_3 <= data_out(5 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000011",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_549_addr_3_req_0,
          ackL => ptr_deref_549_addr_3_ack_0,
          reqR => ptr_deref_549_addr_3_req_1,
          ackR => ptr_deref_549_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared load operator group (0) : ptr_deref_571_load_0 ptr_deref_540_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_571_load_0_req_0;
      reqL(0) <= ptr_deref_540_load_0_req_0;
      ptr_deref_571_load_0_ack_0 <= ackL(1);
      ptr_deref_540_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_571_load_0_req_1;
      reqR(0) <= ptr_deref_540_load_0_req_1;
      ptr_deref_571_load_0_ack_1 <= ackR(1);
      ptr_deref_540_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_571_word_address_0 & ptr_deref_540_word_address_0;
      ptr_deref_571_data_0 <= data_out(15 downto 8);
      ptr_deref_540_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(7),
          mack => memory_space_1_lr_ack(7),
          maddr => memory_space_1_lr_addr(47 downto 42),
          mtag => memory_space_1_lr_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(7),
          mack => memory_space_1_lc_ack(7),
          mdata => memory_space_1_lc_data(63 downto 56),
          mtag => memory_space_1_lc_tag(23 downto 21),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_540_load_1 ptr_deref_571_load_1 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_540_load_1_req_0;
      reqL(0) <= ptr_deref_571_load_1_req_0;
      ptr_deref_540_load_1_ack_0 <= ackL(1);
      ptr_deref_571_load_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_540_load_1_req_1;
      reqR(0) <= ptr_deref_571_load_1_req_1;
      ptr_deref_540_load_1_ack_1 <= ackR(1);
      ptr_deref_571_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_540_word_address_1 & ptr_deref_571_word_address_1;
      ptr_deref_540_data_1 <= data_out(15 downto 8);
      ptr_deref_571_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(6),
          mack => memory_space_1_lr_ack(6),
          maddr => memory_space_1_lr_addr(41 downto 36),
          mtag => memory_space_1_lr_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(6),
          mack => memory_space_1_lc_ack(6),
          mdata => memory_space_1_lc_data(55 downto 48),
          mtag => memory_space_1_lc_tag(20 downto 18),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_571_load_2 ptr_deref_540_load_2 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_571_load_2_req_0;
      reqL(0) <= ptr_deref_540_load_2_req_0;
      ptr_deref_571_load_2_ack_0 <= ackL(1);
      ptr_deref_540_load_2_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_571_load_2_req_1;
      reqR(0) <= ptr_deref_540_load_2_req_1;
      ptr_deref_571_load_2_ack_1 <= ackR(1);
      ptr_deref_540_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_571_word_address_2 & ptr_deref_540_word_address_2;
      ptr_deref_571_data_2 <= data_out(15 downto 8);
      ptr_deref_540_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(5),
          mack => memory_space_1_lr_ack(5),
          maddr => memory_space_1_lr_addr(35 downto 30),
          mtag => memory_space_1_lr_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(5),
          mack => memory_space_1_lc_ack(5),
          mdata => memory_space_1_lc_data(47 downto 40),
          mtag => memory_space_1_lc_tag(17 downto 15),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_571_load_3 ptr_deref_540_load_3 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_571_load_3_req_0;
      reqL(0) <= ptr_deref_540_load_3_req_0;
      ptr_deref_571_load_3_ack_0 <= ackL(1);
      ptr_deref_540_load_3_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_571_load_3_req_1;
      reqR(0) <= ptr_deref_540_load_3_req_1;
      ptr_deref_571_load_3_ack_1 <= ackR(1);
      ptr_deref_540_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_571_word_address_3 & ptr_deref_540_word_address_3;
      ptr_deref_571_data_3 <= data_out(15 downto 8);
      ptr_deref_540_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(4),
          mack => memory_space_1_lr_ack(4),
          maddr => memory_space_1_lr_addr(29 downto 24),
          mtag => memory_space_1_lr_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(4),
          mack => memory_space_1_lc_ack(4),
          mdata => memory_space_1_lc_data(39 downto 32),
          mtag => memory_space_1_lc_tag(14 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_549_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_549_load_0_req_0;
      ptr_deref_549_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_549_load_0_req_1;
      ptr_deref_549_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_549_word_address_0;
      ptr_deref_549_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(3),
          mack => memory_space_1_lr_ack(3),
          maddr => memory_space_1_lr_addr(23 downto 18),
          mtag => memory_space_1_lr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(3),
          mack => memory_space_1_lc_ack(3),
          mdata => memory_space_1_lc_data(31 downto 24),
          mtag => memory_space_1_lc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_549_load_1 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_549_load_1_req_0;
      ptr_deref_549_load_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_549_load_1_req_1;
      ptr_deref_549_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_549_word_address_1;
      ptr_deref_549_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(2),
          mack => memory_space_1_lr_ack(2),
          maddr => memory_space_1_lr_addr(17 downto 12),
          mtag => memory_space_1_lr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(2),
          mack => memory_space_1_lc_ack(2),
          mdata => memory_space_1_lc_data(23 downto 16),
          mtag => memory_space_1_lc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_549_load_2 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_549_load_2_req_0;
      ptr_deref_549_load_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_549_load_2_req_1;
      ptr_deref_549_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_549_word_address_2;
      ptr_deref_549_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(1),
          mack => memory_space_1_lr_ack(1),
          maddr => memory_space_1_lr_addr(11 downto 6),
          mtag => memory_space_1_lr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(1),
          mack => memory_space_1_lc_ack(1),
          mdata => memory_space_1_lc_data(15 downto 8),
          mtag => memory_space_1_lc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_549_load_3 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_549_load_3_req_0;
      ptr_deref_549_load_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_549_load_3_req_1;
      ptr_deref_549_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_549_word_address_3;
      ptr_deref_549_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 6,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(5 downto 0),
          mtag => memory_space_1_lr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 3,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared store operator group (0) : ptr_deref_535_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_535_store_0_req_0;
      ptr_deref_535_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_535_store_0_req_1;
      ptr_deref_535_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_535_word_address_0;
      data_in <= ptr_deref_535_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(3),
          mack => memory_space_1_sr_ack(3),
          maddr => memory_space_1_sr_addr(23 downto 18),
          mdata => memory_space_1_sr_data(31 downto 24),
          mtag => memory_space_1_sr_tag(11 downto 9),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(3),
          mack => memory_space_1_sc_ack(3),
          mtag => memory_space_1_sc_tag(11 downto 9),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_535_store_1 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_535_store_1_req_0;
      ptr_deref_535_store_1_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_535_store_1_req_1;
      ptr_deref_535_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_535_word_address_1;
      data_in <= ptr_deref_535_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(2),
          mack => memory_space_1_sr_ack(2),
          maddr => memory_space_1_sr_addr(17 downto 12),
          mdata => memory_space_1_sr_data(23 downto 16),
          mtag => memory_space_1_sr_tag(8 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(2),
          mack => memory_space_1_sc_ack(2),
          mtag => memory_space_1_sc_tag(8 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_535_store_2 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_535_store_2_req_0;
      ptr_deref_535_store_2_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_535_store_2_req_1;
      ptr_deref_535_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_535_word_address_2;
      data_in <= ptr_deref_535_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(1),
          mack => memory_space_1_sr_ack(1),
          maddr => memory_space_1_sr_addr(11 downto 6),
          mdata => memory_space_1_sr_data(15 downto 8),
          mtag => memory_space_1_sr_tag(5 downto 3),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(1),
          mack => memory_space_1_sc_ack(1),
          mtag => memory_space_1_sc_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_535_store_3 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_535_store_3_req_0;
      ptr_deref_535_store_3_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_535_store_3_req_1;
      ptr_deref_535_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_535_word_address_3;
      data_in <= ptr_deref_535_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 6,
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(5 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(2 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : simple_obj_ref_527_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_527_inst_req_0;
      simple_obj_ref_527_inst_ack_0 <= ack(0);
      simple_obj_ref_527_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => foo_out_pipe_read_req(0),
          oack => foo_out_pipe_read_ack(0),
          odata => foo_out_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : simple_obj_ref_556_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_556_inst_req_0;
      simple_obj_ref_556_inst_ack_0 <= ack(0);
      data_in <= type_cast_558_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => output_data_pipe_write_req(0),
          oack => output_data_pipe_write_ack(0),
          odata => output_data_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_565_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_565_inst_req_0;
      simple_obj_ref_565_inst_ack_0 <= ack(0);
      data_in <= type_cast_567_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_582_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_582_inst_req_0;
      simple_obj_ref_582_inst_ack_0 <= ack(0);
      data_in <= type_cast_584_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_put_pipe_write_req(0),
          oack => free_queue_put_pipe_write_ack(0),
          odata => free_queue_put_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity test_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    input_data_pipe_write_data: in std_logic_vector(31 downto 0);
    input_data_pipe_write_req : in std_logic_vector(0 downto 0);
    input_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    output_data_pipe_read_data: out std_logic_vector(31 downto 0);
    output_data_pipe_read_req : in std_logic_vector(0 downto 0);
    output_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of test_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(47 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(47 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(287 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(143 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(47 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(47 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(383 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(143 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(27 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(27 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(167 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(223 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(83 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(27 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(27 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(83 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  -- interface signals to connect to memory space memory_space_4
  -- interface signals to connect to memory space memory_space_5
  -- interface signals to connect to memory space memory_space_6
  -- interface signals to connect to memory space memory_space_7
  -- interface signals to connect to memory space memory_space_8
  -- interface signals to connect to memory space memory_space_9
  -- declarations related to module foo
  component foo is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(15 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(15 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(95 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(47 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(15 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(127 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(47 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(47 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(23 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(7 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(23 downto 0);
      foo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      foo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      foo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      foo_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      foo_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      foo_out_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module foo
  signal foo_tag_in    : std_logic_vector(0 downto 0);
  signal foo_tag_out   : std_logic_vector(0 downto 0);
  signal foo_start : std_logic;
  signal foo_fin   : std_logic;
  -- declarations related to module free_queue_manager
  component free_queue_manager is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(1 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(1 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(1 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(1 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(1 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(11 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(11 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(71 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(35 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(11 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(11 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(95 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(35 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(47 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(23 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(7 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(23 downto 0);
      free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_manager
  signal free_queue_manager_tag_in    : std_logic_vector(0 downto 0);
  signal free_queue_manager_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_manager_start : std_logic;
  signal free_queue_manager_fin   : std_logic;
  -- declarations related to module input_module
  component input_module is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(11 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(11 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(71 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(35 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(11 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(11 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(95 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(35 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(47 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(23 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(7 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(23 downto 0);
      free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      foo_in_pipe_write_req : out  std_logic_vector(0 downto 0);
      foo_in_pipe_write_ack : in   std_logic_vector(0 downto 0);
      foo_in_pipe_write_data : out  std_logic_vector(31 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module input_module
  signal input_module_tag_in    : std_logic_vector(0 downto 0);
  signal input_module_tag_out   : std_logic_vector(0 downto 0);
  signal input_module_start : std_logic;
  signal input_module_fin   : std_logic;
  -- declarations related to module mem_load_x_x
  component mem_load_x_x is -- 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(7 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module mem_load_x_x
  signal mem_load_x_x_address :  std_logic_vector(31 downto 0);
  signal mem_load_x_x_data :  std_logic_vector(7 downto 0);
  signal mem_load_x_x_in_args    : std_logic_vector(31 downto 0);
  signal mem_load_x_x_out_args   : std_logic_vector(7 downto 0);
  signal mem_load_x_x_tag_in    : std_logic_vector(0 downto 0);
  signal mem_load_x_x_tag_out   : std_logic_vector(0 downto 0);
  signal mem_load_x_x_start : std_logic;
  signal mem_load_x_x_fin   : std_logic;
  -- declarations related to module mem_store_x_x
  component mem_store_x_x is -- 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(7 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module mem_store_x_x
  signal mem_store_x_x_address :  std_logic_vector(31 downto 0);
  signal mem_store_x_x_data :  std_logic_vector(7 downto 0);
  signal mem_store_x_x_in_args    : std_logic_vector(39 downto 0);
  signal mem_store_x_x_tag_in    : std_logic_vector(0 downto 0);
  signal mem_store_x_x_tag_out   : std_logic_vector(0 downto 0);
  signal mem_store_x_x_start : std_logic;
  signal mem_store_x_x_fin   : std_logic;
  -- declarations related to module output_module
  component output_module is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(47 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(23 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(7 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(23 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(3 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(23 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(11 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(3 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(3 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(11 downto 0);
      foo_out_pipe_read_req : out  std_logic_vector(0 downto 0);
      foo_out_pipe_read_ack : in   std_logic_vector(0 downto 0);
      foo_out_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_data_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module output_module
  signal output_module_tag_in    : std_logic_vector(0 downto 0);
  signal output_module_tag_out   : std_logic_vector(0 downto 0);
  signal output_module_start : std_logic;
  signal output_module_fin   : std_logic;
  -- aggregate signals for write to pipe foo_in
  signal foo_in_pipe_write_data: std_logic_vector(31 downto 0);
  signal foo_in_pipe_write_req: std_logic_vector(0 downto 0);
  signal foo_in_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe foo_in
  signal foo_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal foo_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal foo_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe foo_out
  signal foo_out_pipe_write_data: std_logic_vector(31 downto 0);
  signal foo_out_pipe_write_req: std_logic_vector(0 downto 0);
  signal foo_out_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe foo_out
  signal foo_out_pipe_read_data: std_logic_vector(31 downto 0);
  signal foo_out_pipe_read_req: std_logic_vector(0 downto 0);
  signal foo_out_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_get
  signal free_queue_get_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_get
  signal free_queue_get_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_put
  signal free_queue_put_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_put
  signal free_queue_put_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_request
  signal free_queue_request_pipe_write_data: std_logic_vector(15 downto 0);
  signal free_queue_request_pipe_write_req: std_logic_vector(1 downto 0);
  signal free_queue_request_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe free_queue_request
  signal free_queue_request_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_data
  signal input_data_pipe_read_data: std_logic_vector(31 downto 0);
  signal input_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_data
  signal output_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal output_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module foo
  foo_instance:foo-- 
    port map(-- 
      start => foo_start,
      fin => foo_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(47 downto 32),
      memory_space_1_lr_ack => memory_space_1_lr_ack(47 downto 32),
      memory_space_1_lr_addr => memory_space_1_lr_addr(287 downto 192),
      memory_space_1_lr_tag => memory_space_1_lr_tag(143 downto 96),
      memory_space_1_lc_req => memory_space_1_lc_req(47 downto 32),
      memory_space_1_lc_ack => memory_space_1_lc_ack(47 downto 32),
      memory_space_1_lc_data => memory_space_1_lc_data(383 downto 256),
      memory_space_1_lc_tag => memory_space_1_lc_tag(143 downto 96),
      memory_space_1_sr_req => memory_space_1_sr_req(27 downto 20),
      memory_space_1_sr_ack => memory_space_1_sr_ack(27 downto 20),
      memory_space_1_sr_addr => memory_space_1_sr_addr(167 downto 120),
      memory_space_1_sr_data => memory_space_1_sr_data(223 downto 160),
      memory_space_1_sr_tag => memory_space_1_sr_tag(83 downto 60),
      memory_space_1_sc_req => memory_space_1_sc_req(27 downto 20),
      memory_space_1_sc_ack => memory_space_1_sc_ack(27 downto 20),
      memory_space_1_sc_tag => memory_space_1_sc_tag(83 downto 60),
      foo_in_pipe_read_req => foo_in_pipe_read_req(0 downto 0),
      foo_in_pipe_read_ack => foo_in_pipe_read_ack(0 downto 0),
      foo_in_pipe_read_data => foo_in_pipe_read_data(31 downto 0),
      foo_out_pipe_write_req => foo_out_pipe_write_req(0 downto 0),
      foo_out_pipe_write_ack => foo_out_pipe_write_ack(0 downto 0),
      foo_out_pipe_write_data => foo_out_pipe_write_data(31 downto 0),
      tag_in => foo_tag_in,
      tag_out => foo_tag_out-- 
    ); -- 
  -- module will be run forever 
  foo_tag_in <= (others => '0');
  foo_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => foo_start, fin => foo_fin);
  -- module free_queue_manager
  free_queue_manager_instance:free_queue_manager-- 
    port map(-- 
      start => free_queue_manager_start,
      fin => free_queue_manager_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(23 downto 12),
      memory_space_1_lr_ack => memory_space_1_lr_ack(23 downto 12),
      memory_space_1_lr_addr => memory_space_1_lr_addr(143 downto 72),
      memory_space_1_lr_tag => memory_space_1_lr_tag(71 downto 36),
      memory_space_1_lc_req => memory_space_1_lc_req(23 downto 12),
      memory_space_1_lc_ack => memory_space_1_lc_ack(23 downto 12),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 96),
      memory_space_1_lc_tag => memory_space_1_lc_tag(71 downto 36),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(1 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(3 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(15 downto 8),
      memory_space_1_sr_ack => memory_space_1_sr_ack(15 downto 8),
      memory_space_1_sr_addr => memory_space_1_sr_addr(95 downto 48),
      memory_space_1_sr_data => memory_space_1_sr_data(127 downto 64),
      memory_space_1_sr_tag => memory_space_1_sr_tag(47 downto 24),
      memory_space_1_sc_req => memory_space_1_sc_req(15 downto 8),
      memory_space_1_sc_ack => memory_space_1_sc_ack(15 downto 8),
      memory_space_1_sc_tag => memory_space_1_sc_tag(47 downto 24),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(1 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      free_queue_put_pipe_read_req => free_queue_put_pipe_read_req(0 downto 0),
      free_queue_put_pipe_read_ack => free_queue_put_pipe_read_ack(0 downto 0),
      free_queue_put_pipe_read_data => free_queue_put_pipe_read_data(31 downto 0),
      free_queue_request_pipe_read_req => free_queue_request_pipe_read_req(0 downto 0),
      free_queue_request_pipe_read_ack => free_queue_request_pipe_read_ack(0 downto 0),
      free_queue_request_pipe_read_data => free_queue_request_pipe_read_data(7 downto 0),
      free_queue_get_pipe_write_req => free_queue_get_pipe_write_req(0 downto 0),
      free_queue_get_pipe_write_ack => free_queue_get_pipe_write_ack(0 downto 0),
      free_queue_get_pipe_write_data => free_queue_get_pipe_write_data(31 downto 0),
      tag_in => free_queue_manager_tag_in,
      tag_out => free_queue_manager_tag_out-- 
    ); -- 
  -- module will be run forever 
  free_queue_manager_tag_in <= (others => '0');
  free_queue_manager_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => free_queue_manager_start, fin => free_queue_manager_fin);
  -- module input_module
  input_module_instance:input_module-- 
    port map(-- 
      start => input_module_start,
      fin => input_module_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(11 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(11 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(71 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(35 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(11 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(11 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(35 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(7 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(7 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(47 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(23 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(7 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(7 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(23 downto 0),
      free_queue_get_pipe_read_req => free_queue_get_pipe_read_req(0 downto 0),
      free_queue_get_pipe_read_ack => free_queue_get_pipe_read_ack(0 downto 0),
      free_queue_get_pipe_read_data => free_queue_get_pipe_read_data(31 downto 0),
      input_data_pipe_read_req => input_data_pipe_read_req(0 downto 0),
      input_data_pipe_read_ack => input_data_pipe_read_ack(0 downto 0),
      input_data_pipe_read_data => input_data_pipe_read_data(31 downto 0),
      foo_in_pipe_write_req => foo_in_pipe_write_req(0 downto 0),
      foo_in_pipe_write_ack => foo_in_pipe_write_ack(0 downto 0),
      foo_in_pipe_write_data => foo_in_pipe_write_data(31 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(0 downto 0),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(0 downto 0),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(7 downto 0),
      tag_in => input_module_tag_in,
      tag_out => input_module_tag_out-- 
    ); -- 
  -- module will be run forever 
  input_module_tag_in <= (others => '0');
  input_module_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => input_module_start, fin => input_module_fin);
  -- module mem_load_x_x
  mem_load_x_x_start <= '0';
  mem_load_x_x_instance:mem_load_x_x-- 
    port map(-- 
      address => mem_load_x_x_address,
      data => mem_load_x_x_data,
      start => mem_load_x_x_start,
      fin => mem_load_x_x_fin,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(7 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => mem_load_x_x_tag_in,
      tag_out => mem_load_x_x_tag_out-- 
    ); -- 
  -- module mem_store_x_x
  mem_store_x_x_start <= '0';
  mem_store_x_x_instance:mem_store_x_x-- 
    port map(-- 
      address => mem_store_x_x_address,
      data => mem_store_x_x_data,
      start => mem_store_x_x_start,
      fin => mem_store_x_x_fin,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(0 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(7 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(0 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => mem_store_x_x_tag_in,
      tag_out => mem_store_x_x_tag_out-- 
    ); -- 
  -- module output_module
  output_module_instance:output_module-- 
    port map(-- 
      start => output_module_start,
      fin => output_module_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(31 downto 24),
      memory_space_1_lr_ack => memory_space_1_lr_ack(31 downto 24),
      memory_space_1_lr_addr => memory_space_1_lr_addr(191 downto 144),
      memory_space_1_lr_tag => memory_space_1_lr_tag(95 downto 72),
      memory_space_1_lc_req => memory_space_1_lc_req(31 downto 24),
      memory_space_1_lc_ack => memory_space_1_lc_ack(31 downto 24),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(95 downto 72),
      memory_space_1_sr_req => memory_space_1_sr_req(19 downto 16),
      memory_space_1_sr_ack => memory_space_1_sr_ack(19 downto 16),
      memory_space_1_sr_addr => memory_space_1_sr_addr(119 downto 96),
      memory_space_1_sr_data => memory_space_1_sr_data(159 downto 128),
      memory_space_1_sr_tag => memory_space_1_sr_tag(59 downto 48),
      memory_space_1_sc_req => memory_space_1_sc_req(19 downto 16),
      memory_space_1_sc_ack => memory_space_1_sc_ack(19 downto 16),
      memory_space_1_sc_tag => memory_space_1_sc_tag(59 downto 48),
      foo_out_pipe_read_req => foo_out_pipe_read_req(0 downto 0),
      foo_out_pipe_read_ack => foo_out_pipe_read_ack(0 downto 0),
      foo_out_pipe_read_data => foo_out_pipe_read_data(31 downto 0),
      free_queue_put_pipe_write_req => free_queue_put_pipe_write_req(0 downto 0),
      free_queue_put_pipe_write_ack => free_queue_put_pipe_write_ack(0 downto 0),
      free_queue_put_pipe_write_data => free_queue_put_pipe_write_data(31 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(1 downto 1),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(1 downto 1),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(15 downto 8),
      output_data_pipe_write_req => output_data_pipe_write_req(0 downto 0),
      output_data_pipe_write_ack => output_data_pipe_write_ack(0 downto 0),
      output_data_pipe_write_data => output_data_pipe_write_data(31 downto 0),
      tag_in => output_module_tag_in,
      tag_out => output_module_tag_out-- 
    ); -- 
  -- module will be run forever 
  output_module_tag_in <= (others => '0');
  output_module_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => output_module_start, fin => output_module_fin);
  foo_in_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => foo_in_pipe_read_req,
      read_ack => foo_in_pipe_read_ack,
      read_data => foo_in_pipe_read_data,
      write_req => foo_in_pipe_write_req,
      write_ack => foo_in_pipe_write_ack,
      write_data => foo_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  foo_out_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => foo_out_pipe_read_req,
      read_ack => foo_out_pipe_read_ack,
      read_data => foo_out_pipe_read_data,
      write_req => foo_out_pipe_write_req,
      write_ack => foo_out_pipe_write_ack,
      write_data => foo_out_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_get_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_get_pipe_read_req,
      read_ack => free_queue_get_pipe_read_ack,
      read_data => free_queue_get_pipe_read_data,
      write_req => free_queue_get_pipe_write_req,
      write_ack => free_queue_get_pipe_write_ack,
      write_data => free_queue_get_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_put_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_put_pipe_read_req,
      read_ack => free_queue_put_pipe_read_ack,
      read_data => free_queue_put_pipe_read_data,
      write_req => free_queue_put_pipe_write_req,
      write_ack => free_queue_put_pipe_write_ack,
      write_data => free_queue_put_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_request_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_request_pipe_read_req,
      read_ack => free_queue_request_pipe_read_ack,
      read_data => free_queue_request_pipe_read_data,
      write_req => free_queue_request_pipe_write_req,
      write_ack => free_queue_request_pipe_write_ack,
      write_data => free_queue_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => input_data_pipe_read_req,
      read_ack => input_data_pipe_read_ack,
      read_data => input_data_pipe_read_data,
      write_req => input_data_pipe_write_req,
      write_ack => input_data_pipe_write_ack,
      write_data => input_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => output_data_pipe_read_req,
      read_ack => output_data_pipe_read_ack,
      read_data => output_data_pipe_read_data,
      write_req => output_data_pipe_write_req,
      write_ack => output_data_pipe_write_ack,
      write_data => output_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  RegisterBank_memory_space_0: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: memory_subsystem -- 
    generic map(-- 
      num_loads => 48,
      num_stores => 28,
      addr_width => 6,
      data_width => 8,
      tag_width => 3,
      number_of_banks => 2,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_2: register_bank -- 
    generic map(-- 
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
use work.Utility_Package.all;
use work.Vhpi_Foreign.all;
entity test_system_Test_Bench is -- 
  -- 
end entity;
architecture VhpiLink of test_system_Test_Bench is -- 
  component test_system is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      input_data_pipe_write_data: in std_logic_vector(31 downto 0);
      input_data_pipe_write_req : in std_logic_vector(0 downto 0);
      input_data_pipe_write_ack : out std_logic_vector(0 downto 0);
      output_data_pipe_read_data: out std_logic_vector(31 downto 0);
      output_data_pipe_read_req : in std_logic_vector(0 downto 0);
      output_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  signal clk: std_logic := '0';
  signal reset: std_logic := '1';
  signal foo_tag_in: std_logic_vector(0 downto 0);
  signal foo_tag_out: std_logic_vector(0 downto 0);
  signal foo_start : std_logic := '0';
  signal foo_fin   : std_logic := '0';
  signal free_queue_manager_tag_in: std_logic_vector(0 downto 0);
  signal free_queue_manager_tag_out: std_logic_vector(0 downto 0);
  signal free_queue_manager_start : std_logic := '0';
  signal free_queue_manager_fin   : std_logic := '0';
  signal input_module_tag_in: std_logic_vector(0 downto 0);
  signal input_module_tag_out: std_logic_vector(0 downto 0);
  signal input_module_start : std_logic := '0';
  signal input_module_fin   : std_logic := '0';
  signal output_module_tag_in: std_logic_vector(0 downto 0);
  signal output_module_tag_out: std_logic_vector(0 downto 0);
  signal output_module_start : std_logic := '0';
  signal output_module_fin   : std_logic := '0';
  -- write to pipe input_data
  signal input_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal input_data_pipe_write_req : std_logic_vector(0 downto 0) := (others => '0');
  signal input_data_pipe_write_ack : std_logic_vector(0 downto 0);
  -- read from pipe output_data
  signal output_data_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_data_pipe_read_req : std_logic_vector(0 downto 0) := (others => '0');
  signal output_data_pipe_read_ack : std_logic_vector(0 downto 0);
  -- 
begin --
  -- clock/reset generation 
  clk <= not clk after 5 ns;
  process
  begin --
    Vhpi_Initialize;
    wait until clk = '1';
    reset <= '0';
    while true loop --
      wait until clk = '0';
      Vhpi_Listen;
      Vhpi_Send;
      --
    end loop;
    wait;
    --
  end process;
  -- connect all the top-level modules to Vhpi
  process
  variable val_string, obj_ref: VhpiString;
  begin --
    wait until reset = '0';
    while true loop -- 
      wait until clk = '0';
      wait for 1 ns; 
      obj_ref := Pack_String_To_Vhpi_String("input_data req");
      Vhpi_Get_Port_Value(obj_ref,val_string);
      input_data_pipe_write_req <= Unpack_String(val_string,1);
      obj_ref := Pack_String_To_Vhpi_String("input_data 0");
      Vhpi_Get_Port_Value(obj_ref,val_string);
      input_data_pipe_write_data <= Unpack_String(val_string,32);
      wait until clk = '1';
      obj_ref := Pack_String_To_Vhpi_String("input_data ack");
      val_string := Pack_SLV_To_Vhpi_String(input_data_pipe_write_ack);
      Vhpi_Set_Port_Value(obj_ref,val_string);
      -- 
    end loop;
    --
  end process;
  process
  variable val_string, obj_ref: VhpiString;
  begin --
    wait until reset = '0';
    while true loop -- 
      wait until clk = '0';
      wait for 1 ns; 
      obj_ref := Pack_String_To_Vhpi_String("output_data req");
      Vhpi_Get_Port_Value(obj_ref,val_string);
      output_data_pipe_read_req <= Unpack_String(val_string,1);
      wait until clk = '1';
      obj_ref := Pack_String_To_Vhpi_String("output_data ack");
      val_string := Pack_SLV_To_Vhpi_String(output_data_pipe_read_ack);
      Vhpi_Set_Port_Value(obj_ref,val_string);
      obj_ref := Pack_String_To_Vhpi_String("output_data 0");
      val_string := Pack_SLV_To_Vhpi_String(output_data_pipe_read_data);
      Vhpi_Set_Port_Value(obj_ref,val_string);
      -- 
    end loop;
    --
  end process;
  test_system_instance: test_system -- 
    port map ( -- 
      clk => clk,
      reset => reset,
      input_data_pipe_write_data  => input_data_pipe_write_data, 
      input_data_pipe_write_req  => input_data_pipe_write_req, 
      input_data_pipe_write_ack  => input_data_pipe_write_ack,
      output_data_pipe_read_data  => output_data_pipe_read_data, 
      output_data_pipe_read_req  => output_data_pipe_read_req, 
      output_data_pipe_read_ack  => output_data_pipe_read_ack ); -- 
  -- 
end VhpiLink;
