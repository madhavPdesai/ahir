------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
package GlobalConstants is
    constant global_debug_flag: boolean := false;
    constant global_pipe_report_flag: boolean := true;
    constant global_use_vivado_bbank_dual_port : boolean := true;
    constant global_use_vivado_distributed_ram_queue : boolean := true;

    -- clock gating using Xilinx IP?
    constant use_xilinx_bufce: boolean := true;

    --
    -- for guarded statements... increase this with care!
    --
    constant max_single_bit_queue_depth_per_stage : integer := 16;  -- this is huge.. make it smaller for effect (carefully)

    -- threshold for deciding if a pipe is deep or shallow
    -- pipes shallower than this are implemented using FF's
    -- this or deeper pipes with DPRAM.  Note: this is a hack!
    constant global_pipe_shallowness_threshold : integer := 10;  


    -- use the optimized unload buffer implementation if possible.
    -- this saves a substantial amount of logic, but  can result
    -- in a slight (2.5%) performance reduction.  use it for the
    -- minimizing resource usage.
    --
    -- DANGER ALERT: do not turn this to true under any circumstances.
    --               A bug hunt is in progress.
    --
    constant global_use_optimized_unload_buffer : boolean := false;

end package GlobalConstants;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package Types is

  type ApInt is array(integer range <>) of std_logic;
  type ApIntArray is array(integer range <>, integer range <>) of std_logic;
 
  type ApFloat is array(integer range <>) of std_logic;
  type ApFloatArray is array(integer range <>, integer range <>) of std_logic;
  
  type BooleanArray is array(integer range <>) of boolean;
  type IntegerArray is array(integer range <>) of integer;
  type NaturalArray is array(integer range <>) of natural;

  type StdLogicArray2D is array (integer range <>,integer range <>) of std_logic;
  type IStdLogicVector is array (integer range <>) of std_logic; -- note: integer range

  constant slv_zero: std_logic_vector(0 downto 0) := "0";
  constant sl_zero: std_logic := '0';
  constant slv_one: std_logic_vector(0 downto 0) := "1";
  constant sl_one: std_logic := '1';

  constant loop_pipeline_buffering: integer := 4;
end package Types;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;

package Utilities is

  function Digit_To_Char(val: integer) return character;
  function Convert_To_String(val : integer) return STRING; -- convert val to string.
  function Convert_To_String(val : boolean) return STRING; -- convert val to string.
  function Convert_To_String(val : std_logic_vector) return STRING; -- convert val to string.
  function Convert_Bool_To_String(val : boolean) return STRING; -- convert bool to string.
  function Convert_SLV_To_String(val : std_logic_vector) return STRING; -- convert val to string.
  function Convert_SLV_To_Hex_String(val : std_logic_vector) return STRING; -- convert val to string.  
  function To_Hex_Char (constant val: std_logic_vector)    return character;
  
  function Ceil (constant x, y : integer)   return integer;

  function Ceil_Log2( constant x : integer)  return integer;
  function LogWidth (constant x: integer) return integer;

  function Max (constant x : NaturalArray)    return natural;
  function Sum (constant x : IntegerArray) return integer;

  function Maximum(x,y: integer)   return integer;
  function Minimum(x,y: integer)   return integer;  
  
  -- wrap around incr/decr
  function IncrWrap(x: integer; M: integer) return integer;
  function DecrWrap(x: integer; M: integer) return integer;

  function All_Entries_Same ( x : NaturalArray) return boolean;
  function Is_At_Most_One_Hot(x: BooleanArray) return Boolean;


  function Reverse(x: unsigned) return unsigned;
  procedure TruncateOrPad(signal rhs: in std_logic_vector; signal lhs : out std_logic_vector);

  function TieLowSlvConstant (constant W: integer) return std_logic_vector;
  function TieHighSlvConstant (constant W: integer) return std_logic_vector;

end Utilities;


package body Utilities is

  function Digit_To_Char(val: integer) return character is
	variable ret_val : character;
  begin
	case val is
		when 0 => ret_val := '0';
		when 1 => ret_val := '1';
		when 2 => ret_val := '2';
		when 3 => ret_val := '3';
		when 4 => ret_val := '4';
		when 5 => ret_val := '5';
		when 6 => ret_val := '6';
		when 7 => ret_val := '7';
		when 8 => ret_val := '8';
		when 9 => ret_val := '9';
		when others => ret_val := 'X';
	end case;
	return(ret_val);
  end Digit_To_Char;

    -- Thanks to: D. Calvet calvet@hep.saclay.cea.fr
    -- modified to support negative values
  function Convert_To_String(val : integer) return STRING is
	variable result : STRING(12 downto 1) := (others => '0'); -- smallest natural, longest string
	variable pos    : NATURAL := 1;
	variable tmp : integer;
	variable digit  : NATURAL;
	variable is_negative : boolean;
  begin
	tmp := val;
	if val < 0 then
	  tmp := -val;
	end if;
	is_negative := val < 0;
	
	loop
		digit := abs(tmp MOD 10);
	    	tmp := tmp / 10;
	    	result(pos) := Digit_To_Char(digit);
	    	pos := pos + 1;
	    	exit when ((tmp = 0) or (pos = (result'high-1)));
	end loop;
	
	if is_negative then
	  result(pos) := '-';
	  pos := pos + 1;
	end if;
	
	return result((pos-1) downto 1);
  end Convert_To_String;
  

  function Convert_Bool_To_String(val : boolean) return STRING is
	variable ret_var : string (1 to 5); -- convert bool to string.
  begin
    if(val) then ret_var := " true";
    else ret_var := "false"; end if;
    return(ret_var);
  end Convert_Bool_To_String;

  function Convert_To_String(val : boolean) return STRING is
	variable ret_var : string (1 to 5); -- convert bool to string.
  begin
	ret_var := Convert_Bool_To_String(val);
	return(ret_var);
  end  Convert_To_String;
   

  function Convert_SLV_To_String(val : std_logic_vector) return STRING is
	alias lval: std_logic_vector(1 to val'length) is val;
        variable ret_var: string( 1 to lval'length);
   begin
        for I in lval'range loop
                if(lval(I) = '1') then
			ret_var(I) := '1';
		elsif (lval(I) = '0') then
			ret_var(I) := '0';
		else
			ret_var(I) := 'X';
		end if;
        end loop;
        return(ret_var);
   end Convert_SLV_To_String;
    
  function Convert_To_String(val : std_logic_vector) return STRING is
	alias lval: std_logic_vector(1 to val'length) is val;
        variable ret_var: string( 1 to lval'length);
  begin
	ret_var := Convert_SLV_To_String(val);
	return(ret_var);
  end  Convert_To_String;

  function To_Hex_Char (constant val: std_logic_vector)   return character  is
    alias lval: std_logic_vector(1 to val'length) is val;
    variable tvar : std_logic_vector(1 to 4);
    variable ret_val : character;
  begin
    if(lval'length >= 4) then
      tvar := lval(1 to 4);
    else
      tvar := (others => '0');
      tvar(1 to lval'length) := lval;
    end if;

    case tvar is
      when "0000" => ret_val := '0';
      when "0001" => ret_val := '1';
      when "0010" => ret_val := '2';                     
      when "0011" => ret_val := '3';
      when "0100" => ret_val := '4';
      when "0101" => ret_val := '5';
      when "0110" => ret_val := '6';                     
      when "0111" => ret_val := '7';
      when "1000" => ret_val := '8';
      when "1001" => ret_val := '9';
      when "1010" => ret_val := 'a';                     
      when "1011" => ret_val := 'b';
      when "1100" => ret_val := 'c';
      when "1101" => ret_val := 'd';
      when "1110" => ret_val := 'e';                     
      when "1111" => ret_val := 'f';                                                               
      when others => ret_val := '?';
    end case;

    return(ret_val);
  end To_Hex_Char;
        
  function Convert_SLV_To_Hex_String(val : std_logic_vector) return STRING is
    alias lval: std_logic_vector(val'length downto 1) is val;
    variable ret_var: string( 1 to Ceil(lval'length,4));
    variable hstr  : std_logic_vector(4 downto 1);
    variable I : integer;
  begin

    I := 0;

    while I < (lval'length/4) loop
      hstr := lval(4*(I+1) downto (4*I)+1);
      ret_var(ret_var'length - I) := To_Hex_Char(hstr);
      I := (I + 1);
    end loop;  -- I

    hstr := (others => '0');
    if(ret_var'length > (lval'length/4)) then
      hstr((lval'length-((lval'length/4)*4)) downto 1) := lval(lval'length downto (4*(lval'length/4))+1);
      ret_var(1) := To_Hex_Char(hstr);
    end if;

    return(ret_var);
  end Convert_SLV_To_Hex_String;
  
  function Ceil (
    constant x, y : integer)
    return integer is
    variable ret_var : integer;
  begin
    ret_var := x/y;
    if((ret_var*y) < x) then
      ret_var := ret_var + 1;
    end if;
    return(ret_var);
  end Ceil;

  -- dont touch this?
  function Ceil_Log2
    ( constant x : integer)
    return integer is
    variable ret_var : integer;
  begin
    ret_var := 0;
    if(x > 1) then
      while((2**ret_var) < x) loop
        ret_var := ret_var + 1;
      end loop;
    end if;
    return(ret_var);
  end Ceil_Log2;

  -- x is assumed to be > 0
  function LogWidth
    ( constant x : integer)
    return integer is
    variable ret_val : integer;
    variable pow_val : integer;
  begin
    assert (x > 0) report "In LogWidth, argument must be > 0" severity error;
    ret_val := 1;

    if(x > 1) then
      while true loop
         ret_val := ret_val + 1;
         pow_val := 2**ret_val;
         if(pow_val > x) then
            exit;
         end if;
      end loop; 
    end if;

    return(ret_val);
  end LogWidth;

  function Max
    (constant x : NaturalArray)
    return natural is
    variable t, max_var : natural;
  begin
    max_var := 0;
    for I in x'low(1) to x'high(1) loop
      t := x(I);
      if( t > max_var) then
        max_var := t;
      end if;
    end loop;  -- I
    return(max_var);
  end function;

  function Sum(constant x : IntegerArray)
    return integer is
    variable ret_var : integer;
  begin
    ret_var := 0;
    for I in x'low(1) to x'high(1) loop
      ret_var := x(I) + ret_var;
    end loop;
    return(ret_var);
  end function;

  function Maximum(x,y: integer)   return integer is
    begin
      if(x > y) then
        return x;
      else
        return y;
      end if;
    end function Maximum;
    
  function Minimum(x,y: integer)   return integer is
    begin
      if(x > y) then
        return y;
      else
        return x;
      end if;
    end function Minimum;
    
  function IncrWrap(x: integer; M: integer) return integer is
    variable ret_val: integer;
  begin
    ret_val := 0;
    if(x < M) then
      ret_val := (x + 1);
    end if;
    return ret_val;
  end IncrWrap;

  function DecrWrap(x: integer; M: integer) return integer is
	variable ret_val: integer;
  begin
    ret_val := M;
    if(x > 0) then
      ret_val := (x - 1);
    end if;
    return ret_val;
  end DecrWrap;


  function All_Entries_Same ( x : NaturalArray) return boolean is
    variable ret_var : boolean;
    variable t : natural;
    alias lx : NaturalArray(x'length - 1 downto 0) is x;
  begin
    ret_var := true;
    if(lx'length > 1) then
      t := lx(lx'high);
      for I in lx'high-1 downto lx'low loop
        if(t /= lx(I)) then
          ret_var := false;
          exit;
        end if;
      end loop;  -- I
    end if;
    return(ret_var);
  end All_Entries_Same;

  function Is_At_Most_One_Hot(x: BooleanArray) return Boolean is
    variable ret_var : boolean;
    alias lx : BooleanArray(1 to x'length) is x;
    variable count : integer;
  begin
    count := 0;
    for I  in lx'range loop
      if(lx(I)) then
        count := count + 1;
      end if;
    end loop;  -- I
    if(count > 1) then
      ret_var := false;
    else
      ret_var := true;
    end if;
    return(ret_var);
  end Is_At_Most_One_Hot;


  
  function Reverse(x: unsigned) return unsigned is
	alias lx: unsigned(1 to x'length) is x;
	variable ret_var : unsigned(x'length downto 1);
  begin
	for  I in 1 to x'length loop
		ret_var(I) := lx(I);
	end loop;
	return(ret_var);
  end function Reverse;

  procedure TruncateOrPad(signal rhs: in std_logic_vector; signal lhs : out std_logic_vector) is
	alias arhs : std_logic_vector(rhs'length downto 1) is rhs;
	alias alhs : std_logic_vector(lhs'length downto 1) is lhs;
        constant L : integer := Minimum(rhs'length, lhs'length);
  begin
	alhs(L downto 1) <= arhs(L downto 1);
  end procedure TruncateOrPad;

  function TieLowSlvConstant (constant W: integer) return std_logic_vector is
	variable ret_var : std_logic_vector(1 to W) ;
  begin
	ret_var := (others => '0');
	return(ret_var);
  end TieLowSlvConstant;

  function TieHighSlvConstant (constant W: integer) return std_logic_vector is
	variable ret_var : std_logic_vector(1 to W) ;
  begin
	ret_var := (others => '1');
	return(ret_var);
  end TieHighSlvConstant;
  
end Utilities;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Utilities.all;

library aHiR_ieee_proposed;
-- use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

package Subprograms is

  function ApIntZero( l: integer) return ApInt;
  function ApFloatZero( characteristic,mantissa: integer) return ApFloat;

  function To_Boolean ( inp : ApInt) return boolean;
  function To_Boolean (  x : std_logic) return Boolean;
  function To_BooleanArray( inp: std_logic_vector) return BooleanArray;
  function To_Std_Logic ( x : boolean)   return std_logic;

  -- missing in std_logic_1164.
  function To_Std_Logic(x: bit) return std_logic;

  function To_ApInt ( inp : boolean) return ApInt;
  function To_ApInt ( inp : signed) return ApInt;
  function To_Apint ( inp : unsigned) return ApInt;
  function To_ApInt ( inp : std_logic_vector) return ApInt;
  function To_ApInt ( inp : IStdLogicVector) return ApInt;

  -- already present in float_pkg in aHiR_ieee_proposed
  --function To_Float ( x                       : std_logic_vector;
  --                    constant exponent_width : integer;
  --                    constant fraction_width : integer)
  --  return Unresolved_Float;
  
  function To_Float ( inp : ApFloat) return float;

  function To_Signed ( inp : ApInt) return signed;
  function To_Signed ( inp : std_logic_vector) return signed;
  function To_Unsigned ( inp : ApInt) return unsigned;
  function To_Unsigned ( inp : std_logic_vector) return unsigned;
  function To_Unsigned(constant W : in integer; inp : std_logic_vector) return unsigned;


  function To_SLV ( x: ApInt) return std_logic_vector;
  function To_SLV ( x: IStdLogicVector) return std_logic_vector;
  function To_SLV ( x: ApFloat) return std_logic_vector;
  function To_SLV( x : BooleanArray) return std_logic_vector;
  function To_SLV( x : Boolean) return std_logic_vector;  
  function To_SLV( x : Signed) return std_logic_vector;
  function To_SLV( x : Unsigned) return std_logic_vector;
  function Float_To_SLV( x : UNRESOLVED_float) return std_logic_vector;  
  
  function To_SLV (x : StdLogicArray2D) return std_logic_vector; 
  function To_SLV_Shuffle(x : StdLogicArray2D) return std_logic_vector;

  function To_ISLV(inp: ApInt) return IStdLogicVector;
  function To_ISLV(inp: ApFloat) return IStdLogicVector;
  function To_ISLV(inp : BooleanArray) return IStdLogicVector;
  function To_ISLV(inp : std_logic_vector) return IStdLogicVector;
  function To_ISLV(inp: Float) return IStdLogicVector;
  
  function To_StdLogicArray2D( inp: ApIntArray) return StdLogicArray2D;
  function To_StdLogicArray2D( inp: ApFloatArray) return StdLogicArray2D;
  function To_StdLogicArray2D( inp: std_logic_vector) return StdLogicArray2D;
  function To_StdLogicArray2D( inp: std_logic_vector; word_size: integer) return StdLogicArray2D;

  function To_StdLogicArray2D_Shuffle( inp: std_logic_vector; word_size: integer) return StdLogicArray2D;

  function To_ApIntArray(inp : StdLogicArray2D) return ApIntArray;
  function To_ApIntArray (inp : ApInt)   return ApIntArray;
  function To_ApIntArray (inp : integer; width : integer)   return ApIntArray;

  function To_ApFloatArray(inp : StdLogicArray2D) return ApFloatArray;
  function To_ApFloatArray (inp : ApFloat)   return ApFloatArray;

  function "&" (x : ApInt; y : ApInt) return ApInt;
  function "&" (x : ApFloat; y : ApFloat) return ApFloat;
  -- function "&" (x : std_logic_vector; y : std_logic_vector) return std_logic_vector;

  procedure Unflatten (signal z : out ApIntArray; x : in  ApInt);
  procedure Unflatten (signal z : out ApFloatArray; x : in  ApFloat);
  procedure Unflatten (signal z : out StdLogicArray2D; x : in std_logic_vector);

  function zero_pad (x : IStdLogicVector; constant h, l : integer)
    return IStdLogicVector;

  function zero_pad (x : std_logic_vector; constant h, l : integer)
    return std_logic_vector;

  function zero_pad (x : ApInt; constant h, l : integer)
    return ApInt;

  function zero_pad (x : ApFloat; constant h, l : integer)
    return ApFloat;

  function Stack( x, y : StdLogicArray2D) return StdLogicArray2D;
  procedure Split(x : in  StdLogicArray2D; y, z : out StdLogicArray2D);

  function To_ApFloat( x : float)   return ApFloat;
  function To_ApFloat( x : std_logic_vector)   return ApFloat;
  function To_ApFloat( x : std_logic_vector;  characteristic, mantissa: integer)   return ApFloat;
  function To_ApFloat( x : ApInt;  characteristic, mantissa: integer)   return ApFloat;
  function To_ApFloat ( inp : IStdLogicVector) return ApFloat;
  function To_ApFloat (x : real; characteristic, mantissa : integer) return ApFloat;
  function To_ApFloat (x : integer; characteristic, mantissa : integer) return ApFloat;

  function Extract( x : StdLogicArray2D;  idx : integer) return std_logic_vector;
  function Extract( x: ApIntArray;  idx: integer) return ApInt;
  function Extract( x: ApFloatArray;  idx: integer) return ApFloat;


  procedure Extract(source: in std_logic_vector; index: in integer; target: out std_logic_vector);
  procedure Insert(target: out std_logic_vector; index: in integer; source: in std_logic_vector);


  procedure Insert(x: out StdLogicArray2D; idx: in integer; w: in std_logic_vector );
  procedure Insert(x: out ApIntArray; idx: in integer; w: in ApInt );
  procedure Insert(x: out ApFloatArray; idx: in integer; w: in ApFloat );


  function PriorityEncode(x: BooleanArray) return BooleanArray;
  function PriorityEncode(x: std_logic_vector) return std_logic_vector;

  function OrReduce(x: BooleanArray) return boolean;
  function OrReduce(x: std_logic_vector) return std_logic;
  function OrReduce(x: unsigned) return std_logic;

  function AndReduce(x: BooleanArray) return boolean;
  function AndReduce(x: std_logic_vector) return std_logic;

  function XorReduce(x: std_logic_vector) return std_logic;

  -- generic encoders/decoders
  function GenericEncode(x: std_logic_vector) return std_logic_vector;
  function GenericDecode(x: std_logic_vector) return std_logic_vector;

  function MuxOneHot (
    constant din : StdLogicArray2D;     -- input data
    constant sel : std_logic_vector)    -- select vector (one hot)
    return std_logic_vector;

  function MuxOneHot(x: std_logic_vector; sel: BooleanArray) return std_logic_vector;
  

  function Swap_Bytes(x: std_logic_vector) return std_logic_vector;

end package Subprograms;


package body Subprograms is

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function ApIntZero( l: integer) return ApInt is
    variable ret_var : ApInt(l-1 downto 0);
  begin
    ret_var := (others => '0');
    return(ret_var);
  end ApIntZero;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function ApFloatZero( characteristic,mantissa: integer) return ApFloat is
    variable ret_var : ApFloat(characteristic downto -mantissa);
  begin
    ret_var := (others => '0');
    return(ret_var);
  end ApFloatZero;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Boolean ( inp : ApInt) return boolean is
  begin
    if(inp(inp'left) = '1') then
      return(true);
    else
      return(false);
    end if;
  end To_Boolean;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Boolean (  x : std_logic) return Boolean is
  begin
    if( x = '1') then
      return(true);
    else
      return(false);
    end if;
  end To_Boolean;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_BooleanArray( inp: std_logic_vector) return BooleanArray is
    alias linp : std_logic_vector(1 to inp'length) is inp;
    variable ret_var : BooleanArray(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := To_Boolean(linp(I));
    end loop;  -- I
    return(ret_var);
  end To_BooleanArray;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Std_Logic ( x : boolean)   return std_logic is
  begin
    if(x) then
      return('1');
    else
      return('0');
    end if;
  end To_Std_Logic;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Std_Logic(x: bit) return std_logic is
	variable ret_var : std_logic;
  begin
	if(x = '1') then 
		ret_var := '1';
	else
		ret_var := '0';
	end if;
	return(ret_var);
  end To_Std_Logic;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApInt ( inp : boolean) return ApInt is
    variable ret_var : ApInt(0 downto 0);
  begin
    if(inp) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end To_ApInt;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApInt ( inp : signed) return ApInt is
    alias linp : signed(1 to inp'length) is inp;
    variable ret_var : ApInt(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_ApInt;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Apint ( inp : unsigned) return ApInt is
    alias linp : unsigned(1 to inp'length) is inp;
    variable ret_var : ApInt(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_ApInt;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApInt ( inp : std_logic_vector) return ApInt is
    alias linp : std_logic_vector(1 to inp'length) is inp;
    variable ret_var : ApInt(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_ApInt;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApInt ( inp : IStdLogicVector) return ApInt is
    alias linp: IStdLogicVector(inp'high downto inp'low) is inp;
    variable ret_var :ApInt(inp'high downto inp'low);
  begin
    for I in linp'range loop
      ret_var(I) := linp(I);
    end loop;
    return(ret_var);
  end To_ApInt;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  --function To_Float ( x                       : std_logic_vector;
  --                    constant exponent_width : integer;
  --                    constant fraction_width : integer)
  --  return Unresolved_Float is
  --  alias lx : std_logic_vector(0 to x'length-1) is x;
  --  variable ret_var : Unresolved_Float(exponent_width downto -fraction_width);
  --begin
  --  for I in 0 to x'length loop
  --    ret_var(exponent_width-I) := lx(I);
  --  end loop;
  --  return(ret_var);
  --end To_Float;
  
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Float ( inp : ApFloat) return float is
    -- note : Apfloat is always of the form (exp downto -mantessa)
    alias linp : ApFloat(inp'high downto inp'low) is inp;
    variable ret_var : float(inp'high downto inp'low);
  begin
    for I in inp'range loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_Float;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Signed ( inp : ApInt) return signed is
    alias linp : ApInt(1 to inp'length) is inp;
    variable ret_var : signed(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_Signed;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Signed ( inp : std_logic_vector) return signed is
    alias linp : std_logic_vector(1 to inp'length) is inp;
    variable ret_var : signed(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_Signed;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Unsigned ( inp : ApInt) return unsigned is
    alias linp : ApInt(1 to inp'length) is inp;
    variable ret_var : unsigned(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_Unsigned;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Unsigned ( inp : std_logic_vector) return unsigned is
    alias linp : std_logic_vector(1 to inp'length) is inp;
    variable ret_var : unsigned(1 to inp'length);
  begin
    for I in 1 to inp'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_Unsigned;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_Unsigned(constant W : in integer; inp : std_logic_vector) return unsigned is
    alias linp : std_logic_vector(inp'length downto 1) is inp;
    variable ret_var : unsigned(Minimum(W,inp'length) downto 1);
  begin
    for I in 1 to ret_var'length loop
      ret_var(I) := linp(I);
    end loop;  -- I
    return(ret_var);
  end To_Unsigned;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV( x: ApInt) return std_logic_vector is
    alias lx: ApInt(x'length-1 downto 0) is x;
    variable rv: std_logic_vector(x'length-1 downto 0);
  begin
    for I in 1 to x'length loop
      rv(I-1) := lx(I-1);
    end loop;
    return(rv);
  end function To_SLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV( x: IStdLogicVector) return std_logic_vector is
    alias lx: IStdLogicVector(x'length-1 downto 0) is x;
    variable rv: std_logic_vector(x'length-1 downto 0);
  begin
    for I in 1 to x'length loop
      rv(I-1) := lx(I-1);
    end loop;
    return(rv);
  end function To_SLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV ( x: ApFloat) return std_logic_vector is
    alias lx: ApFloat(x'length-1 downto 0) is x;
    variable rv: std_logic_vector(x'length-1 downto 0);
  begin
    for I in 1 to x'length loop
      rv(I-1) := lx(I-1);
    end loop;
    return(rv);
  end function To_SLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV ( x: BooleanArray) return std_logic_vector is
    alias lx: BooleanArray(x'length-1 downto 0) is x;
    variable rv: std_logic_vector(x'length-1 downto 0);
  begin
    for I in 1 to x'length loop
      if(lx(I-1)) then
        rv(I-1) := '1';
      else
        rv(I-1) := '0';
      end if;
    end loop;
    return(rv);
  end function To_SLV;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV ( x: Boolean) return std_logic_vector is
    variable rv: std_logic_vector(0 downto 0);
  begin
    if(x) then
      rv(0) := '1';
    else
      rv(0) := '0';
    end if;
    return(rv);
  end function To_SLV;

  
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV ( x: Signed) return std_logic_vector is
    alias lx: Signed(1 to x'length) is x;
    variable rv: std_logic_vector(1 to x'length);
  begin
    for I in 1 to x'length loop
      rv(I) := lx(I);
    end loop;
    return(rv);
  end function To_SLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV ( x: Unsigned) return std_logic_vector is
    alias lx: Unsigned(1 to x'length) is x;
    variable rv: std_logic_vector(1 to x'length);
  begin
    for I in 1 to x'length loop
      rv(I) := lx(I);
    end loop;
    return(rv);
  end function To_SLV;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function Float_To_SLV (x: UNRESOLVED_float) return std_logic_vector is
    alias lx: UNRESOLVED_float(1 to x'length) is x;
    variable rv: std_logic_vector(1 to x'length);
  begin
    for I in 1 to x'length loop
      rv(I) := lx(I);
    end loop;
    return(rv);
  end function Float_To_SLV;
  

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ISLV(inp: ApInt) return IStdLogicVector is
    alias linp: ApInt(inp'high downto inp'low) is inp;
    variable ret_var :IStdLogicVector(inp'high downto inp'low);
  begin
    for I in linp'range loop
      ret_var(I) := linp(I);
    end loop;
    return(ret_var);
  end To_ISLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ISLV(inp: ApFloat) return IStdLogicVector is
    alias linp: ApFloat(inp'high downto inp'low) is inp;
    variable ret_var :IStdLogicVector(inp'high downto inp'low);
  begin
    for I in linp'range loop
      ret_var(I) := linp(I);
    end loop;
    return(ret_var);
  end To_ISLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ISLV(inp : BooleanArray) return IStdLogicVector is
    alias linp: BooleanArray(inp'high downto inp'low) is inp;
    variable ret_var :IStdLogicVector(inp'high downto inp'low);
  begin
    for I in linp'range loop
      ret_var(I) := To_Std_Logic(linp(I));
    end loop;
    return(ret_var);
  end To_ISLV;

    -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ISLV(inp : std_logic_vector) return IStdLogicVector is
    alias linp: std_logic_vector(inp'high downto inp'low) is inp;
    variable ret_var :IStdLogicVector(inp'high downto inp'low);
  begin
    for I in linp'range loop
      ret_var(I) := linp(I);
    end loop;
    return(ret_var);
  end To_ISLV;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ISLV(inp: Float) return IStdLogicVector is
    variable ret_var :IStdLogicVector(inp'high downto inp'low);
  begin
    for I in inp'range loop
      ret_var(I) := inp(I);
    end loop;
    return(ret_var);
  end To_ISLV;
  

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- purpose: convert a 2D array to SLV
  function To_SLV (
    x : StdLogicArray2D)
    return std_logic_vector is
    variable ret_var  : std_logic_vector((x'length(1)*x'length(2))-1 downto 0);
    variable lx : StdLogicArray2D(x'length(1)-1 downto 0, x'length(2)-1 downto 0);
  begin  -- To_SLV
    lx := x;
    for I in lx'range(1) loop
      for J in lx'range(2) loop
        ret_var((I*x'length(1))+J) := lx(I,J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end To_SLV;
  
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_SLV_Shuffle(x : StdLogicArray2D) return std_logic_vector is
    variable ret_var  : std_logic_vector((x'length(1)*x'length(2))-1 downto 0);
    variable lx : StdLogicArray2D(x'length(1)-1 downto 0, x'length(2)-1 downto 0);
    variable I : integer;
  begin
    lx := x;
    I := 0;
    while I < lx'length(1)/2 loop
      for J in lx'high(2) downto lx'low(2) loop
        ret_var((2*I*x'length(2))+J) := lx(I,J);
        ret_var((((2*I)+1)*x'length(2))+J) := lx(I+(x'length(1)/2),J);
      end loop;  -- J
      I := I + 1;
    end loop;  -- I
    return(ret_var);
  end To_SLV_Shuffle;
  
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_StdLogicArray2D( inp: ApIntArray) return StdLogicArray2D is
    variable ret_var : StdLogicArray2D(inp'range(1), inp'range(2));
  begin
    for I in ret_var'range(1) loop
      for J in ret_var'range(2) loop
        ret_var(I,J) := inp(I,J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end To_StdLogicArray2D;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_StdLogicArray2D( inp: ApFloatArray) return StdLogicArray2D is
    variable ret_var : StdLogicArray2D(inp'range(1), inp'range(2));
  begin
    for I in ret_var'range(1) loop
      for J in ret_var'range(2) loop
        ret_var(I,J) := inp(I,J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end To_StdLogicArray2D;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_StdLogicArray2D( inp: std_logic_vector) return StdLogicArray2D is
    alias linp: std_logic_vector(inp'length-1 downto 0) is inp;
    variable ret_var : StdLogicArray2D(0 downto 0, inp'length-1 downto 0);
  begin
    for I in linp'range loop
      ret_var(0,I) := linp(I);
    end loop;
    return(ret_var);
  end To_StdLogicArray2D;
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------

  function To_StdLogicArray2D( inp: std_logic_vector; word_size: integer) return StdLogicArray2D is
    variable ret_var : StdLogicArray2D((inp'length/word_size)-1 downto 0, word_size-1 downto 0);
    alias linp : std_logic_vector(inp'length-1 downto 0) is inp;
  begin
    for I in ret_var'range(1) loop
      for J in word_size-1 downto 0 loop
        ret_var(I,J) := linp((I*word_size)+J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end To_StdLogicArray2D;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  
  function To_StdLogicArray2D_Shuffle( inp: std_logic_vector; word_size: integer) return StdLogicArray2D is
    variable ret_var : StdLogicArray2D((inp'length/word_size)-1 downto 0, word_size-1 downto 0);
    alias linp : std_logic_vector(inp'length-1 downto 0) is inp;
    variable I : integer;
  begin
    I := 0;
    while I <  (ret_var'length(1)/2)-1 loop
      for J in word_size-1 downto 0 loop
        ret_var(I,J) := linp((2*I*word_size)+J);
        ret_var(I+ret_var'length(1),J) := linp((((2*I)+1)*word_size) + J);
      end loop;  -- J
      I := I + 1;
    end loop;  -- I
    return(ret_var);
  end To_StdLogicArray2D_Shuffle;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  
  function To_ApIntArray(inp : StdLogicArray2D) return ApIntArray is
    variable linp  : StdLogicArray2D(inp'high(1) downto inp'low(1), inp'high(2) downto inp'low(2));
    variable ret_var : ApIntArray(inp'high(1) downto inp'low(1), inp'high(2) downto inp'low(2));
  begin
    linp := inp;
    for I in linp'range(1) loop
      for J in linp'range(2) loop
        ret_var(I,J) := linp(I,J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end To_ApIntArray;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApIntArray (inp : ApInt)   return ApIntArray is
    variable ret_var : ApIntArray(0 downto 0, inp'range);
  begin
    for I in inp'range loop
      ret_var(0,I) := inp(I);
    end loop;  -- I
    return(ret_var);
  end To_ApIntArray;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApIntArray(inp : integer; width: integer) return ApIntArray is
  begin
    return To_ApIntArray(To_ApInt(to_signed(inp, width)));
  end To_ApIntArray;

  -----------------------------------------------------------------------------
  function To_ApFloatArray(inp : StdLogicArray2D) return ApFloatArray is
    variable linp  : StdLogicArray2D(inp'high(1) downto inp'low(1), inp'high(2) downto inp'low(2));
    variable ret_var : ApFloatArray(inp'high(1) downto inp'low(1), inp'high(2) downto inp'low(2));
  begin
    linp := inp;
    for I in linp'range(1) loop
      for J in linp'range(2) loop
        ret_var(I,J) := linp(I,J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end To_ApFloatArray;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloatArray (inp : ApFloat)   return ApFloatArray is
    variable ret_var : ApFloatArray(0 downto 0, inp'range);
  begin
    for I in inp'range loop
      ret_var(0,I) := inp(I);
    end loop;  -- I
    return(ret_var);
  end To_ApFloatArray;


  -----------------------------------------------------------------------------
  function Stack ( x, y : StdLogicArray2D) return StdLogicArray2D is
    variable lx  : StdLogicArray2D(x'length(1)-1 downto 0, x'high(2) downto x'low(2));
    variable ly  : StdLogicArray2D(y'length(1)-1 downto 0, y'high(2) downto y'low(2));
    variable ret_var:  StdLogicArray2D(x'length(1) + y'length(1) - 1 downto 0, x'high(2) downto x'low(2));
  begin
    lx := x;
    ly := y;
    assert x'high(2) = y'high(2) and x'low(2) = y'low(2) report "high/low index mismatch in Stack"
      severity error;

    for I in lx'range(1) loop
      for J  in x'high(2) downto x'low(2) loop
        ret_var(I,J) := lx(I,J);
      end loop;  -- J
    end loop;  -- I

    for I in ly'range(1) loop
      for J  in y'high(2) downto y'low(2) loop
        ret_var(I+x'length(1),J) := ly(I,J);
      end loop;  -- J
    end loop;  -- I
    return(ret_var);
  end Stack;



  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  procedure Split(x : in  StdLogicArray2D; y, z : out StdLogicArray2D) is
    variable lx  : StdLogicArray2D(x'length(1)-1 downto 0, x'high(2) downto x'low(2));
    variable ly  : StdLogicArray2D(y'length(1)-1 downto 0, y'high(2) downto y'low(2));
    variable lz  : StdLogicArray2D(z'length(1)-1 downto 0, z'high(2) downto z'low(2));
  begin
    assert x'length = (y'length + z'length) report "length mismatch in Split" severity error;
    assert x'high(2) = y'high(2) and x'high(2) = z'high(2) and x'low(2) = y'low(2) and x'low(2) = z'low(2)
      report "high/low mismatch in Split" severity error;

    lx := x;
    for I in ly'range(1) loop
      for J  in y'high(2) downto y'low(2) loop
        ly(I,J) := lx(I,J);
      end loop;  -- J
    end loop;  -- I

    for I in lz'range(1) loop
      for J  in z'high(2) downto z'low(2) loop
        lz(I,J) := lx(I+ly'length(1),J);
      end loop;  -- J
    end loop;  -- I

    y := ly;
    z := lz;
  end Procedure Split;

  -----------------------------------------------------------------------------
  -- Rearrange a really long ApInt into an ApIntArray.
  -- Used by the data-path along with the concatentation operator "&"
  -- to populate an ApIntArray using various ApInt's.
  -----------------------------------------------------------------------------
  procedure Unflatten_var (z : out StdLogicArray2D; x : in  std_logic_vector) is
    alias lx : std_logic_vector(0 to x'length - 1) is x;
    variable p : integer := 0;
  begin
    assert z'length(1) * z'length(2) = x'length
      report "z and x don't match"
      severity error;
    
    p := 0;
    
    for i in z'range(1) loop
      for j in z'range(2) loop
        z(i, j) := lx(p);
        p := p + 1;
      end loop;  -- j
    end loop;  -- i
  end procedure Unflatten_var;

  procedure Unflatten (signal z : out ApIntArray; x : in  ApInt) is
    variable lz : StdLogicArray2D(z'range(1), z'range(2));
  begin
    Unflatten_var(lz, To_SLV(x));
    z <= To_ApIntArray(lz);
  end procedure Unflatten;

  procedure Unflatten (signal z : out ApFloatArray; x : in  ApFloat) is
    variable lz : StdLogicArray2D(z'range(1), z'range(2));
  begin
    Unflatten_var(lz, To_SLV(x));
    z <= To_ApFloatArray(lz);
  end procedure Unflatten;

  procedure Unflatten (signal z : out StdLogicArray2D; x : in std_logic_vector) is
    variable lz : StdLogicArray2D(z'range(1), z'range(2));
  begin
    Unflatten_var(lz, x);
    z <= lz;
  end procedure Unflatten;
  -----------------------------------------------------------------------------
  
  -----------------------------------------------------------------------------
  -- Concatenation operator for ApInt
  -----------------------------------------------------------------------------
  --function "&" (x : std_logic_vector; y : std_logic_vector) return std_logic_vector is
    --variable z : std_logic_vector(0 to x'length + y'length - 1);
  --begin
    --z(0 to x'length - 1) := x;
    --z(x'length to z'length - 1) := y;
    --return z;
  --end function "&";

  function "&" (x : ApInt; y : ApInt) return ApInt is
  begin
    return To_ApInt(To_SLV(x) & To_SLV(y));
  end function "&";

  function "&" (x : ApFloat; y : ApFloat) return ApFloat is
  begin
    return To_ApFloat(To_SLV(x) & To_SLV(y));
  end function "&";
  -----------------------------------------------------------------------------
  
  -----------------------------------------------------------------------------
  -- pad a given value with zeroes on either side.
  -----------------------------------------------------------------------------
  function zero_pad_ascending (x : IStdLogicVector; constant h, l : integer)
    return IStdLogicVector is
    variable z : IStdLogicVector(l to h);
  begin
    assert x'ascending report "expected an SLV with ascending range" severity error;
    assert x'high <= h and x'low >= l report "input out of range" severity error;

    if z'low < x'low then
      z(z'low to x'low - 1) := (others => '0');
    end if;

    if z'high > x'high then
      z(x'high + 1 to z'high) := (others => '0');
    end if;

    z(x'low to x'high) := x;

    return z;
  end zero_pad_ascending;

  function zero_pad_descending (x : IStdLogicVector; constant h, l : integer)
    return IStdLogicVector is
    variable z : IStdLogicVector(h downto l);
  begin
    assert not x'ascending report "expected an SLV with descending range" severity error;
    assert x'high <= h and x'low >= l report "input out of range" severity error;

    if z'low < x'low then
      z(x'low - 1 downto z'low) := (others => '0');
    end if;

    if z'high > x'high then
      z(z'high downto x'high + 1) := (others => '0');
    end if;

    z(x'high downto x'low) := x;

    return z;
  end zero_pad_descending;

  function zero_pad (x : IStdLogicVector; constant h, l : integer)
    return IStdLogicVector is
  begin
    if x'ascending then
      return zero_pad_ascending(x, h, l);
    else
      return zero_pad_descending(x, h, l);
    end if;
  end zero_pad;
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- pad ApInt and ApFloat values
  -----------------------------------------------------------------------------
  function zero_pad (
    x             : ApInt;
    constant h, l : integer)
    return ApInt is
  begin
    return To_ApInt(zero_pad(To_ISLV(x), h, l));
  end zero_pad;
  
  function zero_pad (
    x             : ApFloat;
    constant h, l : integer)
    return ApFloat is
  begin
    return To_ApFloat(zero_pad(To_ISLV(x), h, l));
  end zero_pad;

  function zero_pad (
    x             : std_logic_vector;
    constant h, l : integer)
    return std_logic_vector is
  begin
    return To_SLV(zero_pad(To_ISLV(x), h, l));
  end zero_pad;
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloat( x : float)   return ApFloat is
    variable rv: ApFloat(x'high downto x'low);
  begin
    for I in x'range loop
      rv(I) := x(I);
    end loop;
    return(rv);
  end function To_ApFloat;


  -----------------------------------------------------------------------------
  function To_ApFloat( x : std_logic_vector)   return ApFloat is
    alias lx: std_logic_vector(0 to x'length-1) is x;
    variable rv: ApFloat(0 to x'length-1);
  begin
    for I in lx'range loop
      rv(I) := lx(I);
    end loop;
    return(rv);
  end function To_ApFloat;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloat( x : std_logic_vector;  characteristic, mantissa: integer)   return ApFloat is
    --alias lx: std_logic_vector(characteristic downto mantissa) is x;
    -- will not work because mantissa will be negative
    variable rv: ApFloat(characteristic downto mantissa);
    variable J: integer;
  begin
    assert (x'length = characteristic-mantissa+1)
      report "Length Mismatch in To_ApFloat" severity error;

    J := characteristic;
    for I  in x'range loop
      rv(J) := x(I);
      J := J-1;
    end loop;  -- I
    return(rv);
  end To_ApFloat;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloat( x : ApInt;  characteristic, mantissa: integer)   return ApFloat is
    alias lx: ApInt(characteristic downto mantissa) is x;
    variable rv: ApFloat(characteristic downto mantissa);
  begin
    for I  in lx'range loop
      rv(I) := lx(I);
    end loop;  -- I
    return(rv);
  end To_ApFloat;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloat ( inp : IStdLogicVector) return ApFloat is
    alias linp: IStdLogicVector(inp'high downto inp'low) is inp;
    variable ret_var :ApFloat(inp'high downto inp'low);
  begin
    for I in linp'range loop
      ret_var(I) := linp(I);
    end loop;
    return(ret_var);
  end To_ApFloat;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloat( x : real; characteristic, mantissa : integer)   return ApFloat is
  begin
    return to_apfloat(to_float(x, characteristic, mantissa));
  end function To_ApFloat;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function To_ApFloat( x : integer; characteristic, mantissa : integer)   return ApFloat is
  begin
    return to_apfloat(to_float(x, characteristic, mantissa));
  end function To_ApFloat;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function Extract( x : StdLogicArray2D;  idx : integer) return std_logic_vector is
    variable rv: IStdLogicVector(x'range(2));
  begin
    for I in x'range(2) loop
      rv(I) := x(idx,I);
    end loop;
    return To_SLV(rv);
  end function Extract;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function Extract( x: ApIntArray;  idx: integer) return ApInt is
    variable rv: ApInt(x'range(2));
  begin
    rv := To_ApInt(Extract(To_StdLogicArray2D(x),idx));
    return(rv);
  end function Extract;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function Extract( x: ApFloatArray;  idx: integer) return ApFloat is
    variable rv: ApFloat(x'range(2));
  begin
    rv := To_ApFloat(Extract(To_StdLogicArray2D(x),idx));
    return(rv);
  end function Extract;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  procedure Extract(source: in std_logic_vector; index: in integer; target: out std_logic_vector) is
  begin
    target := source(((index+1)*target'length)-1 downto (index*target'length));
  end procedure;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  procedure Insert(target: out std_logic_vector; index: in integer; source: in std_logic_vector) is
  begin
    target(((index+1)*source'length)-1 downto (index*source'length)) := source;
  end procedure;

  
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  procedure Insert(x: out StdLogicArray2D; idx: in integer; w: in std_logic_vector ) is
    alias lw: std_logic_vector(0 to w'length-1) is w;
    variable xI: integer;
  begin
    for I in lw'range loop
      if(x'ascending(2)) then
        xI := x'left(2) + I;
      else
        xI := x'left(2) - I;
      end if;
      x(idx,xI) := lw(I);
    end loop;
  end procedure Insert;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  procedure Insert(x: out ApIntArray; idx: in integer; w: in ApInt ) is
    alias lw: ApInt(0 to w'length-1) is w;
    variable xI: integer;
  begin
    for I in lw'range loop
      if(x'ascending(2)) then
        xI := x'left(2) + I;
      else
        xI := x'left(2) - I;
      end if;
      x(idx,xI) := lw(I);
    end loop;
  end procedure Insert;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  procedure Insert(x: out ApFloatArray; idx: in integer; w: in ApFloat ) is
    alias lw: ApFloat(0 to w'length-1) is w;
    variable xI: integer;
  begin
    for I in lw'range loop
      if(x'ascending(2)) then
        xI := x'left(2) + I;
      else
        xI := x'left(2) - I;
      end if;
      x(idx,xI) := lw(I);
    end loop;
  end procedure Insert;


  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function PriorityEncode(x: BooleanArray) return BooleanArray is
    alias lx  : BooleanArray(1 to x'length) is x;
    variable ret_var  : BooleanArray(1 to x'length);
  begin
    if(lx'length = 1) then
      ret_var(1) := lx(1);
    else
      ret_var := (others => false);
      if(OrReduce(lx(1 to (x'length/2)))) then
        ret_var(1 to (x'length/2)) := PriorityEncode(lx(1 to x'length/2));
      elsif(OrReduce(lx((x'length/2)+1 to x'length))) then
        ret_var((x'length/2)+1 to x'length) := PriorityEncode(lx((x'length/2)+1 to x'length));
      end if;
    end if;
    return(ret_var);
  end PriorityEncode;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function PriorityEncode(x: std_logic_vector) return std_logic_vector is
    alias lx  : std_logic_vector(1 to x'length) is x;
    variable ret_var  : std_logic_vector(1 to x'length);
  begin
    ret_var := (others => '0');
    for I in 1 to lx'length loop
       if(lx(I) = '1') then
           ret_var(I) := '1';
           exit;
       end if;
    end loop; 
    return(ret_var);
  end PriorityEncode;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function OrReduce(x: BooleanArray) return boolean is
    alias lx  : BooleanArray(1 to x'length) is x;
    variable ret_var  : Boolean;
  begin
    if(lx'length = 1) then
      ret_var := lx(1);
    else
      ret_var:= OrReduce(lx(1 to x'length/2)) or OrReduce(lx((x'length/2)+1 to x'length));
    end if;
    return(ret_var);
  end OrReduce;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function OrReduce(x: std_logic_vector) return std_logic is
	alias lx: std_logic_vector(1 to x'length) is x;
	variable ret_var: std_logic;
  begin
        ret_var := '0';	
	for I in 1 to x'length loop
		ret_var := ret_var or lx(I);
	end loop;
	return(ret_var);
  end OrReduce;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function OrReduce(x: unsigned) return std_logic is
	alias lx: unsigned(1 to x'length) is x;
	variable ret_var: std_logic;
  begin
        ret_var := '0';	
	for I in 1 to x'length loop
		ret_var := ret_var or lx(I);
	end loop;
	return(ret_var);
  end OrReduce;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function AndReduce(x: BooleanArray) return boolean is
    alias lx  : BooleanArray(1 to x'length) is x;
    variable ret_var  : Boolean;
  begin
    if(lx'length = 1) then
      ret_var := lx(1);
    else
      ret_var:= AndReduce(lx(1 to x'length/2)) and AndReduce(lx((x'length/2)+1 to x'length));
    end if;
    return(ret_var);
  end AndReduce;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function AndReduce(x: std_logic_vector) return std_logic is
  begin
    return(To_Std_Logic(AndReduce(To_BooleanArray(x))));
  end AndReduce;

  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  function XorReduce(x: std_logic_vector) return std_logic is
    alias lx  : std_logic_vector(1 to x'length) is x;
    variable ret_var  : std_logic;
  begin
    if(lx'length = 1) then
      ret_var := lx(1);
    else
      ret_var:= XorReduce(lx(1 to x'length/2)) xor XorReduce(lx((x'length/2)+1 to x'length));
    end if;
    return(ret_var);
  end XorReduce;

  -----------------------------------------------------------------------------
  -- sel is one-hot coded, build a balanced mux to
  -- pick row indicated by sel from din
  -----------------------------------------------------------------------------
  -- a utility function.
  function MuxOneHotBase (
    constant din  : StdLogicArray2D;
    constant sel  : std_logic_vector;
    constant h, l : integer)
    return std_logic_vector is
    variable ret_val : std_logic_vector(din'length(2)-1 downto 0);
    variable mid_point  : integer;
  begin
    ret_val := (others => '0');
    if(h > l) then
      mid_point := l + ((h-l)/2);
      ret_val := MuxOneHotBase(din,sel,h,mid_point+1) or
                 MuxOneHotBase(din,sel,mid_point,l);
    else
      if(sel(l) = '1') then 
      	ret_val := Extract(din,l);
      end if;
    end if;
    return(ret_val);
  end MuxOneHotBase;


  function MuxOneHot (
      constant din : StdLogicArray2D;     -- input data
      constant sel : std_logic_vector)    -- select vector (one hot)
      return std_logic_vector is
      variable ret_var : std_logic_vector(din'length(2)-1 downto 0);
      variable dinv : StdLogicArray2D(din'length(1)-1 downto 0, din'length(2)-1 downto 0);
      alias selv : std_logic_vector(sel'length-1 downto 0) is sel;
    begin
      dinv := din;
      assert sel'length = din'length(1) report "mismatched select and data dimensions" severity failure;
      ret_var := MuxOneHotBase(dinv,selv,dinv'high(1),dinv'low(1));
      return(ret_var);
    end MuxOneHot;

  function MuxOneHot(x: std_logic_vector; sel: BooleanArray) return std_logic_vector is
	variable ret_var : std_logic_vector(1 to ((x'length)/(sel'length)));
	variable mid_point : integer;
	alias lsel : BooleanArray(1 to sel'length) is sel;
	alias lx : std_logic_vector(1 to x'length) is x;
	constant word_size: integer := x'length/sel'length;
  begin
	assert( word_size*sel'length = x'length)
		report "word size not an integer" severity failure;

        if(sel'length = 1) then
		if(lsel(1)) then
            		ret_var := x;
		else
			ret_var := (others => '0');
		end if;
	else
		mid_point := sel'length/2;
		ret_var :=  MuxOneHot(lx(1 to (mid_point*word_size)), lsel(1 to mid_point)) or
                           MuxOneHot(lx((mid_point*word_size)+1 to x'length), lsel(mid_point+1 to sel'length));
	end if;
	return(ret_var);
  end MuxOneHot;
      
  function Swap_Bytes(x: std_logic_vector) return std_logic_vector is
     alias lx: std_logic_vector(1 to x'length) is x;
     variable ret_var: std_logic_vector(1 to x'length);
     variable J: integer;
     constant num_bytes: integer := (x'length/8);
  begin
     assert((x'length/8)*8 = x'length) report "Swap_Bytes argument length must be a multiple of 8" severity error;
     for I in 0 to num_bytes-1 loop
	J := (num_bytes-1) - I;
	ret_var((I*8)+1 to (I+1)*8) := lx((J*8)+1 to (J+1)*8);
     end loop;  
     return(ret_var);
  end Swap_Bytes;

  -- to be called only if x'length > 1
  function GenericEncode (x: std_logic_vector)
	return std_logic_vector is
      alias lx: std_logic_vector(x'length-1 downto 0) is x;
      variable ret_var: std_logic_vector(Ceil_Log2(x'length)-1 downto 0);
      variable TMP: unsigned(Ceil_Log2(x'length)-1 downto 0);
  begin
      ret_var := (others => '0');
      for I in 1 to x'length loop
	TMP := to_unsigned(I-1, Ceil_Log2(x'length));
        for J in 0 to Ceil_Log2(x'length)-1 loop
           if(TMP(J) = '1') then
             ret_var(J) := ret_var(J) or lx(I-1);
           end if;
        end loop;
      end loop;
      return(ret_var);
  end GenericEncode;

  function GenericDecode(x: std_logic_vector) return std_logic_vector is
     alias lx: std_logic_vector(x'length-1 downto 0) is x;
     variable ret_var: std_logic_vector((2**x'length)-1 downto 0);
     variable I : integer range 0 to (2**x'length)-1;
  begin
     ret_var := (others => '0');
     I := to_integer(to_unsigned(lx));
     ret_var(I) := '1';
     return(ret_var);
  end GenericDecode;
      
end package body Subprograms;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;                  
use aHiR_ieee_proposed.float_pkg.all;


package BaseComponents is

  -----------------------------------------------------------------------------
  -- control path components
  -----------------------------------------------------------------------------
  
  component place
    generic (
      capacity : integer := 1;
      marking : integer := 0;
      name : string);

    port (
      preds : in  BooleanArray;
      succs : in  BooleanArray;
      token : out boolean;
      clk   : in  std_logic;
      reset : in  std_logic); 
  end component;

  component place_with_bypass
    generic (
      capacity : integer := 1;
      marking : integer := 0;
      name : string );

    port (
      preds : in  BooleanArray;
      succs : in  BooleanArray;
      token : out boolean;
      clk   : in  std_logic;
      reset : in  std_logic); 
  end component;

  component transition
    generic (name: string);
    port (
      preds      : in BooleanArray;
      symbol_in  : in boolean;
      symbol_out : out boolean); 
  end component;

  component out_transition
    generic (name: string);
      port (preds      : in   BooleanArray;
              symbol_out : out  boolean);
  end component;

  component level_to_pulse 
    generic (name: string; forward_delay: integer; backward_delay: integer);
    port (clk   : in  std_logic;
          reset : in  std_logic;
          lreq: in std_logic;
          lack: out std_logic;
          preq: out boolean;
          pack: in boolean);
  end component;
  
  component control_delay_element 
    generic (name: string; delay_value: integer := 0);
    port (
      req   : in Boolean;
      ack   : out Boolean;
      clk   : in  std_logic;
      reset : in  std_logic);
  end component;

  component pipeline_interlock 
    port (name: string; trigger: in boolean;
          enable : in boolean;
          symbol_out : out  boolean;
          clk: in std_logic;
          reset: in std_logic);
  end component;

  component join is
     generic(number_of_predecessors: integer;
		place_capacity : integer := 1;
		bypass: boolean := true;
      		name : string );
     port (preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
  end component;

  component join2 
    generic (bypass : boolean := true; name: string);
    port ( pred0, pred1      : in   Boolean;
           symbol_out : out  boolean;
           clk: in std_logic;
           reset: in std_logic);
  end component;

  component generic_join2 
    generic( marking_0: integer; marking_1: integer;
		  delay_0: integer; delay_1: integer;
		    capacity_0: integer; capacity_1: integer; 
			name : string);
    port ( pred_0, pred_1      : in   Boolean;
    		symbol_out : out  boolean;
		clk: in std_logic;
		reset: in std_logic);
  end component;

  component join3 
    generic (bypass : boolean := true; name: string);
    port ( pred0, pred1, pred2      : in   Boolean;
           symbol_out : out  boolean;
           clk: in std_logic;
           reset: in std_logic);
  end component;

  component join_with_input is
     generic(number_of_predecessors: integer;
		place_capacity : integer := 1;
		bypass: boolean := false;
      		name : string );
     port (preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
    	symbol_in  : in   boolean;
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
  end component;
  
  component  generic_join 
   generic(number_of_predecessors: integer;
		name: string; place_capacities: IntegerArray; place_markings: IntegerArray; place_delays: IntegerArray);
   port ( preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
  end component;
  
  component auto_run 
    generic (use_delay : boolean);
    port (clk   : in  std_logic;
    	reset : in  std_logic;
	start_req: out std_logic;
        start_ack: in std_logic;
        fin_req: out std_logic;
        fin_ack: in std_logic);
  end component;

  component loop_terminator 
      generic (name: string; max_iterations_in_flight : integer := 4);
      port(loop_body_exit: in boolean;
       loop_continue: in boolean;
       loop_terminate: in boolean;
       loop_back: out boolean;
       loop_exit: out boolean;
       clk: in std_logic;
       reset: in std_logic);
  end component;
  

  component marked_join is
     generic(number_of_predecessors: integer;
		number_of_marked_predecessors: integer;
		place_capacity : integer := 1;
		bypass: boolean := true;
      		name : string;
		marked_predecessor_bypass: BooleanArray);
     port (preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
           marked_preds      : in   BooleanArray(number_of_marked_predecessors-1 downto 0);
           symbol_out : out  boolean;
           clk: in std_logic;
           reset: in std_logic);
  end component;

  component marked_join_with_input is
     generic(number_of_predecessors: integer;
		number_of_marked_predecessors: integer;
		place_capacity : integer := 1;
		bypass: boolean := false;
      		name : string);
     port (preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
           marked_preds      : in   BooleanArray(number_of_marked_predecessors-1 downto 0);
           symbol_in : in boolean;
           symbol_out : out  boolean;
           clk: in std_logic;
           reset: in std_logic);
  end component;

  component phi_sequencer
    generic (place_capacity: integer; nreqs : integer; nenables : integer; name : string);
    port (
      selects : in BooleanArray(0 to nreqs-1); -- one out of nreqs..
      reqs : out BooleanArray(0 to nreqs-1); -- one out of nreqs
      ack  : in Boolean;
      enables: in BooleanArray(0 to nenables-1);   -- all need to arrive to reenable
      done : out Boolean;
      clk, reset: in std_logic);
  end component;

  component phi_sequencer_v2  is
    generic (place_capacity : integer; 
	      ntriggers : integer; 
	      name : string);
    port (
  	triggers : in BooleanArray(0 to ntriggers-1); 	    -- there are nreq triggers.
  	src_sample_starts : out BooleanArray(0 to ntriggers-1);   -- sample starts for sources.
	src_sample_completes: in BooleanArray(0 to ntriggers-1);  -- sample completes from sources.
  	src_update_starts : out BooleanArray(0 to ntriggers-1);   -- update starts for sources.
	src_update_completes: in BooleanArray(0 to ntriggers-1);  -- update completes from sources.
  	phi_sample_req  : in Boolean;			   	  -- incoming sample-req to phi.
	phi_sample_ack  : out Boolean;				  -- outgoing sample-ack from phi.
  	phi_update_req  : in Boolean;			   	  -- incoming update-req to phi.
	phi_update_ack  : out Boolean;				  -- outgoing update-ack from phi.
  	phi_mux_select_reqs    : out BooleanArray(0 to ntriggers-1);	  -- phi-select mux select reqs.
	phi_mux_ack: in Boolean;				  -- ack from mux signifying select complete.
  	clk, reset: in std_logic);
   end component;

   component conditional_fork is
       generic (name: string; place_capacity: integer := 1; 
			ntriggers: integer);
       port  (triggers: in BooleanArray(0 to ntriggers-1);
			in_transition: in Boolean;
			out_transitions: out BooleanArray(0 to ntriggers-1);
			clk: in std_logic; reset: in std_logic);
   end component;

  component transition_merge 
      generic (name: string);
      port (
	   preds      : in   BooleanArray;
          symbol_out : out  boolean);
  end component;
  
  component access_regulator_base 
    generic (name : string; num_slots: integer := 1);
    port (
      -- the req-ack pair being regulated.
      req   : in Boolean;
      ack   : out Boolean;
      -- the regulated versions of req/ack
      regulated_req : out Boolean;
      regulated_ack : in Boolean;
      -- transitions on the next two will
      -- open up a slot.
      release_req   : in Boolean;
      release_ack   : in Boolean;
      clk   : in  std_logic;
      reset : in  std_logic);
  end component;

  component access_regulator 
    generic (name: string; num_reqs : integer := 1; num_slots: integer := 1; pipeline_depth: integer := 1);
    port (
      -- the req-ack pair being regulated.
      req   : in BooleanArray(num_reqs-1 downto 0);
      ack   : out BooleanArray(num_reqs-1 downto 0);
      -- the regulated versions of req/ack
      regulated_req : out BooleanArray(num_reqs-1 downto 0);
      regulated_ack : in BooleanArray(num_reqs-1 downto 0);
      -- transitions on the next two will
      -- open up a slot.
      release_req   : in BooleanArray(num_reqs-1 downto 0);
      release_ack   : in BooleanArray(num_reqs-1 downto 0);
      clk   : in  std_logic;
      reset : in  std_logic);
   end component;

  -----------------------------------------------------------------------------
  -- miscellaneous
  -----------------------------------------------------------------------------

  component RigidRepeater
    generic(name: string;
	   data_width: integer := 32);
    port(clk: in std_logic;
         reset: in std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         req_in: in std_logic;
         ack_out: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         req_out : out std_logic;
         ack_in: in std_logic);
  end component RigidRepeater;
  

  -----------------------------------------------------------------------------
  -- operator base components
  -----------------------------------------------------------------------------
  component GenericCombinationalOperator 
  generic
    (
      name: string;
	   operator_id   : string;          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer;    -- width of input2
      num_inputs    : integer := 2;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer;          -- width of output.
      constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
      constant_width: integer;
      use_constant  : boolean := false
      );
  port (
    data_in       : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
    result      : out std_logic_vector(owidth-1 downto 0)
    );
  end component GenericCombinationalOperator;

  component UnsharedOperatorBase 
    generic
      (
        name: string;
	   operator_id   : string;          -- operator id
        input1_is_int : Boolean := true; -- false means float
        input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
        input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
        iwidth_1      : integer;    -- width of input1
        input2_is_int : Boolean := true; -- false means float
        input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
        input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
        iwidth_2      : integer;    -- width of input2
        num_inputs    : integer := 2;    -- can be 1 or 2.
        output_is_int : Boolean := true;  -- false means that the output is a float
        output_characteristic_width : integer := 0;
        output_mantissa_width       : integer := 0;
        owidth        : integer;          -- width of output.
        constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
        constant_width: integer;
        use_constant  : boolean := false  -- if true, the second operand is
                                          -- assumed to be the generic
        );
    port (
      -- req -> ack follow pulse protocol
      reqL:  in Boolean;
      ackL : out Boolean;
      reqR : in Boolean;
      ackR:  out Boolean;
      -- operands.
      dataL      : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
      dataR      : out std_logic_vector(owidth-1 downto 0);
      clk, reset : in  std_logic);
  end component UnsharedOperatorBase;

  component SplitOperatorBase
    generic
      (
        name: string;
	   operator_id   : string;          -- operator id
        input1_is_int : Boolean := true; -- false means float
        input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
        input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
        iwidth_1      : integer;    -- width of input1
        input2_is_int : Boolean := true; -- false means float
        input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
        input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
        iwidth_2      : integer;    -- width of input2
        num_inputs    : integer := 2;    -- can be 1 or 2.
        output_is_int : Boolean := true;  -- false means that the output is a float
        output_characteristic_width : integer := 0;
        output_mantissa_width       : integer := 0;
        owidth        : integer;          -- width of output.
        constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
        constant_width: integer;
        twidth        : integer;          -- tag width
        use_constant  : boolean := false  -- if true, the second operand is
                                           -- provided by the generic.
        );
    port (
      -- req/ack follow level protocol
      reqR: out std_logic;
      ackR: in std_logic;
      reqL: in std_logic;
      ackL : out  std_logic;
      -- tagL is passed out to tagR
      tagL       : in  std_logic_vector(twidth-1 downto 0);
      -- input array consists of m sets of 1 or 2 possibly concatenated
      -- operands.
      dataL      : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
      dataR      : out std_logic_vector(owidth-1 downto 0);
      -- tagR is received from tagL, concurrent
      -- with dataR
      tagR       : out std_logic_vector(twidth-1 downto 0);
      clk, reset : in  std_logic);
  end component SplitOperatorBase;


  component SplitOperatorShared
    generic
      (
        name : string;
        operator_id   : string;          -- operator id
        input1_is_int : Boolean := true; -- false means float
        input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
        input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
        iwidth_1      : integer;    -- width of input1
        input2_is_int : Boolean := true; -- false means float
        input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
        input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
        iwidth_2      : integer;    -- width of input2
        num_inputs    : integer := 2;    -- can be 1 or 2.
        output_is_int : Boolean := true;  -- false means that the output is a float
        output_characteristic_width : integer := 0;
        output_mantissa_width       : integer := 0;
        owidth        : integer;          -- width of output.
        constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
        constant_width: integer;
        use_constant  : boolean := false;
        no_arbitration: boolean := false;
        min_clock_period: boolean := false;
        num_reqs : integer;  -- how many requesters?
	use_input_buffering: boolean;
        detailed_buffering_per_input: IntegerArray;
        detailed_buffering_per_output: IntegerArray;
	full_rate: boolean := false
        );

    port (
      -- req/ack follow level protocol
      reqL                     : in BooleanArray(num_reqs-1 downto 0);
      ackR                     : out BooleanArray(num_reqs-1 downto 0);
      ackL                     : out BooleanArray(num_reqs-1 downto 0);
      reqR                     : in  BooleanArray(num_reqs-1 downto 0);
      -- input data consists of concatenated pairs of ips
      dataL                    : in std_logic_vector(((iwidth_1 + iwidth_2)*num_reqs)-1 downto 0);
      -- output data consists of concatenated pairs of ops.
      dataR                    : out std_logic_vector((owidth*num_reqs)-1 downto 0);
      -- with dataR
      clk, reset              : in std_logic);
  end component SplitOperatorShared;


  component SplitOperatorSharedTB 
    generic
      ( name: string;
	   g_num_req: integer := 2;
        operator_id: string := "ApIntSle";
        verbose_mode: boolean := false;
        input_data_width: integer := 8;
        output_data_width: integer := 1;
        num_ips : integer := 2;
        tb_id : string
        );
  end component SplitOperatorSharedTB;

  -----------------------------------------------------------------------------
  -- register operator
  -----------------------------------------------------------------------------
  component RegisterBase 
      generic(name: string;
	   in_data_width: integer; out_data_width : integer);
      port(din: in std_logic_vector(in_data_width-1 downto 0);
           dout: out std_logic_vector(out_data_width-1 downto 0);
           req: in boolean;
           ack: out boolean;
           clk,reset: in std_logic);
  end component RegisterBase;

  component SynchResetRegisterSlv is
    generic(name: string; data_width: integer);
    port(din: in std_logic_vector(data_width-1 downto 0);
       dout: out std_logic_vector(data_width-1 downto 0);
       clk,reset: in std_logic);
  end component SynchResetRegisterSlv;

  component SynchResetRegisterUnsigned is
    generic(name: string; data_width: integer);
    port(din: in unsigned(data_width-1 downto 0);
       dout: out unsigned(data_width-1 downto 0);
       clk,reset: in std_logic);
  end component SynchResetRegisterUnsigned;


  -----------------------------------------------------------------------------
  -- queue, fifo, lifo
  -----------------------------------------------------------------------------
  component QueueBaseCore is
  generic(name : string := "Anon"; 
		queue_depth: integer := 3; 
		reverse_bypass_flag: boolean := false;
		data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       empty, full: out std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component QueueBaseCore;
  
  component QueueBase 
    generic(name : string; queue_depth: integer := 2; data_width: integer := 32; save_one_slot: Boolean := false);
    port(clk: in std_logic;
         reset: in std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         push_req: in std_logic;
         push_ack: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         pop_ack : out std_logic;
         pop_req: in std_logic);
  end component QueueBase;

  component QueueBaseSaveSlot
    generic(name : string; queue_depth: integer := 2; data_width: integer := 32);
    port(clk: in std_logic;
         reset: in std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         push_req: in std_logic;
         push_ack: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         pop_ack : out std_logic;
         pop_req: in std_logic);
  end component QueueBaseSaveSlot;

  component QueueWithBypass is
    generic(name : string; queue_depth: integer := 1; data_width: integer := 32);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component QueueWithBypass;

  component QueueBaseWithBypass
    generic(name : string; queue_depth: integer := 2; data_width: integer := 32);
    port(clk: in std_logic;
         reset: in std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         push_req: in std_logic;
         push_ack: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         pop_ack : out std_logic;
         pop_req: in std_logic);
  end component QueueBaseWithBypass;

  component QueueBaseWithEmptyFull
    generic(name : string; queue_depth: integer := 2; reverse_bypass_flag: boolean := false; data_width: integer := 32);
    port(clk: in std_logic;
         reset: in std_logic;
         empty, full: out std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         push_req: in std_logic;
         push_ack: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         pop_ack : out std_logic;
         pop_req: in std_logic);
  end component QueueBaseWithEmptyFull;

  component QueueEmptyFullLogic is
	port (clk, reset: in std_logic;
		read,write,eq_flag: in boolean;
		full, empty: out boolean);
  end component;


  --
  -- a special purpose queue which keeps a 1-bit data value.
  --
  component SingleBitQueueBase is
    generic(name : string; queue_depth: integer := 1; bypass_flag: boolean := false);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(0 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(0 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component SingleBitQueueBase;

  component SynchFifoWithDPRAM
    generic(name: string; queue_depth: integer := 3; data_width: integer := 72);
    port(clk: in std_logic;
         reset: in std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         push_req: in std_logic;
         push_ack : out std_logic;
         nearly_full: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         pop_ack : out std_logic;
         pop_req: in std_logic);
  end component SynchFifoWithDPRAM;

  component SynchLifo 
    generic(name : string; queue_depth: integer := 3; data_width: integer := 72);
    port(clk: in std_logic;
         reset: in std_logic;
         data_in: in std_logic_vector(data_width-1 downto 0);
         push_req: in std_logic;
         push_ack : out std_logic;
         nearly_full: out std_logic;
         data_out: out std_logic_vector(data_width-1 downto 0);
         pop_ack : out std_logic;
         pop_req: in std_logic);
  end component SynchLifo;
  
  component SynchToAsynchReadInterface 
    generic (
      name: string;
      data_width : integer);
    port (
      clk : in std_logic;
      reset  : in std_logic;
      synch_req : in std_logic;
      synch_ack : out std_logic;
      asynch_req : out std_logic;
      asynch_ack: in std_logic;
      synch_data: in std_logic_vector(data_width-1 downto 0);
      asynch_data : out std_logic_vector(data_width-1 downto 0));
    
  end component SynchToAsynchReadInterface;

  component ShiftRegisterQueue is
    generic(name : string ; queue_depth: integer := 1; data_width: integer := 32);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component;


  component ShiftRegisterSingleBitQueue is
    generic(name : string; queue_depth: integer; number_of_stages: integer; bypass_flag: boolean := false);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(0 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(0 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component ShiftRegisterSingleBitQueue;

  -----------------------------------------------------------------------------
  -- pipe
  -----------------------------------------------------------------------------
  component PipeBase 
    
    generic (name : string;
	     num_reads: integer;
             num_writes: integer;
             data_width: integer;
             lifo_mode: boolean := false;
             depth: integer := 1;
	     signal_mode: boolean := false;
 	     shift_register_mode: boolean := false;
	     save_slot: boolean := false;
	     bypass: boolean := false;
	     full_rate : boolean := false);
    port (
      read_req       : in  std_logic_vector(num_reads-1 downto 0);
      read_ack       : out std_logic_vector(num_reads-1 downto 0);
      read_data      : out std_logic_vector((num_reads*data_width)-1 downto 0);
      write_req       : in  std_logic_vector(num_writes-1 downto 0);
      write_ack       : out std_logic_vector(num_writes-1 downto 0);
      write_data      : in std_logic_vector((num_writes*data_width)-1 downto 0);
      clk, reset : in  std_logic);
    
  end component PipeBase;

  component PipelineRegister is
  generic (name : string;
           data_width: integer);
  port (
    read_req       : in  std_logic;
    read_ack       : out std_logic;
    read_data      : out std_logic_vector(data_width-1 downto 0);
    write_req       : in  std_logic;
    write_ack       : out std_logic;
    write_data      : in std_logic_vector((data_width-1) downto 0);
    clk, reset : in  std_logic);
   end component PipelineRegister;

  -----------------------------------------------------------------------------
  -- phi,branch,select
  -----------------------------------------------------------------------------

  component PhiBase 
    generic (
      name: string;
      num_reqs   : integer;
      data_width : integer;
      bypass_flag: boolean := false);
    port (
      req                 : in  BooleanArray(num_reqs-1 downto 0);
      ack                 : out Boolean;
      idata               : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
      odata               : out std_logic_vector(data_width-1 downto 0);
      clk, reset          : in std_logic);
  end component PhiBase;

  
  component PhiPipelined is
    generic (
      name       : string;
      num_reqs   : integer;
      buffering  : integer;
      data_width : integer);
    port (
      sample_req                 : in  BooleanArray(num_reqs-1 downto 0);
      sample_ack                 : out Boolean;
      update_req                 : in Boolean;
      update_ack                 : out Boolean;
      idata                      : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
      odata                      : out std_logic_vector(data_width-1 downto 0);
      clk, reset                 : in std_logic);
  end component;


  component BranchBase
    generic (
      name: string;
      condition_width : integer;
      bypass_flag: boolean := false);
    port (condition: in std_logic_vector(condition_width-1 downto 0);
          clk,reset: in std_logic;
          req: in Boolean;
          ack0: out Boolean;
          ack1: out Boolean);
  end component;

  component SelectBase 
    generic(name: string; data_width: integer; flow_through: boolean := false);
    port(x,y: in std_logic_vector(data_width-1 downto 0);
         sel: in std_logic_vector(0 downto 0);
         req: in boolean;
         z: out std_logic_vector(data_width-1 downto 0);
         ack: out boolean;
         clk,reset: in std_logic);
  end component SelectBase;

  component Slicebase 
    generic(name: string; in_data_width : integer; high_index: integer; low_index : integer; flow_through : boolean := false);
    port(din: in std_logic_vector(in_data_width-1 downto 0);
         dout: out std_logic_vector(high_index-low_index downto 0);
         req: in boolean;
         ack: out boolean;
         clk,reset: in std_logic);
  end component Slicebase;

  component SliceSplitProtocol is
    generic(name: string; 
	in_data_width : integer; 
	high_index: integer; 
	low_index : integer; 
	buffering : integer;
	flow_through: boolean := false; 
	full_rate: boolean := false
	);
    port(din: in std_logic_vector(in_data_width-1 downto 0);
       dout: out std_logic_vector(high_index-low_index downto 0);
       sample_req: in boolean;
       sample_ack: out boolean;
       update_req: in boolean;
       update_ack: out boolean;
       clk,reset: in std_logic);
  end component;

  -----------------------------------------------------------------------------
  -- mux/demux
  -----------------------------------------------------------------------------
  
  component InputMuxBase 
    generic ( name: string; iwidth: integer;
              owidth: integer;
              twidth: integer;
              nreqs: integer;
              no_arbitration: Boolean;
              registered_output: Boolean);
    port (
      -- req/ack follow pulse protocol
      reqL                 : in  BooleanArray(nreqs-1 downto 0);
      ackL                 : out BooleanArray(nreqs-1 downto 0);
      dataL                : in  std_logic_vector(iwidth-1 downto 0);
      -- output side req/ack level protocol
      reqR                 : out std_logic;
      ackR                 : in  std_logic;
      dataR                : out std_logic_vector(owidth-1 downto 0);
      -- tag specifies the requester index 
      tagR                : out std_logic_vector(twidth-1 downto 0);
      clk, reset          : in std_logic);
  end component InputMuxBase;

  component InputMuxBaseNoData 
    generic ( name: string; twidth: integer;
              nreqs: integer;
              no_arbitration: Boolean);
    port (
      -- req/ack follow pulse protocol
      reqL                 : in  BooleanArray(nreqs-1 downto 0);
      ackL                 : out BooleanArray(nreqs-1 downto 0);
      -- output side req/ack level protocol
      reqR                 : out std_logic;
      ackR                 : in  std_logic;
      -- tag specifies the requester index 
      tagR                : out std_logic_vector(twidth-1 downto 0);
      clk, reset          : in std_logic);
  end component InputMuxBaseNoData;



  component OutputDeMuxBaseNoData
    generic(name : string;
	    twidth: integer;
            nreqs: integer;
	    detailed_buffering_per_output: IntegerArray);
    port (
      -- req/ack follow level protocol
      reqL                 : in  std_logic;
      ackL                 : out std_logic;
      -- tag identifies index to which demux
      -- should happen
      tagL                 : in std_logic_vector(twidth-1 downto 0);
      -- reqR/ackR follow pulse protocol
      -- and are of length n
      reqR                : in BooleanArray(nreqs-1 downto 0);
      ackR                : out  BooleanArray(nreqs-1 downto 0);
      clk, reset          : in std_logic);
  end component OutputDeMuxBaseNoData;

  component OutputDeMuxBase
    generic(name: string; iwidth: integer;
            owidth: integer;
            twidth: integer;
            nreqs: integer;
            no_arbitration: Boolean;
            pipeline_flag : Boolean := true);
    port (
      -- req/ack follow level protocol
      reqL                 : in  std_logic;
      ackL                 : out std_logic;
      dataL                : in  std_logic_vector(iwidth-1 downto 0);
      -- tag identifies index to which demux
      -- should happen
      tagL                 : in std_logic_vector(twidth-1 downto 0);
      -- reqR/ackR follow pulse protocol
      -- and are of length n
      reqR                : in BooleanArray(nreqs-1 downto 0);
      ackR                : out  BooleanArray(nreqs-1 downto 0);
      -- dataR is array(n,m) 
      dataR               : out std_logic_vector(owidth-1 downto 0);
      clk, reset          : in std_logic);
  end component OutputDeMuxBase;
  

  component OutputDeMuxBaseWithBuffering
    generic(name : string;
            iwidth: integer;
            owidth: integer;
            twidth: integer;
            nreqs : integer;
            detailed_buffering_per_output: IntegerArray;
	    full_rate : boolean);
    port (
      -- req/ack follow level protocol
      reqL                 : in  std_logic;
      ackL                 : out std_logic;
      dataL                : in  std_logic_vector(iwidth-1 downto 0);
      -- tag identifies index to which demux
      -- should happen
      tagL                 : in std_logic_vector(twidth-1 downto 0);
      -- reqR/ackR follow pulse protocol
      -- and are of length n
      reqR                : in BooleanArray(nreqs-1 downto 0);
      ackR                : out  BooleanArray(nreqs-1 downto 0);
      -- dataR is array(n,m) 
      dataR               : out std_logic_vector(owidth-1 downto 0);
      clk, reset          : in std_logic);
  end component OutputDeMuxBaseWithBuffering;
  

  -----------------------------------------------------------------------------
  -- call arbiters
  -- there are four forms for the four possibilities of the
  -- called function (in-args+out-args, in-args, out-args, no args)
  -----------------------------------------------------------------------------
  component CallArbiter
    generic(name: string; num_reqs: integer;
            call_data_width: integer;
            return_data_width: integer;
            tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
      -- call port connected to the called module
      call_mreq   : out std_logic;
      call_mack   : in  std_logic;
      call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
      call_mtag   : out std_logic_vector(tag_length-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks : out std_logic_vector(num_reqs-1 downto 0);
      return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
      -- return from function
      -- function to assert mreq arbiter to return mack
      -- ( NOTE: It has to be this way, the arbiter should
      -- accept the return value if it has room)
      return_mreq : in std_logic;
      return_mack : out std_logic;
      return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
      return_mtag : in  std_logic_vector(tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiter;

  component CallArbiterNoInargs
    generic(name: string; num_reqs: integer;
            return_data_width: integer;
            tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      -- call port connected to the called module
      call_mreq   : out std_logic;
      call_mack   : in  std_logic;
      call_mtag   : out std_logic_vector(tag_length-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks : out std_logic_vector(num_reqs-1 downto 0);
      return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
      -- return from function
      -- function to assert mreq arbiter to return mack
      -- ( NOTE: It has to be this way, the arbiter should
      -- accept the return value if it has room)
      return_mreq : in std_logic;
      return_mack : out std_logic;
      return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
      return_mtag : in  std_logic_vector(tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterNoInargs;

  component CallArbiterNoOutargs
    generic(name: string; num_reqs: integer;
            call_data_width: integer;
            tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
      -- call port connected to the called module
      call_mreq   : out std_logic;
      call_mack   : in  std_logic;
      call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
      call_mtag   : out std_logic_vector(tag_length-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks : out std_logic_vector(num_reqs-1 downto 0);
      -- return from function
      -- function to assert mreq arbiter to return mack
      -- ( NOTE: It has to be this way, the arbiter should
      -- accept the return value if it has room)
      return_mreq : in std_logic;
      return_mack : out std_logic;
      return_mtag : in  std_logic_vector(tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterNoOutargs;



  component CallArbiterNoInargsNoOutargs
    generic(name: string; num_reqs: integer;
            tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      -- call port connected to the called module
      call_mreq   : out std_logic;
      call_mack   : in  std_logic;
      call_mtag   : out std_logic_vector(tag_length-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks : out std_logic_vector(num_reqs-1 downto 0);
      -- return from function
      -- function to assert mreq arbiter to return mack
      -- ( NOTE: It has to be this way, the arbiter should
      -- accept the return value if it has room)
      return_mreq : in std_logic;
      return_mack : out std_logic;
      return_mtag : in  std_logic_vector(tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterNoInargsNoOutargs;


  component CallArbiterUnitary
    generic(name: string; num_reqs: integer;
            call_data_width: integer;
            return_data_width: integer;
            caller_tag_length: integer;
            callee_tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
      call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks   : out std_logic_vector(num_reqs-1 downto 0);
      return_data   : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
      return_tag    : out  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- ports connected to the called module
      call_start   : out std_logic;
      call_fin   : in  std_logic;
      call_in_args  : out std_logic_vector(call_data_width-1 downto 0);
      call_in_tag   : out std_logic_vector(callee_tag_length-1 downto 0);
      -- from the called module
      call_out_args : in  std_logic_vector(return_data_width-1 downto 0);
      call_out_tag : in  std_logic_vector(callee_tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterUnitary;


  component CallArbiterUnitaryNoInargs
    generic(name: string; num_reqs: integer;
            return_data_width: integer;
            caller_tag_length: integer;
            callee_tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks   : out std_logic_vector(num_reqs-1 downto 0);
      return_data   : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
      return_tag    : out  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- ports connected to the called module
      call_start   : out std_logic;
      call_fin   : in  std_logic;
      call_in_tag   : out std_logic_vector(callee_tag_length-1 downto 0);
      -- from the called module
      call_out_args : in  std_logic_vector(return_data_width-1 downto 0);
      call_out_tag : in  std_logic_vector(callee_tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterUnitaryNoInargs;

  component CallArbiterUnitaryNoOutargs
    generic(name: string; num_reqs: integer;
            call_data_width: integer;
            caller_tag_length: integer;
            callee_tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
      call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks   : out std_logic_vector(num_reqs-1 downto 0);
      return_tag    : out  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- ports connected to the called module
      call_start   : out std_logic;
      call_fin   : in  std_logic;
      call_in_args  : out std_logic_vector(call_data_width-1 downto 0);
      call_in_tag   : out std_logic_vector(callee_tag_length-1 downto 0);
      -- from the called module
      call_out_tag : in  std_logic_vector(callee_tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterUnitaryNoOutargs;


  component CallArbiterUnitaryNoInargsNoOutargs
    generic(name: string; num_reqs: integer;
            caller_tag_length: integer;
            callee_tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks   : out std_logic_vector(num_reqs-1 downto 0);
      return_tag    : out  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- ports connected to the called module
      call_start   : out std_logic;
      call_fin   : in  std_logic;
      call_in_tag   : out std_logic_vector(callee_tag_length-1 downto 0);
      -- from the called module
      call_out_tag : in  std_logic_vector(callee_tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component CallArbiterUnitaryNoInargsNoOutargs;

  component CallMediator
    port (
      call_req: in std_logic;
      call_ack: out std_logic;
      enable_call_data: out std_logic;
      return_req: in std_logic;
      return_ack: out std_logic;
      enable_return_data: out std_logic;
      start: out std_logic;
      fin: in std_logic;
      clk: in std_logic;
      reset: in std_logic);
  end component CallMediator;

  -----------------------------------------------------------------------------
  --   NobodyLeftBehind..
  --   this is a small utility which ensures that there is no starvation
  --   in the system.. needs to be used as a filter between reqs and priority
  --   encoding.  currently used in split-call arbiters.
  -----------------------------------------------------------------------------
  component  NobodyLeftBehind 
     generic (name: string;  num_reqs : integer := 1);
     port (
       clk,reset : in std_logic;
       reqIn : in std_logic_vector(num_reqs-1 downto 0);
       ackOut: out std_logic_vector(num_reqs-1 downto 0);
       reqOut : out std_logic_vector(num_reqs-1 downto 0);
       ackIn : in std_logic_vector(num_reqs-1 downto 0));
  end component;

  -----------------------------------------------------------------------------
  -- split call arbiters..
  --   Modules will now have a split request-complete handshake
  --   (just like operators)
  -----------------------------------------------------------------------------
  component SplitCallArbiter
    generic(name: string; num_reqs: integer;
	  call_data_width: integer;
	  return_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
      call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- call port connected to the called module
      call_mreq   : out std_logic;
      call_mack   : in  std_logic;
      call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
      call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks : out std_logic_vector(num_reqs-1 downto 0);
      return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
      return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- return from function
      return_mreq : out std_logic;
      return_mack : in std_logic;
      return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
      return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component SplitCallArbiter;

  component SplitCallArbiterNoInargs
  generic(name: string; num_reqs: integer;
	  return_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
  end component SplitCallArbiterNoInargs;

  component SplitCallArbiterNoOutargs
    generic(name: string; num_reqs: integer;
	  call_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
  end component SplitCallArbiterNoOutargs;



  component SplitCallArbiterNoInargsNoOutargs
    generic(name: string; num_reqs: integer;
            caller_tag_length: integer;
            callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
  end component SplitCallArbiterNoInargsNoOutargs;


  -----------------------------------------------------------------------------
  -- IO ports
  -----------------------------------------------------------------------------
  component InputPort
    generic (name: string; num_reqs: integer;
             data_width: integer;
             no_arbitration: boolean);
    port (
      -- pulse interface with the data-path
      req        : in  BooleanArray(num_reqs-1 downto 0);
      ack        : out BooleanArray(num_reqs-1 downto 0);
      data       : out std_logic_vector((num_reqs*data_width)-1 downto 0);
      -- ready/ready interface with outside world
      oreq       : out std_logic;
      oack       : in  std_logic;
      odata      : in  std_logic_vector(data_width-1 downto 0);
      clk, reset : in  std_logic);
  end component;

  component InputPortNoData
    generic (name: string; num_reqs: integer;
             no_arbitration: boolean);
    port (
      -- pulse interface with the data-path
      req        : in  BooleanArray(num_reqs-1 downto 0);
      ack        : out BooleanArray(num_reqs-1 downto 0);
      -- ready/ready interface with outside world
      oreq       : out std_logic;
      oack       : in  std_logic;
      clk, reset : in  std_logic);
  end component;


  component InputPortLevel
    generic (name: string; num_reqs: integer; 
             data_width: integer;  
             no_arbitration: boolean);
    port (
      -- ready/ready interface with the requesters
      req       : in  std_logic_vector(num_reqs-1 downto 0);
      ack       : out std_logic_vector(num_reqs-1 downto 0);
      data      : out std_logic_vector((num_reqs*data_width)-1 downto 0);
      -- ready/ready interface with outside world
      oreq       : out std_logic;
      oack       : in  std_logic;
      odata      : in  std_logic_vector(data_width-1 downto 0);
      clk, reset : in  std_logic);
  end component InputPortLevel;


  component InputPortLevelNoData 
    generic (name: string; num_reqs: integer; 
             no_arbitration: boolean);
    port (
      -- ready/ready interface with the requesters
      req       : in  std_logic_vector(num_reqs-1 downto 0);
      ack       : out std_logic_vector(num_reqs-1 downto 0);
      -- ready/ready interface with outside world
      oreq       : out std_logic;
      oack       : in  std_logic;
      clk, reset : in  std_logic);
  end component;

  component InputPortSingleReader is
  generic (name : string;
	   data_width: integer);
  port (
    -- pulse interface with the data-path
    sample_req        : in  BooleanArray(0 downto 0); -- sacrificial.
    sample_ack        : out BooleanArray(0 downto 0); -- sacrificial.
    update_req        : in  BooleanArray(0 downto 0);
    update_ack        : out BooleanArray(0 downto 0);
    data              : out std_logic_vector((data_width-1) downto 0);
    -- ready/ready interface with outside world
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : in  std_logic_vector((data_width-1) downto 0);
    clk, reset : in  std_logic);
  end component;

  component OutputPort
    generic(name: string; num_reqs: integer;
            data_width: integer;
            no_arbitration: boolean);
    port (
      req        : in  BooleanArray(num_reqs-1 downto 0);
      ack        : out BooleanArray(num_reqs-1 downto 0);
      data       : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
      oreq       : out std_logic;
      oack       : in  std_logic;
      odata      : out std_logic_vector(data_width-1 downto 0);
      clk, reset : in  std_logic);
  end component;


  component OutputPortNoData
    generic(name: string; num_reqs: integer;
            no_arbitration: boolean);
    port (
      req        : in  BooleanArray(num_reqs-1 downto 0);
      ack        : out BooleanArray(num_reqs-1 downto 0);
      oreq       : out std_logic;
      oack       : in  std_logic;
      clk, reset : in  std_logic);
  end component;
  
  component OutputPortLevel
    generic(name: string; num_reqs: integer;
            data_width: integer;
            no_arbitration: boolean);
    port (
      req       : in  std_logic_vector(num_reqs-1 downto 0);
      ack       : out std_logic_vector(num_reqs-1 downto 0);
      data      : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
      oreq       : out std_logic;
      oack       : in  std_logic;
      odata      : out std_logic_vector(data_width-1 downto 0);
      clk, reset : in  std_logic);
  end component;

  component OutputPortLevelNoData 
    generic(name: string; num_reqs: integer;
            no_arbitration: boolean);
    port (
      req       : in  std_logic_vector(num_reqs-1 downto 0);
      ack       : out std_logic_vector(num_reqs-1 downto 0);
      oreq       : out std_logic;
      oack       : in  std_logic;
      clk, reset : in  std_logic);
  end component;

  component OutputPortSingleWriter is
  generic(name : string;
	  data_width: integer);
  port (
    sample_req        : in  BooleanArray(0 downto 0);
    sample_ack        : out BooleanArray(0 downto 0);
    update_req        : in  BooleanArray(0 downto 0); -- sacrificial
    update_ack        : out BooleanArray(0 downto 0); -- sacrificial
    data       : in  std_logic_vector((data_width-1) downto 0);
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : out std_logic_vector((data_width-1) downto 0);
    clk, reset : in  std_logic);
  end component;
  -----------------------------------------------------------------------------
  -- load/store
  -----------------------------------------------------------------------------
  component LoadReqShared
    generic
      (
	name: string; 	addr_width: integer;
      	num_reqs : integer; -- how many requesters?
	tag_length: integer;
	no_arbitration: Boolean;
	time_stamp_width: integer;
        min_clock_period: Boolean
        );
    port (
      -- req/ack follow pulse protocol
      reqL                     : in BooleanArray(num_reqs-1 downto 0);
      ackL                     : out BooleanArray(num_reqs-1 downto 0);
      -- concatenated address corresponding to access
      dataL                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
      -- address to memory
      maddr                   : out std_logic_vector(addr_width-1 downto 0);
      mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);
      mreq                    : out std_logic;
      mack                    : in std_logic;
      -- clock, reset (active high)
      clk, reset              : in std_logic);
  end component LoadReqShared;

  component StoreReqShared
    generic
      (
	name: string;
	addr_width: integer;
	data_width : integer;
	time_stamp_width: integer;
      	num_reqs : integer; -- how many requesters?
	tag_length: integer;
        min_clock_period : boolean;
	no_arbitration: Boolean
        );
    port (
      -- req/ack follow pulse protocol
      reqL                     : in BooleanArray(num_reqs-1 downto 0);
      ackL                     : out BooleanArray(num_reqs-1 downto 0);
      -- address corresponding to access
      addr                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
      data                    : in std_logic_vector((data_width*num_reqs)-1 downto 0);
      -- address to memory
      maddr                   : out std_logic_vector(addr_width-1 downto 0);
      mdata                   : out std_logic_vector(data_width-1 downto 0);
      mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);
      mreq                    : out std_logic;
      mack                    : in std_logic;
      -- clock, reset (active high)
      clk, reset              : in std_logic);
  end component StoreReqShared;


  component LoadCompleteShared
    generic
      (
        name : string;
        data_width: integer;
        tag_length:  integer;
        num_reqs : integer;
        no_arbitration: boolean;
        detailed_buffering_per_output : IntegerArray
        );
    port (
      -- req/ack follow level protocol
      reqR                     : in BooleanArray(num_reqs-1 downto 0);
      ackR                     : out BooleanArray(num_reqs-1 downto 0);
      dataR                    : out std_logic_vector((data_width*num_reqs)-1 downto 0);
      -- output data consists of concatenated pairs of ops.
      mdata                    : in std_logic_vector(data_width-1 downto 0);
      mreq                     : out std_logic;
      mack                     : in  std_logic;
      mtag                     : in std_logic_vector(tag_length-1 downto 0);
      -- with dataR
      clk, reset              : in std_logic);
  end component LoadCompleteShared;

  component StoreCompleteShared
    generic (name: string; 
	     num_reqs: integer;
             tag_length: integer;
	     detailed_buffering_per_output: IntegerArray);
    port (
      -- in requester array, pulse protocol
      -- more than one requester can be active
      -- at any time
      reqR : in BooleanArray(num_reqs-1 downto 0);
      -- out ack array, pulse protocol
      -- more than one ack can be sent back
      -- at any time.
      --
      -- Note: req -> ack delay can be 0
      ackR : out BooleanArray(num_reqs-1 downto 0);
      -- mreq goes out to memory as 
      -- a response to mack.
      mreq : out std_logic;
      mack : in  std_logic;
      -- mtag to distinguish the 
      -- requesters.
      mtag : in std_logic_vector(tag_length-1 downto 0);
      -- rising edge of clock is used
      clk : in std_logic;
      -- synchronous reset, active high
      reset : in std_logic);
  end component StoreCompleteShared;


  -----------------------------------------------------------------------------
  -- protocol translation, priority encoding
  -----------------------------------------------------------------------------
  component Pulse_To_Level_Translate_Entity 
    generic (name: string);
    port( rL : in boolean;
          rR : out std_logic;
          aL : out boolean;
          aR : in std_logic;
          clk : in std_logic;
          reset : in std_logic);
  end component;

  component Stall_To_Pulse_Translate_Entity is
    generic (name : string);
    port(
	stall_out : out std_logic;
        rR : in  boolean;
        valid_in : in std_logic;
        aR : out boolean;
        clk : in std_logic;
        reset : in std_logic);
  end component;

  component Sample_Pulse_To_Level_Translate_Entity 
    generic (name: string);
    port( rL : in boolean;
          rR : out std_logic;
          aL : out boolean;
          aR : in std_logic;
          clk : in std_logic;
          reset : in std_logic);
  end component;

  component Level_To_Pulse_Translate_Entity is
    generic (name: string);
    port( rL : out std_logic;
        rR : in  boolean;
        aL : in std_logic;
        aR : out boolean;
        clk : in std_logic;
        reset : in std_logic);
  end component;

  component Request_Priority_Encode_Entity
    generic (name:string; num_reqs : integer := 1);
    port (
      clk,reset : in std_logic;
      reqR : in std_logic_vector;
      ackR: out std_logic_vector;
      forward_enable: out std_logic_vector;
      req_s : out std_logic;
      ack_s : in std_logic);
  end component;

  -----------------------------------------------------------------------------
  -- BinaryEncoder: introduced because Xilinx ISE 13.1 barfs on To_Unsigned
  -----------------------------------------------------------------------------
  component BinaryEncoder
    generic (name: string; iwidth: integer := 3; owidth: integer := 3);
    port(din: in std_logic_vector(iwidth-1 downto 0);
         dout: out std_logic_vector(owidth-1 downto 0));
  end component;


  -----------------------------------------------------------------------------
  -- floating point operators (pipelined)
  -----------------------------------------------------------------------------
  
  component GenericFloatToFloat is
    generic (name: string;
	   tag_width : integer;
           in_exponent_width: integer;
           in_fraction_width : integer;
           out_exponent_width: integer;
           out_fraction_width : integer;
           round_style : round_type := float_round_style;  -- rounding option
           addguard       : NATURAL := float_guard_bits;  -- number of guard bits
           check_error : BOOLEAN    := float_check_error;  -- check for errors
           denormalize_in : BOOLEAN := float_denormalize;  -- Use IEEE extended FP           
           denormalize : BOOLEAN    := float_denormalize  -- Use IEEE extended FP           
           );
    port(
      INF: in std_logic_vector((in_exponent_width+in_fraction_width) downto 0);
      OUTF: out std_logic_vector((out_exponent_width+out_fraction_width) downto 0);
      clk,reset: in std_logic;
      tag_in: in std_logic_vector(tag_width-1 downto 0);
      tag_out: out std_logic_vector(tag_width-1 downto 0);
      env_rdy, accept_rdy: in std_logic;
      f2fi_rdy, f2fo_rdy: out std_logic);
  end component;

  component GenericFloatingPointAdderSubtractor
    generic (name: string;
	     tag_width : integer;
             exponent_width: integer;
             fraction_width : integer;
             round_style : round_type := float_round_style;  -- rounding option
             addguard       : NATURAL := float_guard_bits;  -- number of guard bits
             check_error : BOOLEAN    := float_check_error;  -- check for errors
             denormalize : BOOLEAN    := float_denormalize;  -- Use IEEE extended FP           
             use_as_subtractor: BOOLEAN
      );
    port(
      INA, INB: in std_logic_vector((exponent_width+fraction_width) downto 0);
      OUTADD: out std_logic_vector((exponent_width+fraction_width) downto 0);
      clk,reset: in std_logic;
      tag_in: in std_logic_vector(tag_width-1 downto 0);
      tag_out: out std_logic_vector(tag_width-1 downto 0);
      env_rdy, accept_rdy: in std_logic;
      addi_rdy, addo_rdy: out std_logic);
  end component;

  component GenericFloatingPointMultiplier
    generic (name: string;
	     tag_width : integer;
             exponent_width: integer;
             fraction_width : integer;
             round_style : round_type := float_round_style;  -- rounding option
             addguard       : NATURAL := float_guard_bits;  -- number of guard bits
             check_error : BOOLEAN    := float_check_error;  -- check for errors
             denormalize : BOOLEAN    := float_denormalize  -- Use IEEE extended FP           
             );
    port(
      INA, INB: in std_logic_vector((exponent_width+fraction_width) downto 0);
      OUTMUL: out std_logic_vector((exponent_width+fraction_width) downto 0);
      clk,reset: in std_logic;
      tag_in: in std_logic_vector(tag_width-1 downto 0);
      tag_out: out std_logic_vector(tag_width-1 downto 0);
      env_rdy, accept_rdy: in std_logic;
      muli_rdy, mulo_rdy: out std_logic);
  end component;
  
  component SinglePrecisionMultiplier 
    generic (name: string;
	     tag_width : integer);
    port(
      INA, INB: in std_logic_vector(31 downto 0);
      OUTM: out std_logic_vector(31 downto 0);
      clk,reset: in std_logic;
      tag_in: in std_logic_vector(tag_width-1 downto 0);
      tag_out: out std_logic_vector(tag_width-1 downto 0);
      NaN, oflow, uflow: out std_logic := '0';
      env_rdy, accept_rdy: in std_logic;
      muli_rdy, mulo_rdy: out std_logic);
  end component;

  component DoublePrecisionMultiplier 
    generic (name: string;
	     tag_width : integer);
    port(
      INA, INB: in std_logic_vector(63 downto 0);   
      OUTM: out std_logic_vector(63 downto 0);
      clk,reset: in std_logic;
      tag_in: in std_logic_vector(tag_width-1 downto 0);
      tag_out: out std_logic_vector(tag_width-1 downto 0);
      NaN, oflow, uflow: out std_logic := '0';
      env_rdy, accept_rdy: in std_logic;
      muli_rdy, mulo_rdy: out std_logic);
  end component;

  component PipelinedFPOperator 
    generic (
      name : string;
      operator_id : string;
      exponent_width : integer := 8;
      fraction_width : integer := 23;
      no_arbitration: boolean := true;
      num_reqs : integer := 3; -- how many requesters?
      use_input_buffering: boolean;
      detailed_buffering_per_input : IntegerArray;
      detailed_buffering_per_output : IntegerArray;
      full_rate: boolean
      );
    port (
      -- req/ack follow level protocol
      reqL                     : in BooleanArray(num_reqs-1 downto 0);
      ackR                     : out BooleanArray(num_reqs-1 downto 0);
      ackL                     : out BooleanArray(num_reqs-1 downto 0);
      reqR                     : in  BooleanArray(num_reqs-1 downto 0);
      -- input data consists of concatenated pairs of ips
      dataL                    : in std_logic_vector((2*(exponent_width+fraction_width+1)*num_reqs)-1 downto 0);
      -- output data consists of concatenated pairs of ops.
      dataR                    : out std_logic_vector(((exponent_width+fraction_width+1)*num_reqs)-1 downto 0);
    -- with dataR
    clk, reset              : in std_logic);
  end component;

  component GenericFloatingPointNormalizer is
    generic (name: string;
	     tag_width : integer := 8;
             exponent_width: integer := 11;
             fraction_width : integer := 52;
             round_style : round_type := float_round_style;  -- rounding option
             nguard       : NATURAL := float_guard_bits;  -- number of guard bits
             denormalize : BOOLEAN    := float_denormalize  -- Use IEEE extended FP           
             );
    port(
      fract  :in  unsigned(fraction_width+nguard+1 downto 0);
      expon  :in  signed(exponent_width+1 downto 0);
      sign   :in  std_ulogic;
      sticky :in  std_ulogic;
      tag_in :in  std_logic_vector(tag_width-1 downto 0);
      tag_out:out std_logic_vector(tag_width-1 downto 0);
      in_rdy :in  std_ulogic;
      out_rdy:out std_ulogic;
      stall  :in  std_ulogic;
      clk    :in  std_ulogic;
      reset  :in  std_ulogic;
      normalized_result :out UNRESOLVED_float (exponent_width downto -fraction_width)  -- result
     );
  end component;


  -----------------------------------------------------------------------------
  -- pipelined integer components..
  -----------------------------------------------------------------------------
  component UnsignedMultiplier 
    
    generic (
      name: string;
	     tag_width     : integer;
      operand_width : integer;
      chunk_width   : integer := 8);

    port (
      L, R       : in  unsigned(operand_width-1 downto 0);
      RESULT     : out unsigned((2*operand_width)-1 downto 0);
      clk, reset : in  std_logic;
      in_rdy     : in  std_logic;
      out_rdy    : out std_logic;
      stall      : in std_logic;
      tag_in     : in std_logic_vector(tag_width-1 downto 0);
      tag_out    : out std_logic_vector(tag_width-1 downto 0));
  end component;

  component UnsignedShifter 
  
  generic (
    name: string;
	     shift_right_flag   : boolean;
    tag_width     : integer;
    operand_width : integer;
    shift_amount_width: integer);

  port (
    L       : in  unsigned(operand_width-1 downto 0);
    R       : in  unsigned(shift_amount_width-1 downto 0);
    RESULT     : out unsigned(operand_width-1 downto 0);
    clk, reset : in  std_logic;
    in_rdy     : in  std_logic;
    out_rdy    : out std_logic;
    stall      : in std_logic;
    tag_in     : in std_logic_vector(tag_width-1 downto 0);
    tag_out    : out std_logic_vector(tag_width-1 downto 0));
   end component;

  component UnsignedAdderSubtractor 
  
  generic (
    name: string;
	     tag_width          : integer;
    operand_width      : integer;
    chunk_width        : integer
	);

  port (
    L            : in  unsigned(operand_width-1 downto 0);
    R            : in  unsigned(operand_width-1 downto 0);
    RESULT       : out unsigned(operand_width-1 downto 0);
    subtract_op  : in std_logic;
    clk, reset   : in  std_logic;
    in_rdy       : in  std_logic;
    out_rdy      : out std_logic;
    stall        : in std_logic;
    tag_in       : in std_logic_vector(tag_width-1 downto 0);
    tag_out      : out std_logic_vector(tag_width-1 downto 0));
  end component;



  component GuardInterface is
	generic (name: string;
	     nreqs: integer; delay_flag: boolean);
	port (reqL: in BooleanArray(nreqs-1 downto 0);
	      ackL: out BooleanArray(nreqs-1 downto 0); 
	      reqR: out BooleanArray(nreqs-1 downto 0);
	      ackR: in BooleanArray(nreqs-1 downto 0); 
	      guards: in std_logic_vector(nreqs-1 downto 0); 
	      clk: in std_logic; reset: in std_logic);
  end component;

  component SplitGuardInterfaceBase is
	generic (name: string;
	     buffering:integer);
	port (sr_in: in Boolean;
	      sa_out: out Boolean;
	      sr_out: out Boolean;
	      sa_in: in Boolean;
	      cr_in: in Boolean;
	      ca_out: out Boolean;
	      cr_out: out Boolean;
	      ca_in: in Boolean;
	      guard_interface: in std_logic;
	      clk: in std_logic;
	      reset: in std_logic);
  end component;

  component SplitSampleGuardInterfaceBase is
	generic (name: string;
	     buffering:integer);
	port (sr_in: in Boolean;
	      sa_out: out Boolean;
	      sr_out: out Boolean;
	      sa_in: in Boolean;
	      cr_in: in Boolean;
	      ca_out: out Boolean;
	      cr_out: out Boolean;
	      ca_in: in Boolean;
	      guard_interface: in std_logic;
	      clk: in std_logic;
	      reset: in std_logic);
  end component;

  component SplitUpdateGuardInterfaceBase is
	generic (name: string;
	     buffering:integer);
	port (sr_in: in Boolean;
	      sa_out: out Boolean;
	      sr_out: out Boolean;
	      sa_in: in Boolean;
	      cr_in: in Boolean;
	      ca_out: out Boolean;
	      cr_out: out Boolean;
	      ca_in: in Boolean;
	      guard_interface: in std_logic;
	      clk: in std_logic;
	      reset: in std_logic);
  end component;

  component SgiSampleFsm is
	generic (name: string);
	port (sr_in: in Boolean;
		sr_in_q: out Boolean;
		push_req: out std_logic;
		push_ack: in std_logic;
		clk, reset: in std_logic);
  end component;

  component SgiUpdateFsm is
	generic (name: string);
	port (cr_in: in Boolean;
		cr_out: out Boolean;
		ca_in: in Boolean;
		ca_out: out Boolean;
		pop_req: out std_logic;
		pop_ack: in std_logic;
		pop_data: in std_logic_vector(0 downto 0);
		clk, reset: in std_logic);
  end component;

  component SplitGuardInterface is
	generic (name: string;
	     		nreqs: integer; buffering: IntegerArray; use_guards: BooleanArray;
			sample_only: Boolean; update_only: Boolean);
	port (sr_in: in BooleanArray(nreqs-1 downto 0);
	      sa_out: out BooleanArray(nreqs-1 downto 0); 
	      sr_out: out BooleanArray(nreqs-1 downto 0);
	      sa_in: in BooleanArray(nreqs-1 downto 0); 
	      cr_in: in BooleanArray(nreqs-1 downto 0);
	      ca_out: out BooleanArray(nreqs-1 downto 0); 
	      cr_out: out BooleanArray(nreqs-1 downto 0);
	      ca_in: in BooleanArray(nreqs-1 downto 0); 
	      guards: in std_logic_vector(nreqs-1 downto 0);
	      clk: in std_logic;
	      reset: in std_logic);
  end component;

  
  -----------------------------------------------------------------------------
  -- temporary stuff.
  -----------------------------------------------------------------------------
  component tmpSplitCallArbiter
    generic(num_reqs: integer;
	  call_data_width: integer;
	  return_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
    port ( -- ready/ready handshake on all ports
      -- ports for the caller
      call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
      call_acks   : out std_logic_vector(num_reqs-1 downto 0);
      call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
      call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- call port connected to the called module
      call_mreq   : out std_logic;
      call_mack   : in  std_logic;
      call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
      call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
      -- similarly for return, initiated by the caller
      return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
      return_acks : out std_logic_vector(num_reqs-1 downto 0);
      return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
      return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
      -- return from function
      return_mreq : out std_logic;
      return_mack : in std_logic;
      return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
      return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
      clk: in std_logic;
      reset: in std_logic);
  end component tmpSplitCallArbiter;

  component tmpSplitCallArbiterNoOutargs
    generic(num_reqs: integer;
	  call_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
  end component tmpSplitCallArbiterNoOutargs;

  ----------------------------------------------------------------------------------------
  -- components with per-input buffering
  ----------------------------------------------------------------------------------------

  component UnsharedOperatorWithBuffering 
    generic
    (
      name   : string;
      operator_id   : string;          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer;    -- width of input2
      num_inputs    : integer := 2;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer;          -- width of output.
      constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
      constant_width : integer;
      buffering      : integer;
      use_constant  : boolean := false;
      flow_through : boolean := false;
      full_rate: boolean := false
      );
    port (
      -- req -> ack follow pulse protocol
      reqL:  in Boolean;
      ackL : out Boolean;
      reqR : in Boolean;
      ackR:  out Boolean;
      -- operands.
      dataL      : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
      dataR      : out std_logic_vector(owidth-1 downto 0);
      clk, reset : in  std_logic);
  end component;

  component BinaryLogicalOperator 
  generic
    (
      name  : string;
      operator_id         : string;            -- operator id
      input_width         : integer;           -- input width
      output_width        : integer;           -- the width of the output.
      input_1_buffer_depth: integer;           -- buffering at input 1.
      input_2_buffer_depth: integer;           -- buffering at input 2.
      output_buffer_depth : integer;           -- buffering at output.
	-- both should never be constants.
      input_1_is_constant : boolean := false;
      input_2_is_constant : boolean := false;
      flow_through : boolean := false
      );
  port (
    -- input operands.
    sample_req : in BooleanArray(1 downto 0);  -- sample reqs, one per input.
    sample_ack : out BooleanArray(1 downto 0); -- sample acks, one per output.
    data_in      : in  std_logic_vector((2*input_width)-1 downto 0);
    -- result.
    update_req : in Boolean;  -- req for output update.
    update_ack : out Boolean; -- ack for output update.
    data_out      : out std_logic_vector(output_width-1 downto 0);
    -- clock, reset.
    clk, reset : in  std_logic);
  end component;


  component BinarySharedOperator is
    generic
    (
      name : string;
      operator_id   : string := "ApIntAdd";          -- operator id
      input_1_is_int : Boolean := true; -- false means float
      input_1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input_1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      input_1_width      : integer := 4;    -- width of input1
      input_1_is_constant : BooleanArray;   -- constant case needs to be handled a bit differently..
      input_2_is_int : Boolean := true; -- false means float
      input_2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input_2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      input_2_width      : integer := 0;    -- width of input2
      input_2_is_constant : BooleanArray;  -- constant case needs to be handled a bit differently..
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      output_width        : integer := 4;          -- width of output.
      num_reqs : integer := 3; -- how many requesters?
      input_buffering: integer := 2;
      detailed_buffering_per_output : IntegerArray
    );
  port (
    -- input side.
    sample_req_1                     : in BooleanArray(num_reqs-1 downto 0);
    sample_req_2                     : in BooleanArray(num_reqs-1 downto 0);
    sample_ack_1                     : out BooleanArray(num_reqs-1 downto 0);
    sample_ack_2                     : out BooleanArray(num_reqs-1 downto 0);
    -- output side.
    update_ack                       : out BooleanArray(num_reqs-1 downto 0);
    update_req                       : in  BooleanArray(num_reqs-1 downto 0);
    -- input data consists of concatenated pairs of ips
    data_in_1                    : in std_logic_vector((input_1_width*num_reqs)-1 downto 0);
    data_in_2                    : in std_logic_vector((input_2_width*num_reqs)-1 downto 0);
    -- output data consists of concatenated pairs of ops.
    data_out                    : out std_logic_vector((output_width*num_reqs)-1 downto 0);
    -- with dataR
    clk, reset              : in std_logic);
  end component;


  component LoadReqSharedWithInputBuffers is
    generic
    (
	name : string;
	addr_width: integer := 8;
      	num_reqs : integer := 1; -- how many requesters?
	tag_length: integer := 1;
	no_arbitration: Boolean := false;
        min_clock_period: Boolean := true;
        input_buffering: IntegerArray;
	time_stamp_width: integer := 0
    );
    port (
    -- req/ack follow pulse protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    -- concatenated address corresponding to access
    dataL                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
    -- address to memory
    maddr                   : out std_logic_vector((addr_width)-1 downto 0);
    mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);

    mreq                    : out std_logic;
    mack                    : in std_logic;
    -- clock, reset (active high)
    clk, reset              : in std_logic);
  end component;

  component SelectSplitProtocol is
    generic(name: string; 
	  data_width: integer; 
	  buffering: integer; 
	  flow_through: boolean := false; 
          full_rate: boolean := false);
    port(x,y: in std_logic_vector(data_width-1 downto 0);
       sel: in std_logic_vector(0 downto 0);
       z : out std_logic_vector(data_width-1 downto 0);
       sample_req: in boolean;
       sample_ack: out boolean;
       update_req: in boolean;
       update_ack: out boolean;
       clk,reset: in std_logic);
  end component;

  component StoreReqSharedWithInputBuffers
    generic
    (
	name : string;
	addr_width: integer;
	data_width : integer;
	time_stamp_width : integer;
      	num_reqs : integer; -- how many requesters?
	tag_length: integer;
	no_arbitration: Boolean := false;
        min_clock_period: Boolean := true;
        input_buffering: IntegerArray
    );
    port (
    -- req/ack follow pulse protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    -- address corresponding to access
    addr                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
    data                    : in std_logic_vector((data_width*num_reqs)-1 downto 0);
    -- address to memory
    maddr                   : out std_logic_vector(addr_width-1 downto 0);
    mdata                   : out std_logic_vector(data_width-1 downto 0);
    mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);
    mreq                    : out std_logic;
    mack                    : in std_logic;
    -- clock, reset (active high)
    clk, reset              : in std_logic);
  end component;

  component UnarySharedOperator is
    generic
    (
      name : string;
      operator_id   : string := "ApIntNot";          -- operator id
      input_is_int : Boolean := true; -- false means float
      input_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      input_width      : integer := 4;    -- width of input1
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      output_width        : integer := 4;          -- width of output.
      num_reqs : integer := 3; -- how many requesters?
      detailed_buffering_per_output : IntegerArray
    );
  port (
    -- input side.
    sample_req                     : in BooleanArray(num_reqs-1 downto 0);
    sample_ack                     : out BooleanArray(num_reqs-1 downto 0);
    -- output side.
    update_ack                     : out BooleanArray(num_reqs-1 downto 0);
    update_req                     : in  BooleanArray(num_reqs-1 downto 0);
    -- input data consists of concatenated pairs of ips
    data_in                     : in std_logic_vector((input_width*num_reqs)-1 downto 0);
    -- output data consists of concatenated pairs of ops.
    data_out                    : out std_logic_vector((output_width*num_reqs)-1 downto 0);
    -- with dataR
    clk, reset                  : in std_logic);
  end component;

  component UnaryUnsharedOperator 
    generic
    (
      name          : string;          -- instance name.
      operator_id   : string;          -- operator id
      input_is_int : Boolean := true; -- false means float
      input_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      input_width        : integer;    -- width of input1
      input_is_constant  : boolean; 
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      output_width        : integer;          -- width of output.
      output_buffering : integer := 2
      );
    port (
    -- req -> ack follow pulse protocol
    sample_req:  in Boolean;
    sample_ack:  out Boolean;
    update_req:  in Boolean;
    update_ack:  out Boolean;
    -- operands.
    dataL      : in  std_logic_vector(input_width - 1 downto 0);
    dataR      : out std_logic_vector(output_width-1 downto 0);
    clk, reset : in  std_logic);
  end component;

  -------------------------------------------------------------------------------------
  -- full-rate versions of I/O ports
  -------------------------------------------------------------------------------------
  component InputPortRevised 
    generic(name : string;
	   num_reqs: integer;
	   data_width: integer;
           output_buffering: IntegerArray;
	   nonblocking_read_flag: boolean := false;
	   no_arbitration: boolean := false);
    port (
    -- pulse interface with the data-path
    sample_req        : in  BooleanArray(num_reqs-1 downto 0); -- sacrificial
    sample_ack        : out BooleanArray(num_reqs-1 downto 0); -- sacrificial
    update_req        : in  BooleanArray(num_reqs-1 downto 0);
    update_ack        : out BooleanArray(num_reqs-1 downto 0);
    data       : out std_logic_vector((num_reqs*data_width)-1 downto 0);
    -- ready/ready interface with outside world
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : in  std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
  end component;

  component OutputPortRevised 
    generic(name : string;
	  num_reqs: integer;
	  data_width: integer;
	  no_arbitration: boolean := false;
	  full_rate: boolean;
	  input_buffering : IntegerArray);
    port (
    sample_req        : in  BooleanArray(num_reqs-1 downto 0);
    sample_ack        : out BooleanArray(num_reqs-1 downto 0);
    update_req        : in  BooleanArray(num_reqs-1 downto 0); -- sacrificial
    update_ack        : out BooleanArray(num_reqs-1 downto 0); -- sacrificial
    data       : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : out std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
  end component;

  component InputPort_P2P is
    generic (name : string;
	   data_width: integer;
	   queue_depth: integer;
	   bypass_flag: boolean := false;
	   barrier_flag: boolean := false;
	   nonblocking_read_flag: boolean := false);
    port (
    -- pulse interface with the data-path
     sample_req        : in  Boolean; -- sacrificial.
     sample_ack        : out Boolean; -- sacrificial.
     update_req        : in  Boolean;
     update_ack        : out Boolean;
     data              : out std_logic_vector(data_width-1 downto 0);
    -- ready/ready interface with outside world
     oreq       : out std_logic;
     oack       : in  std_logic;
     odata      : in  std_logic_vector(data_width-1 downto 0);
     clk, reset : in  std_logic);
  end component;

  ---------------------------------------------------------------------------------
  -- some useful miscellaneous stuff
  ---------------------------------------------------------------------------------
  component InputMuxWithBuffering 
    generic (name: string;
	   iwidth: integer := 10;
	   owidth: integer := 10;
	   twidth: integer := 3;
	   nreqs: integer := 1;
	   buffering: IntegerArray;
	   no_arbitration: Boolean := false;
	   full_rate: boolean;
	   registered_output: Boolean := true);
    port (
    -- req/ack follow pulse protocol
    reqL                 : in  BooleanArray(nreqs-1 downto 0);
    ackL                 : out BooleanArray(nreqs-1 downto 0);
    dataL                : in  std_logic_vector(iwidth-1 downto 0);
    -- output side req/ack level protocol
    reqR                 : out std_logic;
    ackR                 : in  std_logic;
    dataR                : out std_logic_vector(owidth-1 downto 0);
    -- tag specifies the requester index 
    tagR                : out std_logic_vector(twidth-1 downto 0);
    clk, reset          : in std_logic);
  end component InputMuxWithBuffering;

  component FullRateRepeater is
    generic(name : string;  data_width: integer := 32);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component FullRateRepeater;

  component NullRepeater is
    generic(name : string;  data_width: integer := 32);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
  end component NullRepeater;

  component LevelRepeater is
    generic(name: string; g_data_width: integer := 32; g_depth: integer := 1);
    port(clk: in std_logic;
       reset: in std_logic;
       enable: in std_logic;
       data_in: in std_logic_vector(g_data_width-1 downto 0);
       valid_in: in std_logic;
       data_out: out std_logic_vector(g_data_width-1 downto 0);
       valid_out : out std_logic;
       stall: in std_logic);
  end component;

  component SquashLevelRepeater is
    generic(name: string; g_data_width: integer := 32; g_depth : integer := 1);
    port(clk: in std_logic;
       		reset: in std_logic;
		enable: in std_logic;
       		data_in: in std_logic_vector(g_data_width-1 downto 0);
       		data_out: out std_logic_vector(g_data_width-1 downto 0);
       		stall_vector: in std_logic_vector(1 to g_depth));
  end component SquashLevelRepeater;

  component ValidPropagator is
    generic(name: string; g_depth : integer := 1);
    port(clk: in std_logic;
       		reset: in std_logic;
       		stall_in: in std_logic;
       		valid_in: in std_logic;
       		valid_out : out std_logic;
       		stall_vector: out std_logic_vector(1 to  g_depth));
  end component ValidPropagator;

  component InterlockBuffer 
    generic (name: string; buffer_size: integer := 2; 
		in_data_width : integer := 32;
		out_data_width : integer := 32;
		flow_through: boolean := false;
		cut_through: boolean  := false;
		bypass_flag : boolean := false); 
    port ( write_req: in boolean;
        write_ack: out boolean;
        write_data: in std_logic_vector(in_data_width-1 downto 0);
        read_req: in boolean;
        read_ack: out boolean;
        read_data: out std_logic_vector(out_data_width-1 downto 0);
        clk : in std_logic;
        reset: in std_logic);
  end component InterlockBuffer;
 
  component InterlockBufferSimplified is
    generic (name: string; buffer_size: integer := 2; data_width : integer := 32);
    port (write_req: in boolean;
        write_ack: out boolean;
        write_data: in std_logic_vector(data_width-1 downto 0);
        read_req: in boolean;
        read_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
        clk : in std_logic;
        reset: in std_logic);
  end component InterlockBufferSimplified;


  component ReceiveBuffer  is
    generic (name: string; buffer_size: integer ; data_width : integer ;
	   		full_rate : boolean );
    port ( write_req: in boolean;
         write_ack: out boolean;
         write_data: in std_logic_vector(data_width-1 downto 0);
         read_req: in std_logic;
         read_ack: out std_logic;
         read_data: out std_logic_vector(data_width-1 downto 0);
         clk : in std_logic;
         reset: in std_logic);
  end component;

  component PulseToLevel 
   port( rL : in boolean;
        rR : out std_logic;
        aL : out boolean;
        aR : in std_logic;
        clk : in std_logic;
        reset : in std_logic);
  end component;

  component PulseToLevelHalfInterlockBuffer 
    generic (name : string; data_width: integer; buffer_size : integer);
    port( sample_req : in boolean;
        sample_ack : out boolean;
        has_room : out std_logic;
        write_enable : in  std_logic;
        write_data : in std_logic_vector(data_width-1 downto 0);
        update_req : in boolean;
        update_ack : out boolean;
        read_data : out std_logic_vector(data_width-1 downto 0);
        clk : in std_logic;
        reset : in std_logic);
  end component;

  component PulseLevelPulseInterlockBuffer 
  generic (name : string; data_width: integer; buffer_size : integer);
  port( write_req : in boolean;
        write_ack : out boolean;
        write_data : in std_logic_vector(data_width-1 downto 0);
        update_req : in boolean;
        update_ack : out boolean;
        has_data    : out std_logic;
        read_enable : in std_logic;
        read_data : out std_logic_vector(data_width-1 downto 0);
        clk : in std_logic;
        reset : in std_logic);
  end component;


  component LevelMux 
    generic(name: string; num_reqs: integer;
	  data_width: integer;
	  no_arbitration: boolean := true);
    port (
    write_req       : in  std_logic_vector(num_reqs-1 downto 0);
    write_ack       : out std_logic_vector(num_reqs-1 downto 0);
    write_data      : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
    read_req        : in  std_logic;
    read_ack        : out std_logic;
    read_data       : out std_logic_vector(data_width-1 downto 0);
    clk, reset      : in  std_logic);
  end component;

  component CounterBase generic(name: string; data_width : integer);
	port(clk, reset: in std_logic; count_out: out std_logic_vector(data_width-1 downto 0));
  end component;

  component UnloadBuffer 
    generic (name: string; buffer_size: integer; data_width : integer; 
				bypass_flag: boolean := false; nonblocking_read_flag: boolean := false;
					use_unload_register: boolean := true);
    port (write_req: in std_logic;
          write_ack: out std_logic;
          write_data: in std_logic_vector(data_width-1 downto 0);
          unload_req: in boolean;
          unload_ack: out boolean;
          read_data: out std_logic_vector(data_width-1 downto 0);
	  has_data: out std_logic;
          clk : in std_logic;
          reset: in std_logic);
  end component UnloadBuffer;
  component UnloadBufferDeep is
    generic (name: string; buffer_size: integer ; data_width : integer ; nonblocking_read_flag : boolean := false);
    port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);
  end component UnloadBufferDeep;
  component UnloadBufferOptimized is
    generic (name: string; buffer_size: integer ; data_width : integer ; 
			bypass_flag, nonblocking_read_flag : boolean := false);
    port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);
  end component UnloadBufferOptimized;
  component UnloadBufferRevised is
    generic (name: string; 
		buffer_size: integer ; 
		data_width : integer ; 
		bypass_flag: boolean := false);
    port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);
  end component;
  component UnloadBufferRevisedNonblocking is
    generic (name: string; 
		buffer_size: integer ; 
		data_width : integer ; 
		bypass_flag: boolean := false);
    port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);
  end component;

  component UnloadRegister is
    generic (name: string; 
		data_width : integer ; 
		bypass_flag: boolean := false;
		nonblocking_read_flag : boolean := false);
    port ( write_req: in std_logic;
           write_ack: out std_logic;
           write_data: in std_logic_vector(data_width-1 downto 0);
           unload_req: in boolean;
           unload_ack: out boolean;
           read_data: out std_logic_vector(data_width-1 downto 0);
           clk : in std_logic;
           reset: in std_logic);
  end component UnloadRegister;

  component UnloadFsm is
  generic (name: string; data_width: integer);
  port ( 
	 write_req: in std_logic;
         write_ack: out std_logic;
         unload_req: in boolean;
         unload_ack: out boolean;
	 data_in :  in std_logic_vector(data_width-1 downto 0);
	 data_out :  out std_logic_vector(data_width-1 downto 0);
         clk : in std_logic;
         reset: in std_logic);
  end component;

  component UnloadFsmNoblock is
  generic (name: string; data_width: integer);
  port ( 
	 write_req: in std_logic;
         write_ack: out std_logic;
         unload_req: in boolean;
         unload_ack: out boolean;
	 data_in :  in std_logic_vector(data_width-1 downto 0);
	 data_out :  out std_logic_vector(data_width-1 downto 0);
         clk : in std_logic;
         reset: in std_logic);
  end component;

  -----------------------------------------------------------------------------------------
  --  System Ports
  -----------------------------------------------------------------------------------------
  component SystemInPort 
   generic (name : string;
	    num_reads: integer;
	    in_data_width: integer;
            out_data_width : integer; 
	    full_rate: boolean := false); 
   port (read_req : in std_logic_vector(num_reads-1 downto 0);
         read_ack : out std_logic_vector(num_reads-1 downto 0);
         read_data: out std_logic_vector((num_reads*out_data_width)-1 downto 0);
         in_data  : in std_logic_vector(in_data_width-1 downto 0);
	 clk : in std_logic;
	 reset : in std_logic);
  end component;

  component SystemOutPort 
   generic (name : string;
	    num_writes: integer;
	    in_data_width: integer;
            out_data_width : integer;
	    full_rate: boolean := false); 
   port (write_req : in std_logic_vector(num_writes-1 downto 0);
         write_ack : out std_logic_vector(num_writes-1 downto 0);
         write_data: in std_logic_vector((num_writes*in_data_width)-1 downto 0);
         out_data  : out std_logic_vector(out_data_width-1 downto 0);
	 clk : in std_logic;
	 reset : in std_logic);
  end component;
 
  component SignalBase is
   generic (name : string;
	    volatile_flag: boolean := false;
	    num_writes: integer;
            data_width : integer); 
   port (
         read_data  : out std_logic_vector(data_width-1 downto 0);
	 write_req : in std_logic_vector(num_writes-1 downto 0);
         write_ack : out std_logic_vector(num_writes-1 downto 0);
         write_data: in std_logic_vector((num_writes*data_width)-1 downto 0);
	 clk : in std_logic;
	 reset : in std_logic);
  end component;

  ----------------------------------------------------------------------------------------------
  -- glue
  ----------------------------------------------------------------------------------------------
  component PipeJoin is
   generic (name : string; data_width_0, data_width_1: integer);
   port (
    write_req_0   : in std_logic;
    write_ack_0   : out std_logic;
    write_data_0   : in std_logic_vector(data_width_0-1 downto 0);
    write_req_1   : in std_logic;
    write_ack_1   : out std_logic;
    write_data_1   : in std_logic_vector(data_width_1-1 downto 0);
    read_req      : in  std_logic;
    read_ack       : out std_logic;
    read_data     : out std_logic_vector((data_width_1 + data_width_0)-1 downto 0);
    clk, reset : in  std_logic);
  end component;

  component PipeMerge is
    generic (name : string; data_width_0, data_width_1: integer);
    port (
      write_req_0   : in std_logic;
      write_ack_0   : out std_logic;
      write_data_0   : in std_logic_vector(data_width_0-1 downto 0);
      write_req_1   : in std_logic;
      write_ack_1   : out std_logic;
      write_data_1   : in std_logic_vector(data_width_1-1 downto 0);
      read_req      : in  std_logic;
      read_ack       : out std_logic;
      read_data     : out std_logic_vector((data_width_1 + data_width_0)-1 downto 0);
      clk, reset : in  std_logic);
  end component;
 
  component PipeMux is
   generic (name : string; data_width: integer);
   port (
    write_req_0   : in std_logic;
    write_ack_0   : out std_logic;
    write_data_0   : in std_logic_vector(data_width-1 downto 0);
    write_req_1   : in std_logic;
    write_ack_1   : out std_logic;
    write_data_1   : in std_logic_vector(data_width-1 downto 0);
    read_req      : in  std_logic;
    read_ack       : out std_logic;
    read_data     : out std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
  end component;

  component PipeSizeMonitor is
   generic (name : string; depth: integer);
   port (
    write_req   : in  std_logic;
    write_ack   : in  std_logic;
    read_req    : in  std_logic;
    read_ack    : in  std_logic;
    has_data    : out Boolean;
    clk, reset  : in  std_logic);
  end component;

  component BypassRegister is
	generic (data_width: integer; bypass: boolean);
	port (clk, reset: in std_logic; 
		enable: in boolean; 
		din: in std_logic_vector(data_width-1 downto 0);
		q: out std_logic_vector(data_width-1 downto 0));
  end component;

  component SingleCycleStartFinFsm is
	port (clk, reset, start_req, fin_req : in std_logic;
		enable, start_ack, fin_ack: out std_logic) ;
  end component SingleCycleStartFinFsm;

  component ram_1024x32_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    enable : in  std_logic_vector(0 downto 0);
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(9 downto 0);
    din : in  std_logic_vector(31 downto 0);
    dout : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component ram_1024x32_Operator;
  component dpram_1w_1r_1024x32_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    read_enable : in  std_logic_vector(0 downto 0);
    write_enable : in  std_logic_vector(0 downto 0);
    read_addr : in  std_logic_vector(9 downto 0);
    write_addr : in  std_logic_vector(9 downto 0);
    write_data : in  std_logic_vector(31 downto 0);
    read_data : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component dpram_1w_1r_1024x32_Operator;

  component module_clock_gate is
	port (reset, start_req, start_ack, fin_req, fin_ack, clock_in: in std_logic;
		clock_out : out std_logic);
  end component module_clock_gate;

  component signal_clock_gate is
	port (reset, clock_in, clock_enable: in std_logic; clock_out : out std_logic);
  end component signal_clock_gate;

  component clock_gater is
	port (clock_in, clock_enable: in std_logic; clock_out : out std_logic);
  end component clock_gater;

end BaseComponents;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- all component declarations necessary for the
-- vhdl generator
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;

package Components is
end Components;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;	
use ieee.std_logic_1164.all;	
use ieee.numeric_std.all;	
	
library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.Utilities.all;
	
library aHiR_ieee_proposed;	
use aHiR_ieee_proposed.math_utility_pkg.all;	
use aHiR_ieee_proposed.fixed_pkg.all;	
use aHiR_ieee_proposed.float_pkg.all;	

package FloatOperatorPackage is

  -----------------------------------------------------------------------------
  -- use the float type directly
  -----------------------------------------------------------------------------
  procedure ApFloatResize_proc(l: in float;
                               constant exponent_width : in integer;
                               constant fraction_width : in integer;                               
                               result : out std_logic_vector);
  procedure ApFloatAdd_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatSub_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatMul_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOeq_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOne_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOgt_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOge_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOlt_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOle_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatOrd_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUno_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUeq_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUne_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUgt_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUge_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUlt_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatUle_proc(l: in float; r : in float; result : out std_logic_vector);
  procedure ApFloatToApIntSigned_proc(l: in float; result : out std_logic_vector);
  procedure ApFloatToApIntUnsigned_proc(l: in float; result : out std_logic_vector);
  procedure ApIntToApFloatSigned_proc(l: in std_logic_vector;
                                      constant exponent_width : in integer;
                                      constant fraction_width : in integer;
                                      result : out std_logic_vector);
  procedure ApIntToApFloatUnsigned_proc(l: in std_logic_vector;
                                      constant exponent_width : in integer;
                                      constant fraction_width : in integer;                                        
                                      result : out std_logic_vector);

  -- TODO
  -- procedures ApFloatToApIntSigned_Proc, ApFloatToApIntUnsigned_Proc,
  --            ApIntSignedToApFloat_Proc, ApIntUnsignedToApFloat_Proc
  procedure TwoInputFloatArithOperation(constant id    : in string;
		  			x, y : in std_logic_vector;
		  			constant exponent_width : in integer;
		  			constant fraction_width : in integer;
					result : out std_logic_vector);
  procedure TwoInputFloatCompareOperation(constant id    : in string;
                                   	x, y : in std_logic_vector;
                                   	constant exponent_width : in integer;
                                   	constant fraction_width : in integer;
                                   	result : out std_logic_vector);
  procedure SingleInputFloatOperation(constant id : in string;
                                      x : in std_logic_vector;
                                      constant exponent_width : in integer;
                                      constant fraction_width : in integer;                                      
                                      result : out std_logic_vector);
  

end package FloatOperatorPackage;

package body FloatOperatorPackage is

  -----------------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatResize_proc (l : in float;
                                constant exponent_width : in integer;
                                constant fraction_width : in integer;
                                result : out std_logic_vector) is					
  begin
     result := To_SLV(RESIZE(l,exponent_width, fraction_width ));
  end ApFloatResize_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatAdd_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApFloatAdd_proc" severity error;
     result := To_SLV(l+r);  
  end ApFloatAdd_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatSub_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApFloatSub_proc" severity error;
     result := To_SLV(l-r);  
  end ApFloatSub_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatMul_proc (l : in float; r : in float; result : out std_logic_vector) is
    variable float_result  : float(l'left downto l'right);
  begin
    assert (l'length = r'length)
      report "input operand length mismatch in ApFloatMul_proc" severity error;
    assert (l'length = result'length)						     
      report "input and output operand length mismatch in ApFloatMul_proc" severity error;
    float_result := l*r;  
    result := To_SLV(float_result);  
  end ApFloatMul_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOeq_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(l=r);  
  end ApFloatOeq_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOne_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(l /= r);  
  end ApFloatOne_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOgt_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(l > r);  
  end ApFloatOgt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOge_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(l >= r);  
  end ApFloatOge_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOlt_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(l < r);  
  end ApFloatOlt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOle_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(l <= r); 
  end ApFloatOle_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatOrd_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(not(Unordered (x => l,y => r))); 
  end ApFloatOrd_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUno_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(Unordered (x => l,y => r)); 
  end ApFloatUno_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUeq_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(eq(l => l, r => r, check_error => false) or Unordered (x => l,y => r)); 
  end ApFloatUeq_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUne_proc (l : in float; r : in float; result : out std_logic_vector) is					
  begin
     result :=  To_SLV(ne(l => l, r => r, check_error => false) or Unordered (x => l,y => r));
  end ApFloatUne_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUgt_proc (l : in float; r : in float; result : out std_logic_vector) is					
	variable cr: boolean;
  begin
     cr :=  gt(l => l, r => r, check_error => false) or Unordered (x => l,y => r);
     result :=  To_SLV(cr);
  end ApFloatUgt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUge_proc (l : in float; r : in float; result : out std_logic_vector) is					
	variable cr: boolean;
  begin
     cr :=  ge(l => l, r => r, check_error => false) or Unordered (x => l,y => r);  
     result(result'low) :=  to_std_logic(cr);
  end ApFloatUge_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUlt_proc (l : in float; r : in float; result : out std_logic_vector) is					
	variable cr: boolean;
  begin
     cr :=  lt(l => l, r => r, check_error => false) or Unordered (x => l,y => r); 
     result(result'low) := to_std_logic(cr);
  end ApFloatUlt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatUle_proc (l : in float; r : in float; result : out std_logic_vector) is					
	variable cr: boolean;
  begin
     cr :=  le(l => l, r => r, check_error => false) or Unordered (x => l,y => r);  
     result(result'low) := to_std_logic(cr);
  end ApFloatUle_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatToApIntSigned_proc (l : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(to_signed(l,result'length));
  end ApFloatToApIntSigned_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApFloatToApIntUnsigned_proc (l : in float; result : out std_logic_vector) is					
  begin
     result := To_SLV(to_unsigned(l,result'length));
  end ApFloatToApIntUnsigned_proc; 				

 ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntToApFloatSigned_proc (l : in std_logic_vector;
                                       constant exponent_width : in integer;
                                       constant fraction_width : in integer;
                                       result : out std_logic_vector) is
  begin
   result := To_SLV(to_float(to_signed(l),exponent_width,fraction_width,round_zero));
  end ApIntToApFloatSigned_proc;
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntToApFloatUnsigned_proc (l : in std_logic_vector;
                                         constant exponent_width : in integer;
                                         constant fraction_width : in integer;                                         
                                         result : out std_logic_vector) is
  begin
   result := To_SLV(to_float(to_unsigned(l),exponent_width, fraction_width,round_zero));
  end ApIntToApFloatUnsigned_proc;
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------	
  procedure TwoInputFloatArithOperation(constant id : in string;
                                   x, y : in std_logic_vector;
                                   constant exponent_width : in integer;
                                   constant fraction_width : in integer;
                                   result : out std_logic_vector) is	
    variable result_var : std_logic_vector(exponent_width+fraction_width downto 0);	
    variable temp_int: integer;
  begin
    result_var:= (others => '0');
    if id = "ApFloatAdd" then					
      ApFloatAdd_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatSub" then					
      ApFloatSub_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatMul" then					
      ApFloatMul_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    else	
      assert false report "Unsupported arithmetic float operator-id " & id severity failure;	
    end if;	
    result := result_var;	
  end TwoInputFloatArithOperation;			

  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------	
  procedure TwoInputFloatCompareOperation(constant id : in string;
                                   x, y : in std_logic_vector;
                                   constant exponent_width : in integer;
                                   constant fraction_width : in integer;
                                   result : out std_logic_vector) is	
    variable result_var : std_logic_vector(0 downto 0);
    variable temp_int: integer;
  begin

    assert(result'length = 1) report "comparison result must be a 1-bit integer" severity error;

    result_var:= (others => '0');
    if id = "ApFloatOeq" then					
      ApFloatOeq_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatOne" then					
      ApFloatOne_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatOgt" then					
      ApFloatOgt_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatOge" then					
      ApFloatOge_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatOlt" then					
      ApFloatOlt_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatOle" then					
      ApFloatOle_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatOrd" then					
      ApFloatOrd_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUno" then					
      ApFloatUno_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUeq" then					
      ApFloatUeq_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUne" then					
      ApFloatUne_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUgt" then					
      ApFloatUgt_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUge" then					
      ApFloatUge_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUlt" then					
      ApFloatUlt_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatUle" then					
      ApFloatUle_proc(To_Float(x,exponent_width,fraction_width), To_Float(y,exponent_width,fraction_width), result_var);
    else	
      assert false report "Unsupported float comparison operator-id " & id severity failure;	
    end if;	
    result(result'low) := result_var(0);	
  end TwoInputFloatCompareOperation;			

  -----------------------------------------------------------------------------
  -----------------------------------------------------------------------------	
  procedure SingleInputFloatOperation(constant id : in string;
                                      x : in std_logic_vector;
                                      constant exponent_width : in integer;
                                      constant fraction_width : in integer;                                      
                                      result : out std_logic_vector) is	
    variable result_var : std_logic_vector(result'length-1 downto 0);	
  begin
    result_var:= (others => '0');
    if id = "ApFloatToApIntSigned" then					
      ApFloatToApIntSigned_proc(To_Float(x,exponent_width,fraction_width), result_var);
    elsif id = "ApFloatToApIntUnsigned" then					
      ApFloatToApIntUnsigned_proc(To_Float(x,exponent_width,fraction_width), result_var);
    elsif id = "ApIntToApFloatSigned" then					
      ApIntToApFloatSigned_proc(x, exponent_width, fraction_width, result_var);
    elsif id = "ApIntToApFloatUnsigned" then					
      ApIntToApFloatUnsigned_proc(x, exponent_width, fraction_width, result_var);
    else	
      assert false report "Unsupported operator-id " & id severity failure;	
    end if;	
    result := result_var;	
  end SingleInputFloatOperation;	
	
  
	
end package body FloatOperatorPackage;	
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;	
use ieee.std_logic_1164.all;	
use ieee.numeric_std.all;	
	
library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.Utilities.all;
	
package OperatorPackage is

  procedure ApConcat_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApBitsel_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntNot_proc(l: in std_logic_vector; result : out std_logic_vector);
  procedure ApIntToApIntSigned_proc(l: in std_logic_vector; result : out std_logic_vector);
  procedure ApIntToApIntUnsigned_proc(l: in std_logic_vector; result : out std_logic_vector);
  procedure ApIntAdd_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntSub_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntAnd_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntNand_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntOr_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntNor_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntXor_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntXnor_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntMul_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntSHL_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntLSHR_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntASHR_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntROL_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntROR_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntEq_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntNe_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntUgt_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntUge_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntUlt_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntUle_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntSgt_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntSge_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntSlt_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);
  procedure ApIntSle_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector);

  -- TODO
  -- procedures ApFloatToApIntSigned_Proc, ApFloatToApIntUnsigned_Proc,
  --            ApIntSignedToApFloat_Proc, ApIntUnsignedToApFloat_Proc

  procedure TwoInputOperation(constant id    : in string; x, y : in std_logic_vector; result : out std_logic_vector);
  procedure SingleInputOperation(constant id : in string; x : in std_logic_vector; result : out std_logic_vector);

  function isTrue(l: in std_logic_vector) return boolean;
  function areEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function uGreaterThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function uGreaterEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function uLessThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function uLessEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function sGreaterThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function sGreaterEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function sLessThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function sLessEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector;
  function Mux2to1 (sel: std_logic_vector; x, y : std_logic_vector) return
		std_logic_vector;

end package OperatorPackage;

package body OperatorPackage is

  -----------------------------------------------------------------------------
  procedure ApConcat_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is
  begin
      result := l & r;
  end procedure;
  -----------------------------------------------------------------------------
  procedure ApBitsel_proc(l: in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is
    variable temp_int: integer;
    alias ll : std_logic_vector (l'length-1 downto 0) is l; 
  begin

      temp_int := To_Integer(To_Unsigned(Ceil_Log2(l'length),r));
      result(result'low) := '0';

      for I in ll'low to ll'high loop
           if (I = temp_int) then
              result(result'low) := ll (I);
           end if;
      end loop;

  end procedure;
  -----------------------------------------------------------------------------
  procedure ApIntNot_proc (l : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = result'length)						     
      report "Length Mismatch inApIntNot_proc" severity error;
    result := To_SLV(not to_signed(l));
  end ApIntNot_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntToApIntSigned_proc (l : in std_logic_vector; result : out std_logic_vector) is					
  begin
     result := To_SLV(RESIZE(to_signed(l), result'length));
  end ApIntToApIntSigned_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntToApIntUnsigned_proc (l : in std_logic_vector; result : out std_logic_vector) is					
  begin
    result := To_SLV(RESIZE(to_unsigned(l), result'length));
  end ApIntToApIntUnsigned_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntAdd_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntAdd_proc" severity error;
    result := To_SLV(to_signed(l)  + to_signed(r));
  end ApIntAdd_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntSub_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntSub_proc" severity error;
    result := To_SLV(to_signed(l)  - to_signed(r));
  end ApIntSub_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntAnd_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntAnd_proc" severity error;
    result := l and r;
  end ApIntAnd_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntNand_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntNand_proc" severity error;
    result := not ( l and r );
  end ApIntNand_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntOr_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntOr_proc" severity error;
    result := l or r;
  end ApIntOr_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntNor_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntNor_proc" severity error;
    result := not (l or r);
  end ApIntNor_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntXor_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntXor_proc" severity error;
    result := l xor r;
  end ApIntXor_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntXnor_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntXnor_proc" severity error;
    result := not (l xor r);
  end ApIntXnor_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntMul_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    assert (l'length = r'length) and (l'length = result'length)						     
      report "Length Mismatch inApIntMul_proc" severity error;
     result := To_SLV(resize((to_unsigned(l)  * to_unsigned(r)),result'length));
  end ApIntMul_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntSHL_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    result := To_SLV(to_unsigned(l) sll to_integer(to_unsigned(Ceil_Log2(l'length)+1, r)));
  end ApIntSHL_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntLSHR_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
     result := To_SLV(to_unsigned(l)  srl to_integer(to_unsigned(Ceil_Log2(l'length)+1, r)));
  end ApIntLSHR_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntASHR_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
     result := To_SLV(shift_right(to_signed(l), to_integer(to_unsigned(Ceil_Log2(l'length)+1,r)))); 
  end ApIntASHR_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntROL_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    result := To_SLV(to_unsigned(l) rol to_integer(to_unsigned(Ceil_Log2(l'length)+1, r)));
  end ApIntROL_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntROR_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    result := To_SLV(to_unsigned(l) ror to_integer(to_unsigned(Ceil_Log2(l'length)+1, r)));
  end ApIntROR_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntEq_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if l = r then
      result(result'low) := '1';
    else
      result(result'low) := '0';
    end if;
  end ApIntEq_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntNe_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if l = r then
      result(result'low) := '0';
    else
      result(result'low) := '1';
    end if;
  end ApIntNe_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntUgt_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_unsigned(l)  > to_unsigned(r) then
      result(result'low) := '1';
    else
      result(result'low) := '0';
    end if;
  end ApIntUgt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntUge_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin

    if to_unsigned(l)  >= to_unsigned(r) then
      result(result'low) := '1';      
    else
      result(result'low) := '0';
    end if;    

  end ApIntUge_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntUlt_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_unsigned(l)  < to_unsigned(r) then
      result(result'low) := '1';            
    else
      result(result'low) := '0';      
    end if;        

  end ApIntUlt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntUle_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_unsigned(l)  <= to_unsigned(r) then
      result(result'low) := '1';            
    else
      result(result'low) := '0';            
    end if;        
  end ApIntUle_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntSgt_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_signed(l)  > to_signed(r) then
      result(result'low) := '1';            
    else
      result(result'low) := '0';                  
    end if;        
  end ApIntSgt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntSge_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_signed(l)  >= to_signed(r) then
      result(result'low) := '1';            
    else
      result(result'low) := '0';                  
    end if;        

  end ApIntSge_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntSlt_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_signed(l) < to_signed(r) then
      result(result'low) := '1';                        
    else
      result(result'low) := '0';                              
    end if;        

  end ApIntSlt_proc; 				
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure ApIntSle_proc (l : in std_logic_vector; r : in std_logic_vector; result : out std_logic_vector) is					
  begin
    if to_signed(l) <= to_signed(r) then
      result(result'low) := '1';                              
    else
      result(result'low) := '0';                              
    end if;        
    
  end ApIntSle_proc;
  ---------------------------------------------------------------------
  -----------------------------------------------------------------------------
  procedure TwoInputOperation(constant id : in string; x, y : in std_logic_vector; result : out std_logic_vector) is	
    variable result_var : std_logic_vector(result'high downto result'low);	
  begin
    if id = "ApConcat" then
      ApConcat_proc(x,y,result_var);
    elsif id = "ApBitsel" then
      ApBitsel_proc(x,y,result_var);
    elsif id = "ApIntAdd" then					
      ApIntAdd_proc(x,y, result_var);
    elsif id = "ApIntSub" then					
      ApIntSub_proc(x, y, result_var);
    elsif id = "ApIntAnd" then					
      ApIntAnd_proc(x, y, result_var);
    elsif id = "ApIntNand" then					
      ApIntNand_proc(x, y, result_var);
    elsif id = "ApIntOr" then					
      ApIntOr_proc(x, y, result_var);
    elsif id = "ApIntNor" then					
      ApIntNor_proc(x, y, result_var);
    elsif id = "ApIntXor" then					
      ApIntXor_proc(x, y, result_var);
    elsif id = "ApIntXnor" then					
      ApIntXnor_proc(x, y, result_var);
    elsif id = "ApIntMul" then					
      ApIntMul_proc(x, y, result_var);
    elsif id = "ApIntSHL" then					
      ApIntSHL_proc(x, y, result_var);
    elsif id = "ApIntLSHR" then					
      ApIntLSHR_proc(x, y, result_var);
    elsif id = "ApIntASHR" then					
      ApIntASHR_proc(x, y, result_var);
    elsif id = "ApIntROL" then					
      ApIntROL_proc(x, y, result_var);
    elsif id = "ApIntROR" then					
      ApIntROR_proc(x, y, result_var);
    elsif id = "ApIntEq" then					
      ApIntEq_proc(x, y, result_var);
    elsif id = "ApIntNe" then					
      ApIntNe_proc(x, y, result_var);
    elsif id = "ApIntUgt" then					
      ApIntUgt_proc(x, y, result_var);
    elsif id = "ApIntUge" then					
      ApIntUge_proc(x, y, result_var);
    elsif id = "ApIntUlt" then					
      ApIntUlt_proc(x, y, result_var);
    elsif id = "ApIntUle" then					
      ApIntUle_proc(x, y, result_var);
    elsif id = "ApIntSgt" then					
      ApIntSgt_proc(x, y, result_var);
    elsif id = "ApIntSge" then					
      ApIntSge_proc(x, y, result_var);
    elsif id = "ApIntSlt" then					
      ApIntSlt_proc(x, y, result_var);
    elsif id = "ApIntSle" then					
      ApIntSle_proc(x, y, result_var);
    else	
      assert false report "Unsupported operator-id " & id severity failure;	
    end if;	
    result := result_var;	
  end TwoInputOperation;			
  -----------------------------------------------------------------------------
	
  -----------------------------------------------------------------------------	
  procedure SingleInputOperation(constant id : in string; x : in std_logic_vector; result : out std_logic_vector) is	
    variable result_var : std_logic_vector(result'high downto result'low);	
  begin
    if id = "ApIntNot" then					
      ApIntNot_proc(x, result_var);
    elsif id = "ApIntToApIntSigned" then					
      ApIntToApIntSigned_proc(x, result_var);
    elsif id = "ApIntToApIntUnsigned" then					
      ApIntToApIntUnsigned_proc(x, result_var);
-- synopsys translate_off
    elsif id = "ApIntDecode" then					
      result_var := GenericDecode(x);
-- synopsys translate_on
    elsif id = "ApIntEncode" then					
      result_var := GenericEncode(x);
    elsif id = "ApIntPriorityEncode" then					
      result_var := PriorityEncode(x);
    elsif id = "ApIntBitreduceOr" then					
      result_var(result_var'low) := OrReduce(x);
    elsif id = "ApIntBitreduceAnd" then					
      result_var(result_var'low) := AndReduce(x);
    elsif id = "ApIntBitreduceXor" then					
      result_var(result_var'low) := XorReduce(x);
    else	
      assert false report "Unsupported operator-id " & id severity failure;	
    end if;	
    result := result_var;	
  end SingleInputOperation;	
	
  -----------------------------------------------------------------------------
   -- useful function forms.	
  -----------------------------------------------------------------------------	
  function isTrue(l: in std_logic_vector) return boolean is
	variable ret_val: boolean;
        variable r_or : std_logic;
	alias ll : std_logic_vector(1 to l'length) is l;
  begin
	
	r_or := '0';
	for I in 1 to l'length loop
		r_or := (r_or or ll(I));
	end loop;

	if(r_or /= '0')  then
		ret_val := true;
	else
		ret_val := false;
	end if;
	return(ret_val);
  end function;

  function areEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if (l = r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
	
  function uGreaterThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_unsigned(l)  > to_unsigned(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;

  function uGreaterEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_unsigned(l)  >= to_unsigned(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
  function uLessThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_unsigned(l)  < to_unsigned(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
  function uLessEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_unsigned(l)  <= to_unsigned(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
  function sGreaterThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_signed(l)  > to_signed(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
  function sGreaterEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_signed(l)  >= to_signed(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
  function sLessThan(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_signed(l)  < to_signed(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;
  function sLessEqual(l: in std_logic_vector; r : in std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(0 downto 0);
  begin
    if to_signed(l)  <= to_signed(r) then
      ret_var(0) := '1';
    else
      ret_var(0) := '0';
    end if;
    return(ret_var);
  end function;

  function Mux2to1 (sel: std_logic_vector; x, y : std_logic_vector) return std_logic_vector is
	variable ret_var : std_logic_vector(1 to x'length);
	alias lsel: std_logic_vector(sel'length downto 1) is sel;
  begin
	assert(x'length = y'length) report "inputs to mux not of same width" severity error;
	if(lsel(1) = '1') then
		ret_var := x;
	else
		ret_var := y;
	end if;
	return(ret_var);
  end Mux2to1;

end package body OperatorPackage;	
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package mem_component_pack is
component mem_demux 
  generic ( name: string;
	    g_data_width: natural;
            g_id_width : natural;
            g_number_of_outputs: natural;
	    g_delay_count: natural);
  port(data_in: in std_logic_vector(g_data_width-1 downto 0);  -- data & id & time-stamp
       sel_in : in std_logic_vector(g_id_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0 );
       req_out: out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clk: in std_logic;
       reset: in std_logic);
end component;

component mem_repeater 
    generic(name: string;
	    g_data_width: natural);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(g_data_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector(g_data_width-1 downto 0);
       req_out : out std_logic;
       ack_in: in std_logic);
end component mem_repeater;

component mem_shift_repeater
    generic(name: string;
	    g_data_width: natural; g_number_of_stages: natural);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(g_data_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector(g_data_width-1 downto 0);
       req_out : out std_logic;
       ack_in: in std_logic);
end component mem_shift_repeater;


component memory_bank 
   generic (
     name: string;
     g_addr_width: natural;
     g_data_width: natural;
     g_write_tag_width : natural;
     g_read_tag_width : natural;
     g_time_stamp_width: natural;
     g_base_bank_addr_width: natural;
     g_base_bank_data_width: natural
	);
   port (
     clk : in std_logic;
     reset: in std_logic;
     write_data     : in  std_logic_vector(g_data_width-1 downto 0);
     write_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     write_tag      : in std_logic_vector(g_write_tag_width-1 downto 0);
     write_tag_out  : out std_logic_vector(g_write_tag_width-1 downto 0);
     write_enable   : in std_logic;
     write_ack   : out std_logic;
     write_result_accept : in std_logic;
     write_result_ready : out std_logic;
     read_data     : out  std_logic_vector(g_data_width-1 downto 0);
     read_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     read_tag      : in std_logic_vector(g_read_tag_width-1 downto 0);
     read_tag_out  : out std_logic_vector(g_read_tag_width-1 downto 0);
     read_enable   : in std_logic;
     read_ack      : out std_logic;
     read_result_accept: in std_logic;
     read_result_ready: out std_logic
     );
end component memory_bank;

component memory_bank_revised is
   generic (
     name: string;
     g_addr_width: natural;
     g_data_width: natural;
     g_write_tag_width : natural;
     g_write_port_id_width : natural;
     g_read_tag_width : natural;
     g_read_port_id_width : natural;
     g_time_stamp_width: natural;
     g_base_bank_addr_width: natural;
     g_base_bank_data_width: natural
	);
   port (
     clk : in std_logic;
     reset: in std_logic;
     write_data     : in  std_logic_vector(g_data_width-1 downto 0);
     write_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     write_tag      : in std_logic_vector(g_write_tag_width-1 downto 0);
     write_time_stamp: in std_logic_vector(g_time_stamp_width-1 downto 0);
     write_tag_out  : out std_logic_vector(g_write_tag_width-1 downto 0);
     write_port_id      : in unsigned(g_write_port_id_width-1 downto 0);
     write_port_id_out  : out unsigned(g_write_port_id_width-1 downto 0);
     write_enable   : in std_logic;
     write_ack   : out std_logic;
     write_result_accept : in std_logic;
     write_result_ready : out std_logic;
     read_data     : out std_logic_vector(g_data_width-1 downto 0);
     read_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     read_tag      : in std_logic_vector(g_read_tag_width-1 downto 0);
     read_time_stamp: in std_logic_vector(g_time_stamp_width-1 downto 0);
     read_tag_out  : out std_logic_vector(g_read_tag_width-1 downto 0);
     read_port_id      : in unsigned(g_read_port_id_width-1 downto 0);
     read_port_id_out  : out unsigned(g_read_port_id_width-1 downto 0);
     read_enable   : in std_logic;
     read_ack      : out std_logic;
     read_result_accept: in std_logic;
     read_result_ready: out std_logic
     );
end component memory_bank_revised;

component memory_bank_base 
   generic ( name: string;
	g_addr_width: natural; 
	g_data_width : natural;
        g_base_bank_addr_width: natural;
        g_base_bank_data_width: natural);
   port (data_in : in std_logic_vector(g_data_width-1 downto 0);
         data_out: out std_logic_vector(g_data_width-1 downto 0);
         addr_in: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         write_bar : in std_logic;
         clk: in std_logic;
         reset : in std_logic
	);
end component memory_bank_base;

component base_bank 
   generic ( name: string;
	g_addr_width: natural; g_data_width : natural);
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component base_bank;

component base_bank_dual_port is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component base_bank_dual_port;

-- single write, read port register file.
component register_file_1w_1r_port is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
         -- write port 0
         datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         -- read port 1 
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;

         clk: in std_logic;
         reset : in std_logic);
end component register_file_1w_1r_port;

-- with write to read bypass.
component register_file_1w_1r_port_with_bypass is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
         -- write port 0
         datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         -- read port 1 
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;

         clk: in std_logic;
         reset : in std_logic);
end component register_file_1w_1r_port_with_bypass;

component fifo_mem_synch_write_asynch_read is
   generic ( name: string; address_width: natural;  data_width : natural;
			mem_size: natural);
   port (
	 write_enable: in std_logic;
	 write_data: in std_logic_vector(data_width-1 downto 0);
	 write_address: in std_logic_vector(address_width-1 downto 0);
	 read_data: out std_logic_vector(data_width-1 downto 0);
	 read_address: in std_logic_vector(address_width-1 downto 0);
         clk: in std_logic);
end component fifo_mem_synch_write_asynch_read;

component base_bank_dual_port_for_vivado is
   generic ( name: string;  g_addr_width: natural := 10; g_data_width : natural := 16);
	port(
		clka : in std_logic;
		clkb : in std_logic;
		ena : in std_logic;
		enb : in std_logic;
		wea : in std_logic;
		web : in std_logic;
		addra : in std_logic_vector(g_addr_width-1 downto 0);
		addrb : in std_logic_vector(g_addr_width-1 downto 0);
		dia : in std_logic_vector(g_data_width-1 downto 0);
		dib : in std_logic_vector(g_data_width-1 downto 0);
		doa : out std_logic_vector(g_data_width-1 downto 0);
		dob : out std_logic_vector(g_data_width-1 downto 0)
		);
end component base_bank_dual_port_for_vivado;

component base_bank_dual_port_for_xst is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component base_bank_dual_port_for_xst;

component base_bank_with_registers
   generic ( name: string;
	g_addr_width: natural; g_data_width : natural);
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component base_bank_with_registers;

component base_bank_dual_port_with_registers is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component base_bank_dual_port_with_registers;

component register_file_1w_1r_port_with_registers  is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component register_file_1w_1r_port_with_registers ;

component merge_box_with_repeater 
  generic (name: string;
	   g_data_width: natural;
           g_number_of_inputs: natural;
           g_number_of_outputs: natural;
           g_time_stamp_width : natural;   -- width of timestamp
           g_tag_width : natural;  -- width of tag
           g_pipeline_flag: integer     -- if 0, dont add pipe-line stage
           );            

  port(data_left: in  std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
       req_in : in std_logic_vector(g_number_of_inputs-1 downto 0);
       ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
       data_right: out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
       req_out : out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clock: in std_logic;
       reset: in std_logic);

end component merge_box_with_repeater;


component merge_tree 
  generic (
    name: string;
    g_number_of_inputs: natural;          
    g_data_width: natural;          -- total width of data
                                          -- (= actual-data & timestamp)
    g_time_stamp_width : natural;   -- width of timestamp
    g_tag_width : natural;          -- width of tag
    g_mux_degree :natural;         -- max-indegree of each pipeline-stage
    g_num_stages : natural;
    g_port_id_width: natural
    );       

  port (
    merge_data_in : in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    merge_req_in  : in std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_data_out: out std_logic_vector(g_data_width-1 downto 0);
    merge_req_out : out std_logic;
    merge_ack_in  : in std_logic;
    clock: in std_logic;
    reset: in std_logic);
  
end component merge_tree;

component demerge_tree 
  
  generic (
     name: string;
    g_demux_degree: natural;
    g_number_of_outputs: natural;
    g_data_width: natural;              -- total width of data
                                        -- (= data & tag & port-id & timestamp)
    g_id_width: natural;
    g_stage_id: natural
    );       

  port (
    demerge_data_out : out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
    demerge_ready_out  : out std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_accept_in   : in std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_data_in: in std_logic_vector(g_data_width-1 downto 0);
    demerge_ack_out : out std_logic;
    demerge_req_in  : in std_logic;
    demerge_sel_in: in std_logic_vector(g_id_width-1 downto 0);
    clock: in std_logic;
    reset: in std_logic);
  
end component demerge_tree;

component demerge_tree_wrap
  
  generic (
     name: string;
    g_demux_degree: natural;
    g_number_of_outputs: natural;
    g_data_width: natural;              -- total width of data
                                        -- (= data & tag & port-id & timestamp)
    g_id_width: natural;
    g_stage_id: natural
    );       

  port (
    demerge_data_out : out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
    demerge_ready_out  : out std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_accept_in   : in std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_data_in: in std_logic_vector(g_data_width-1 downto 0);
    demerge_ack_out : out std_logic;
    demerge_req_in  : in std_logic;
    demerge_sel_in: in std_logic_vector(g_id_width-1 downto 0);
    clock: in std_logic;
    reset: in std_logic);
  
end component demerge_tree_wrap;

component combinational_merge 
  generic (
     name: string;
    g_data_width       : natural;
    g_number_of_inputs: natural;
    g_time_stamp_width : natural);
  port(
    in_data: in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    in_tstamp: in std_logic_vector((g_number_of_inputs*g_time_stamp_width)-1 downto 0);
    out_data: out std_logic_vector(g_data_width-1 downto 0);
    out_tstamp: out std_logic_vector(g_time_stamp_width-1 downto 0);
    in_req: in std_logic_vector(g_number_of_inputs-1 downto 0);
    in_ack: out std_logic_vector(g_number_of_inputs-1 downto 0);
    out_req: out std_logic;
    out_ack: in std_logic);
end component combinational_merge;

component combinational_merge_with_repeater
  generic (
     name: string;
    g_data_width       : natural;
    g_number_of_inputs: natural;
    g_time_stamp_width : natural);
  port(
    clk : in std_logic;
    reset : in std_logic;
    in_data: in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    in_tstamp: in std_logic_vector((g_number_of_inputs*g_time_stamp_width)-1 downto 0);
    out_data: out std_logic_vector(g_data_width-1 downto 0);
    out_tstamp: out std_logic_vector(g_time_stamp_width-1 downto 0);
    in_req: in std_logic_vector(g_number_of_inputs-1 downto 0);
    in_ack: out std_logic_vector(g_number_of_inputs-1 downto 0);
    out_req: out std_logic;
    out_ack: in std_logic);
end component combinational_merge_with_repeater;


component memory_subsystem_core
  generic (
    name: string;
    num_loads       : natural;
    num_stores      : natural;
    addr_width      : natural;
    data_width      : natural;
    tag_width       : natural;
    time_stamp_width    : natural;
    number_of_banks : natural;
    mux_degree      : natural;
    demux_degree    : natural;
    base_bank_addr_width: natural;
    base_bank_data_width: natural);
  port (
    lr_addr_in  : in  std_logic_vector((num_loads*addr_width)-1 downto 0);
    lr_req_in   : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out  : out std_logic_vector(num_loads-1 downto 0);
    lr_tag_in   : in  std_logic_vector((num_loads*tag_width)-1 downto 0);
    lr_time_stamp_in   : in  std_logic_vector((num_loads*time_stamp_width)-1 downto 0);
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);
    lc_req_in   : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out  : out std_logic_vector(num_loads-1 downto 0);
    lc_tag_out  : out std_logic_vector((num_loads*tag_width)-1 downto 0);
    sr_addr_in  : in  std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in  : in  std_logic_vector((num_stores*data_width)-1 downto 0);
    sr_req_in   : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out  : out std_logic_vector(num_stores-1 downto 0);
    sr_tag_in   : in  std_logic_vector((num_stores*tag_width)-1 downto 0);
    sr_time_stamp_in   : in  std_logic_vector((num_stores*time_stamp_width)-1 downto 0);
    sc_req_in   : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out  : out std_logic_vector(num_stores-1 downto 0);
    sc_tag_out  : out std_logic_vector((num_stores*tag_width)-1 downto 0);
    clock       : in  std_logic;
    reset       : in  std_logic);
end component;

component CombinationalMux is
  generic (
     name: string;
    g_data_width       : integer := 32;
    g_number_of_inputs: integer := 2);
  port(
    in_data: in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    out_data: out std_logic_vector(g_data_width-1 downto 0);
    in_req: in std_logic_vector(g_number_of_inputs-1 downto 0);
    in_ack: out std_logic_vector(g_number_of_inputs-1 downto 0);
    out_req: out std_logic;
    out_ack: in std_logic);
end component CombinationalMux;

component PipelinedMux is
  generic (
     name: string;
    g_number_of_inputs: natural;          
    g_data_width: natural;          -- total width of data
                                        -- (= actual-data & tag & port_id)
    g_mux_degree :natural;         -- max-indegree of each pipeline-stage
    g_port_id_width: natural
    );       

  port (
    merge_data_in : in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    merge_req_in  : in std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_data_out: out std_logic_vector(g_data_width-1 downto 0);
    merge_req_out : out std_logic;
    merge_ack_in  : in std_logic;
    clock: in std_logic;
    reset: in std_logic);
  
end component PipelinedMux;

component PipelinedMuxStage is 
  generic (name: string;
	   g_data_width: integer := 10;
           g_number_of_inputs: integer := 8;
           g_number_of_outputs: integer := 1;
           g_tag_width : integer := 3  -- width of tag
           );            

  port(data_left: in  std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
       req_in : in std_logic_vector(g_number_of_inputs-1 downto 0);
       ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
       data_right: out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
       req_out : out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clock: in std_logic;
       reset: in std_logic);

end component PipelinedMuxStage;

component PipelinedDemux is
  generic ( name: string;
	    g_data_width: natural := 10;
            g_destination_id_width : natural := 3;
            g_number_of_outputs: natural := 8);
  port(data_in: in std_logic_vector(g_data_width-1 downto 0);  -- data & destination-id 
       sel_in : in std_logic_vector(g_destination_id_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0 );
       req_out: out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clk: in std_logic;
       reset: in std_logic);
end component;

component spram_generic_reverse_wrapper is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR : in std_logic_vector(address_width-1 downto 0 );
		CLK : in std_logic;
		WRITE_BAR: in std_logic;
		ENABLE_BAR: in std_logic;
		DATAIN  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT  : out std_logic_vector(data_width-1 downto 0));
end component spram_generic_reverse_wrapper;

component dpram_generic_reverse_wrapper is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		WRITE_0_BAR : in std_logic;
		WRITE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAIN_1  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_0  : out std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK : in std_logic);
end component dpram_generic_reverse_wrapper;

component register_file_1w_1r_generic_reverse_wrapper is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK: in std_logic);
end component;

component spmem_column is
   generic ( name: string:="spmem_column"; 
	g_addr_width: natural := 2;
	g_base_bank_addr_width: natural:=4; 
	g_base_bank_data_width : natural := 4);
   port (datain : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         dataout: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component spmem_column;

component spmem_selector_array is
   generic ( name: string:="mem";
		 g_addr_width: natural := 5; 
	      	 g_data_width : natural := 20;
		 g_base_addr_width: natural := 5; 
	      	 g_base_data_width : natural := 20
	   );
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component;

component spmem_selector is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR : in std_logic_vector(address_width-1 downto 0 );
		CLK : in std_logic;
	        RESET: in std_logic;
		WRITE_BAR: in std_logic;
		ENABLE_BAR: in std_logic;
		DATAIN  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT  : out std_logic_vector(data_width-1 downto 0));
end component spmem_selector;

component dpmem_column is
   generic (name: string:="dpmem_column"; 
	g_addr_width: natural := 2;
	g_base_bank_addr_width: natural:=4; 
	g_base_bank_data_width : natural := 4);
   port (datain_0 : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component dpmem_column;

component dpmem_selector_array is
   generic ( name: string:="mem";
		 g_addr_width: natural := 5; 
	      	 g_data_width : natural := 20;
		 g_base_addr_width: natural := 5; 
	      	 g_base_data_width : natural := 20
	   );
   port (datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component;

component dpmem_selector is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		WRITE_0_BAR : in std_logic;
		WRITE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAIN_1  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_0  : out std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK, RESET: in std_logic);
end component dpmem_selector;

component register_file_1w_1r_column is
   generic ( name: string:="register_file_1w_1r_column"; 
	g_addr_width: natural := 2;
	g_base_bank_addr_width: natural:=4; 
	g_base_bank_data_width : natural := 4);
   port (datain_0 : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         dataout_1: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component register_file_1w_1r_column;


component register_file_1w_1r_selector_array is
   generic ( name: string:="mem";
		 g_addr_width: natural := 5; 
	      	 g_data_width : natural := 20;
		 g_base_addr_width: natural := 5; 
	      	 g_base_data_width : natural := 20
	   );
   port (datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end component;

component register_file_1w_1r_selector is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK, RESET: in std_logic);
end component register_file_1w_1r_selector;

end package mem_component_pack;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
                         
package mem_function_pack is
  function Ceil_Log ( x: natural; base: natural) return natural;
  function Ceil_Log2 ( x: natural) return natural;
  function Ceiling (constant x, y : integer) return integer;
  function IsGreaterThan(x, y: std_logic_vector) return boolean;
  function IncrementSLV(constant x : std_logic_vector) return std_logic_vector;
  function Bank_Match(BANK: natural;
                      log2_number_of_banks: natural;
                      addr_in: std_logic_vector)   return boolean;
  function To_Integer(x: std_logic_vector) return natural;
  function Digit_To_Char(val: integer) return character;
  function Minimum(x: integer; y: integer) return integer;
  function Maximum(x: integer; y: integer) return integer;
  function Natural_To_SLV (constant val, size : natural) return std_logic_vector;

  function Convert_To_String(val : natural) return STRING; -- convert val to string.
  function Convert_Integer_To_String(val : integer) return STRING; -- convert val to string.
  function Convert_To_String(val : std_logic_vector) return STRING; -- convert signed to string.

end mem_function_pack;

package body mem_function_pack is
  function Ceil_Log ( x: natural; base: natural ) return natural is
    variable ret_var : integer := 0;
    variable tvar : natural;
  begin
    ret_var := 0;
    if(x > 0) then
      tvar := x;
      while(tvar > 1)loop
        tvar := tvar/base;
        ret_var := ret_var + 1;
      end loop;
      if(base**ret_var < x) then ret_var := ret_var + 1; end if;
    end if;
    return(ret_var);
  end function Ceil_Log;

  function Ceil_Log2 ( x: natural) return natural is
  begin
    return(Ceil_Log(x,2));
  end function Ceil_Log2;
    
  -- purpose: ceiling of x/y
  function Ceiling (
    constant x, y : integer)
    return integer is
    variable ratio : integer;
  begin  -- Ceiling
    ratio := x/y;
    if(y*ratio < x) then
      ratio := ratio + 1;
    end if;
    return ratio;
  end Ceiling;

    -- return true if x > y false otherwise
  function IsGreaterThan(x, y: std_logic_vector) return boolean is
    alias lx : std_logic_vector(1 to x'length) is x;
    alias ly : std_logic_vector(1 to x'length) is y;
    variable ret_val, still_equal : boolean;
  begin
    assert lx'length = ly'length report "mismatched lengths in IsGreaterThan" severity error;
    assert lx'length > 2 report "time-stamp length must be > 2 in IsGreaterThan" severity error;

    ret_val := false;
    
    if((lx(1 to 2) = "00" and ly(1 to 2) = "11") or
       (lx(1 to 2) = "01" and ly(1 to 2) = "00") or
       (lx(1 to 2) = "10" and ly(1 to 2) = "01") or
       (lx(1 to 2) = "11" and ly(1 to 2) = "10")) then
      ret_val := true;
    elsif(lx(1 to 2) = ly(1 to 2)) then
      still_equal := true;
      for I in 3 to lx'length loop
        if(still_equal and (lx(I) = '1') and (ly(I) = '0')) then
          ret_val := true;
          still_equal := false;
        elsif(still_equal and (lx(I) = '0' and ly(I) = '1')) then
          still_equal := false;
        end if;
      end loop;  -- I
    end if;
    return(ret_val);
  end function IsGreaterThan;

  function IncrementSLV(constant x : std_logic_vector) return std_logic_vector
  is
    alias lx : std_logic_vector(1 to x'length) is x;
    variable ret_var : std_logic_vector(1 to x'length);
    variable carry_bit, sum_bit : std_logic;
  begin
    carry_bit := '1';
    for I in x'length downto 1 loop
      sum_bit    := carry_bit xor lx(I);
      carry_bit  := carry_bit and lx(I);
      ret_var(I) := sum_bit;
    end loop;
    return(ret_var);
  end function  IncrementSLV;

  function Bank_Match(BANK: natural;
                      log2_number_of_banks: natural;
                      addr_in: std_logic_vector)
    return boolean is
    alias la : std_logic_vector(1 to addr_in'length) is addr_in;
    variable v : unsigned(1 to log2_number_of_banks);
    variable ret_val : boolean;
  begin
    assert addr_in'length > log2_number_of_banks report "inadequate address length in Bank_Match" severity error;
    ret_val := true;
    if(log2_number_of_banks > 0) then
      for I  in 1 to log2_number_of_banks loop
        v(I) := la((addr_in'length - log2_number_of_banks) + I);
      end loop;  -- I
      if(To_Integer(v) = BANK) then
        ret_val := true;
      else
        ret_val := false;
      end if;
    end if;
    return(ret_val);
  end Bank_Match;

  function To_Integer(x: std_logic_vector) return natural is
	alias lx: std_logic_vector(1 to x'length) is x;
	variable ret_var,two_power: natural;
  begin
        two_power := 1; 
        ret_var := 0;
	for I in x'length downto 1 loop
		if(lx(I) = '1') then
			ret_var := ret_var  + two_power;
		end if;
		two_power := 2*two_power;
	end loop;
	return(ret_var);
  end To_Integer;
  
  function Minimum(x: integer; y: integer) return integer is
       variable ret_var: integer;
    begin
       if(x < y) then ret_var := x; else ret_var := y; end if;
       return(ret_var);
  end Minimum; 

  function Maximum(x: integer; y: integer) return integer is
       variable ret_var: integer;
    begin
       if(x > y) then ret_var := x; else ret_var := y; end if;
       return(ret_var);
  end Maximum; 

  function Natural_To_SLV (constant val, size : natural) return std_logic_vector is
    variable ret_var  : std_logic_vector(size-1 downto 0);
    variable uret_var : unsigned(size-1 downto 0);
    variable scale_val : natural;
  begin
    scale_val := val mod (2**size);
    uret_var := TO_UNSIGNED(scale_val,size);
    for I in 0 to size-1 loop
      ret_var(I) := uret_var(I);
    end loop;  -- I
    return(ret_var);
  end Natural_To_SLV;

  function Convert_To_String(val : NATURAL) return STRING is
	variable result : STRING(10 downto 1) := (others => '0'); -- smallest natural, longest string
	variable pos    : NATURAL := 1;
	variable tmp, digit  : NATURAL;
  begin
    -- synopsys translate_off
	tmp := val;
	loop
		digit := abs(tmp MOD 10);
	    	tmp := tmp / 10;
	    	result(pos) := character'val(character'pos('0') + digit);
	    	pos := pos + 1;
	    	exit when tmp = 0;
	end loop;
    -- synopsys translate_on
	return result((pos-1) downto 1);
  end Convert_To_String;

  function Digit_To_Char(val: integer) return character is
	variable ret_val : character;
  begin
	case val is
		when 0 => ret_val := '0';
		when 1 => ret_val := '1';
		when 2 => ret_val := '2';
		when 3 => ret_val := '3';
		when 4 => ret_val := '4';
		when 5 => ret_val := '5';
		when 6 => ret_val := '6';
		when 7 => ret_val := '7';
		when 8 => ret_val := '8';
		when 9 => ret_val := '9';
		when others => ret_val := 'X';
	end case;
	return(ret_val);
  end Digit_To_Char;


    -- Thanks to: D. Calvet calvet@hep.saclay.cea.fr
    -- modified to support negative values
  function Convert_Integer_To_String(val : integer) return STRING is
	variable result : STRING(12 downto 1) := (others => '0'); -- smallest natural, longest string
	variable pos    : NATURAL := 1;
	variable tmp : integer;
	variable digit  : NATURAL;
	variable is_negative : boolean;
  begin
	tmp := val;
	if val < 0 then
	  tmp := -val;
	end if;
	is_negative := val < 0;
	
	loop
		digit := abs(tmp MOD 10);
	    	tmp := tmp / 10;
	    	result(pos) := Digit_To_Char(digit);
	    	pos := pos + 1;
	    	exit when ((tmp = 0) or (pos = (result'high-1)));
	end loop;
	
	if is_negative then
	  result(pos) := '-';
	  pos := pos + 1;
	end if;
	
	return result((pos-1) downto 1);
  end Convert_Integer_To_String;
  

  function Convert_To_String(val : std_logic_vector) return STRING is
        alias lval: std_logic_vector(1 to val'length) is val;
	variable result : STRING(1 to val'length) := (others => '0'); -- smallest natural, longest string
  begin
        for I in 1 to val'length loop
          if(lval(I) = '0') then result(I) := '0'; else result(I) := '1'; end if;
	end loop;
	return result;
  end Convert_To_String;

end mem_function_pack;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package memory_subsystem_package is

  component memory_subsystem
    generic (
      name: string;
      num_loads       : natural;
      num_stores      : natural;
      addr_width      : natural;
      data_width      : natural;
      tag_width       : natural;
      number_of_banks : natural; -- must be a power of 2!
      mux_degree      : natural;
      demux_degree    : natural;
      base_bank_addr_width: natural;
      base_bank_data_width: natural);
    port (
      lr_addr_in  : in  std_logic_vector((num_loads*addr_width)-1 downto 0);
      lr_req_in   : in  std_logic_vector(num_loads-1 downto 0);
      lr_ack_out  : out std_logic_vector(num_loads-1 downto 0);
      lr_tag_in   : in  std_logic_vector((num_loads*tag_width)-1 downto 0);
      lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);
      lc_req_in   : in  std_logic_vector(num_loads-1 downto 0);
      lc_ack_out  : out std_logic_vector(num_loads-1 downto 0);
      lc_tag_out  : out std_logic_vector((num_loads*tag_width)-1 downto 0);
      sr_addr_in  : in  std_logic_vector((num_stores*addr_width)-1 downto 0);
      sr_data_in  : in  std_logic_vector((num_stores*data_width)-1 downto 0);
      sr_req_in   : in  std_logic_vector(num_stores-1 downto 0);
      sr_ack_out  : out std_logic_vector(num_stores-1 downto 0);
      sr_tag_in   : in  std_logic_vector((num_stores*tag_width)-1 downto 0);
      sc_req_in   : in  std_logic_vector(num_stores-1 downto 0);
      sc_ack_out  : out std_logic_vector(num_stores-1 downto 0);
      sc_tag_out  : out std_logic_vector((num_stores*tag_width)-1 downto 0);
      clock       : in  std_logic;
      reset       : in  std_logic);
  end component;


  component register_bank 
    generic(name: string;
             num_loads             : natural := 5;
            num_stores            : natural := 10;
            addr_width            : natural := 9;
            data_width            : natural := 5;
            tag_width             : natural := 7;
            num_registers         : natural := 1);
    port(
      ------------------------------------------------------------------------------
      -- load request ports
      ------------------------------------------------------------------------------
      lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

      -- req/ack pair:
      -- when both are asserted, time-stamp is set on load request.
      lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
      lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

      -- tag for request, will be returned on completion.
      lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

      ---------------------------------------------------------------------------
      -- load complete ports
      ---------------------------------------------------------------------------
      lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

      -- req/ack pair:
      -- when both are asserted, user should latch data_out.
      lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
      lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

      -- tag of completed request.
      lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

      ------------------------------------------------------------------------------
      -- store request ports
      ------------------------------------------------------------------------------
      sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
      sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

      -- req/ack pair:
      -- when both are asserted, time-stamp is set on store request.
      sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
      sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

      -- tag for request, will be returned on completion.
      sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

      ---------------------------------------------------------------------------
      -- store complete ports
      ---------------------------------------------------------------------------
      -- req/ack pair:
      -- when both are asserted, user assumes that store is done.
      sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
      sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

      -- tag of completed request.
      sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

      ------------------------------------------------------------------------------
      -- clock, reset
      ------------------------------------------------------------------------------
      clock : in std_logic;  -- only rising edge is used to trigger activity.
      reset : in std_logic               -- active high.
      );
  end component register_bank;

  component  dummy_read_only_memory_subsystem 
  generic(name:string;
	  num_loads             : natural := 5;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
   end component dummy_read_only_memory_subsystem;

   component dummy_write_only_memory_subsystem is
  	generic( name:string;
	  num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7);
  	port(
    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
    end component dummy_write_only_memory_subsystem;

component ordered_memory_subsystem is
  generic(name: string;
          num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          time_stamp_width      : natural := 0;
          number_of_banks       : natural := 1;
          mux_degree            : natural := 10;
          demux_degree          : natural := 10;
	  base_bank_addr_width  : natural := 8;
	  base_bank_data_width  : natural := 8);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag + timestamp: tag will be returned on completion..
    lr_tag_in : in std_logic_vector((num_loads*(tag_width+time_stamp_width))-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*(tag_width+time_stamp_width))-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end component ordered_memory_subsystem;

component UnorderedMemorySubsystem is
  generic(name: string;
          num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          -- number_of_banks       : natural := 1; (will always be 1 in this memory)
          mux_degree            : natural := 10;
          demux_degree          : natural := 10;
	  base_bank_addr_width  : natural := 8;
	  base_bank_data_width  : natural := 8);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end component UnorderedMemorySubsystem;


end memory_subsystem_package;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;

package merge_functions is
  type NaturalArray is array (natural range <>) of natural;

  function Total_Intermediate_Width(constant x,y: natural) return natural;
  function Stage_Width (
    constant stage_id     : natural;
    constant mux_degree : natural;
    constant stage0_width : natural)
    return natural;
  function Left_Index (
    constant stage_id     : natural;
    constant mux_degree : natural;
    constant stage0_width : natural)
    return natural;
  function Right_Index (
    constant stage_id     : natural;
    constant mux_degree : natural;
    constant stage0_width : natural)
    return natural;
  
  --constant c_group_left_id : NaturalArray(0 to c_demux_degree-1) := Calculate_Group_Left_Ids(g_number_of_outputs,c_demux_degree);
  function Calculate_Group_Left_Ids (
    constant xwid : natural;
    constant x : natural;
    constant y : natural)
    return NaturalArray;
  
  --constant c_group_right_id : NaturalArray(0 to c_demux_degree-1) := Calculate_Group_Left_Ids(g_number_of_outputs,c_demux_degree);
  function Calculate_Group_Right_Ids (
    constant xwid : natural;
    constant x : natural;
    constant y : natural)
    return NaturalArray;
  
  --constant c_group_sizes : NaturalArray(0 to c_demux_degree-1) := Calculate_Group_Sizes(g_number_of_outputs,c_demux_degree);
  function Calculate_Group_Sizes (
    constant xwid : natural;
    constant x : natural;
    constant y : natural)
    return NaturalArray;

  function Nonzero_Count (
    constant x : NaturalArray)
    return natural;

  procedure Select_Best_Index(time_stamp_vector : in std_logic_vector;
                              data_vector: in std_logic_vector;
			      valid_vector      : in std_logic_vector;
			      best_time_stamp   : out std_logic_vector;
                              best_data : out std_logic_vector;
                              sel_vector: out std_logic_vector;
                              valid_flag: out std_logic);
end merge_functions;

package body merge_functions is

  function Total_Intermediate_Width(constant x,y: natural)
    return natural is
    variable ret_val,tval : natural;
  begin
    ret_val := x;
    tval := x;
    
    while tval > 1 loop
      tval := Ceiling(tval,y);
      ret_val := ret_val + tval;
    end loop;  -- I

    -- for the output.
    ret_val := ret_val + 1;
    return(ret_val);
  end function Total_Intermediate_Width;

  function Stage_Width (
    constant stage_id     : natural;
    constant mux_degree : natural;
    constant stage0_width : natural)
    return natural is
    variable ret_var,tval : natural;
  begin  -- Stage_Width
    ret_var := stage0_width;
    tval := mux_degree;
    if(stage_id > 0) then
      for I  in 1 to stage_id loop
        ret_var := Ceiling(ret_var,tval);
      end loop;  -- I
    end if;
    return(ret_var);
  end Stage_Width;
  
  -- index in intermediate array from which input to stage_id begins
  function Left_Index (
    constant stage_id     : natural;
    constant mux_degree : natural;
    constant stage0_width : natural)
    return natural is
    variable ret_var,offset,tval : natural;
  begin  
    if(stage_id = 0) then
      ret_var := 0;
    else
      ret_var := Right_Index(stage_id-1,mux_degree,stage0_width) + 1;
    end if;
    return(ret_var);
  end Left_Index;

  function Right_Index (
    constant stage_id     : natural;
    constant mux_degree : natural;
    constant stage0_width : natural)
    return natural is
    variable ret_var: natural;
  begin  
    ret_var := Left_Index(stage_id,mux_degree,stage0_width)  +
               Stage_Width(stage_id,mux_degree,stage0_width) - 1;
    return(ret_var);
  end Right_Index;

  function Calculate_Group_Left_Ids (
    constant xwid : natural;
    constant x : natural;
    constant y : natural)
    return NaturalArray is
    variable ret_var  : NaturalArray(0 to y-1);

    constant ysize : natural := Ceil_Log2(y);
    constant xsize : natural := Maximum(xwid,ysize);    

    variable index : natural;
    variable xbin: std_logic_vector(xsize-1 downto 0);
    variable ybin : std_logic_vector(ysize-1 downto 0);
  begin
--    assert false report "left-id called " & Convert_To_String(xwid) & " " &
--		Convert_To_String(x) & " " & Convert_To_String(y) severity note;
    ret_var := (others => x);
    if(xsize >= ysize) then
      for I in x-1 downto 0 loop
        xbin := Natural_To_SLV(I,xsize);
        ybin := xbin(xsize-1 downto xsize-ysize);
        index := To_Integer(ybin);
        if(ret_var(index) = x) then
          ret_var(index) := I;
        end if;
      end loop;  -- I
    end if;
--    for I in 0 to y-1 loop
--      assert false report "group-left-id " & Convert_To_String(ret_var(I)) severity note;
--    end loop;
    return(ret_var);
  end Calculate_Group_Left_Ids;
  

  function Calculate_Group_Right_Ids (
    constant xwid : natural;
    constant x : natural;
    constant y : natural)
    return NaturalArray is
    variable ret_var  : NaturalArray(0 to y-1);

    constant ysize : natural := Ceil_Log2(y);
    constant xsize : natural := Maximum(xwid,ysize);    

    variable index : natural;
    variable xbin: std_logic_vector(xsize-1 downto 0);
    variable ybin : std_logic_vector(ysize-1 downto 0);
  begin
--    assert false report "right-id called " & Convert_To_String(xwid) & " " &
--		Convert_To_String(x) & " " & Convert_To_String(y) severity note;
    ret_var := (others => x);
    if(xsize >= ysize) then
      for I in 0 to x-1 loop
        xbin := Natural_To_SLV(I,xsize);
        ybin := xbin(xsize-1 downto xsize-ysize);
        index := To_Integer(ybin);
        if(ret_var(index) = x) then
          ret_var(index) := I;
        end if;
      end loop;  -- I
    end if;
--    for I in 0 to y-1 loop
--      assert false report "group-right-id " & Convert_To_String(ret_var(I)) severity note;
--    end loop;
    return(ret_var);
  end Calculate_Group_Right_Ids;


  function Calculate_Group_Sizes (
    constant xwid : natural;
    constant x : natural;
    constant y : natural)
    return NaturalArray is
    variable ret_var  : NaturalArray(0 to y-1);

    constant ysize : natural := Ceil_Log2(y);
    constant xsize : natural := Maximum(xwid,ysize);

    variable index : natural;
    variable xbin: std_logic_vector(xsize-1 downto 0);
    variable ybin : std_logic_vector(ysize-1 downto 0);
  begin
--    assert false report "group-sizes called " & Convert_To_String(xwid) & " " &
--		Convert_To_String(x) & " " & Convert_To_String(y) severity note;
    ret_var := (others => 0);
    if(xsize >= ysize) then 
      for I in x-1 downto 0 loop
        xbin := Natural_To_SLV(I,xsize);
        ybin := xbin(xsize-1 downto xsize-ysize);
        index := To_Integer(ybin);
        ret_var(index) := ret_var(index) + 1;
      end loop;  -- I
    end if;
--    for I in 0 to y-1 loop
--      assert false report "group-size " & Convert_To_String(ret_var(I)) severity note;
--    end loop;
    return(ret_var);
  end Calculate_Group_Sizes;

  function Nonzero_Count (
    constant x : NaturalArray)
    return natural is
    variable ret_var : natural;
    alias lx : NaturalArray(1 to x'length) is x;
  begin
    ret_var := 0;
    for I in 1 to x'length loop
      if(lx(I) > 0) then
        ret_var := ret_var + 1;
      end if;
    end loop;  -- I
--    assert false report "non-zero-count " & Convert_To_String(ret_var) severity note;
    return(ret_var);
  end Nonzero_Count;
    
  procedure Select_Best_Index(time_stamp_vector : in std_logic_vector;
                              data_vector: in std_logic_vector;
			      valid_vector      : in std_logic_vector;
			      best_time_stamp   : out std_logic_vector;
                              best_data : out std_logic_vector;
                              sel_vector: out std_logic_vector;
                              valid_flag: out std_logic)
  is
	constant mid_point: integer := valid_vector'length / 2;
        constant time_stamp_width : integer := best_time_stamp'length;
        constant data_width : integer := best_data'length;
        
        alias ltv: std_logic_vector(1 to time_stamp_vector'length) is time_stamp_vector;
        alias ld: std_logic_vector(1 to data_vector'length) is data_vector;
	alias lv: std_logic_vector(1 to valid_vector'length) is valid_vector;

	variable uindex, hindex: integer;
	variable ubest, hbest: std_logic_vector(1 to time_stamp_width);
        variable ud, hd: std_logic_vector(1 to data_width);
        variable sv : std_logic_vector(1 to lv'length) ;
        variable uvalid,hvalid : std_logic;
  begin
        sv := (others => '0');
        valid_flag := '0';
	best_time_stamp := ltv(1 to time_stamp_width);
        best_data := ld(1 to data_width);

	if(valid_vector'length = 1) then
		if(lv(1) = '1') then
                        sv(1) := '1';
                        valid_flag := '1';
		end if;	
	elsif(valid_vector'length = 2) then
		if(lv(1) = '1' and lv(2) = '1') then
			if(IsGreaterThan(ltv(1 to time_stamp_width),ltv(time_stamp_width+1 to (2*time_stamp_width)))) then
				best_time_stamp := ltv(time_stamp_width+1 to 2*time_stamp_width);
                                best_data := ld(data_width+1 to 2*data_width);
                                sv(2) := '1';
			else
                                sv(1) := '1';
			end if;
                        valid_flag := '1';
		elsif(lv(1) = '1') then
                        sv(1) := '1';
                        valid_flag := '1';
		elsif(lv(2) = '1') then
			best_time_stamp := ltv(time_stamp_width+1 to 2*time_stamp_width);
                        best_data := ld(data_width+1 to 2*data_width);
                        sv(2) := '1';
                        valid_flag := '1';
		end if;
	else
		Select_Best_Index(ltv(1 to mid_point*time_stamp_width),
                                  ld(1 to mid_point*data_width),
                                  lv(1 to mid_point),
                                  ubest,
                                  ud,
                                  sv(1 to mid_point),
                                  uvalid);
                
		Select_Best_Index(ltv((mid_point*time_stamp_width)+1 to ltv'length),
                                  ld((mid_point*data_width)+1 to ld'length),
                                  lv(mid_point+1 to lv'length),
                                  hbest,
                                  hd,
                                  sv(mid_point+1 to sv'length),
                                  hvalid);
                
		if(uvalid = '1' and hvalid = '1') then
			if(IsGreaterThan(hbest,ubest)) then
				best_time_stamp := ubest;
                                best_data := ud;
                                sv(mid_point + 1 to sv'length) := (others => '0');
			else
				best_time_stamp := hbest;
                                best_data := hd;
                                sv(1 to mid_point) := (others => '0');
			end if;
                        valid_flag := '1';
		elsif (hvalid = '1' ) then
			best_time_stamp := hbest;
                        best_data := hd;
                        sv(1 to mid_point) := (others => '0');
                        valid_flag := '1';
		elsif(uvalid = '1') then
			best_time_stamp := ubest;
                        best_data := ud;
                        sv(mid_point + 1 to sv'length) := (others => '0');
                        valid_flag := '1';
		end if;
	end if;
        sel_vector := sv;
  end Select_Best_Index;
end merge_functions;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;                  
use aHiR_ieee_proposed.float_pkg.all;


package functionLibraryComponents is

component fpadd32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpadd32;

component fpmul32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpmul32;

component fpsub32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpsub32;

component fpu32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      OP_ID : in std_logic_vector(7 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpu32;


component fpadd64 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpadd64;


component fpsub64 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpsub64;

component fpmul64 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpmul64;


component fpu64 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      OP_ID : in std_logic_vector(7 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component fpu64;

component getClockTime is -- 
    generic (tag_length : integer);
    port ( -- 
      clock_time : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component getClockTime;

component countDownTimer is -- 
    generic (tag_length : integer);
    port ( -- 
      time_count : in  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component countDownTimer;

component umul32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component umul32;

component umul32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end component umul32_Operator;

component ushift32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      shift_right_flag: in std_logic_vector(0 downto 0);
      signed_flag: in std_logic_vector(0 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component ushift32;

component ushift32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      shift_right_flag: in std_logic_vector(0 downto 0);
      signed_flag: in std_logic_vector(0 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end component ushift32_Operator;

component uaddsub32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      carry_in: in std_logic_vector(0 downto 0);
      carry_out: out std_logic_vector(0 downto 0);
      subtract_flag: in std_logic_vector(0 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end component uaddsub32;

component uaddsub32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      carry_in: in std_logic_vector(0 downto 0);
      carry_out: out std_logic_vector(0 downto 0);
      subtract_flag: in std_logic_vector(0 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end component uaddsub32_Operator;

end package;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ApIntComponents is

 component UnsignedAdderSubtractor_n_n_n is
  
  generic (
    name	       : string;
    tag_width          : integer;
    operand_width      : integer;
    chunk_width        : integer
	);

  port (
    slv_L            : in  std_logic_vector(operand_width-1 downto 0);
    slv_R            : in  std_logic_vector(operand_width-1 downto 0);
    slv_RESULT       : out std_logic_vector(operand_width-1 downto 0);
    slv_carry_out    : out std_logic;
    slv_carry_in     : in std_logic;  
    subtract_op      : in std_logic;
    clk, reset       : in  std_logic;
    in_rdy           : in  std_logic;
    out_rdy          : out std_logic;
    stall            : in std_logic;
    tag_in           : in std_logic_vector(tag_width-1 downto 0);
    tag_out          : out std_logic_vector(tag_width-1 downto 0));

 end component;

 component UnsignedMultiplier_n_n_2n is
  
  generic (
    name: string;
    tag_width     : integer;
    operand_width : integer;
    chunk_width   : integer := 16);

  port (
    slv_L, slv_R   : in  std_logic_vector(operand_width-1 downto 0);
    slv_RESULT     : out std_logic_vector((2*operand_width)-1 downto 0);
    clk, reset : in  std_logic;
    in_rdy     : in  std_logic;
    out_rdy    : out std_logic;
    stall      : in std_logic;
    tag_in     : in std_logic_vector(tag_width-1 downto 0);
    tag_out    : out std_logic_vector(tag_width-1 downto 0));
 end component;

 component UnsignedShifter_n_n_n is
  generic (
    name: string;
    tag_width          : integer;
    operand_width      : integer;
    shift_amount_width : integer);

  port (
    slv_L       : in  std_logic_vector(operand_width-1 downto 0);
    slv_R       : in  std_logic_vector(shift_amount_width-1 downto 0);
    slv_RESULT  : out std_logic_vector(operand_width-1 downto 0);
    clk, reset  : in  std_logic;
    in_rdy      : in  std_logic;
    out_rdy     : out std_logic;
    stall       : in std_logic;
    shift_right_flag   : in std_logic;
    signed_flag        : in std_logic;
    tag_in      : in std_logic_vector(tag_width-1 downto 0);
    tag_out     : out std_logic_vector(tag_width-1 downto 0));
 end component;

 component GenericBinaryApIntArithOperatorPipelined is
  generic (
	    name : string;
	    op_id: string;
	    tag_width : integer := 8;
	    in_operand_width: integer;
	    out_result_width: integer
           );
  port(
    inA, inB: in std_logic_vector(in_operand_width-1 downto 0);
    outR: out std_logic_vector(out_result_width-1 downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    pipeline_stall: in std_logic;
    env_rdy: in std_logic;
    op_o_rdy: out std_logic);
 end component;

 component GenericApIntArithOperator is
  generic (
	    name: string;
	    op_id: string;
	    tag_width : integer := 8;
	    in_operand_width: integer;
	    num_non_constant_inputs: integer;
            first_operand_is_constant: boolean;
            second_operand_is_constant: boolean;
	    constant_value: std_logic_vector;
	    out_result_width: integer
           );
  port(
    in_data: in std_logic_vector((num_non_constant_inputs*in_operand_width)-1 downto 0);
    out_data: out std_logic_vector(out_result_width-1 downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    env_rdy, accept_rdy: in std_logic;
    op_i_rdy, op_o_rdy: out std_logic);
 end component;
end package;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;
--use ahir.Utilities.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

package MemCutsPackage is

	-- For a requirement of a memory with MxN (M-rows, N-columns) aspect
	-- ratio, we will first determine uniform columns to implement the
	-- memory.  For each available memory cut, we will find the number
	-- of column-replications that will be filled by it.  For example,
	-- if we have a requirement of 64x24, we could have the following
	-- solutions
	--       column of 16x4 replicated 6 times 
	--       column of 16x4 replicated 2 times, column of 32x16 replicated once
	--  etc.
	--
	
	-- Using the procedure 'opt_find' for a given MxN array, the cut that
	-- maximally covers the N with minimum number of column-replications 
	-- subject to cut utilization of atleast 50% is found out. This procedure
	-- also outputs the number of columns left after filling the N with optimal 
	-- column-replications.
	
	-- To fill the N completely, 'opt_find' is called recursively in the 
	-- function 'find_n_cols', each time passing the number of columns 
	-- yet to be filled. 'find_n_cols' returns an array containg the number
	-- of columns of each available cut required, index-wise.
	
	-- A column memory of size (Mxcut_data_width) for a given cut is build 
	-- using the entity 'mem_column'. This entity is instantiated for
	-- the number of column-replications of each cut. Thus, forming the 
	-- complete MxN array.

	-- functions developed and their description are given in the package body.

	procedure Min_array(x: in IntegerArray;
		    y: in IntegerArray; 
		    min: out integer;
		    index: out integer );
	
	procedure opt_find (constant cut_address_widths: IntegerArray;
		constant cut_data_widths: IntegerArray;
		constant cut_row_heights: IntegerArray;
		addr_width: in natural;  
		data_width: in natural;
		index: out integer; 
		n_cols: out natural;
		extra_cols: out integer);

	-- return the cut that fills the maximum percentage of the
	-- area (with tie break advantage to row filling).
	-- returns a vector of length 3.
	--       index of cut (-1 if not found)
	--       addr_width of cut
        --       data_width of cut
	--       number of rows of cut
	--       number of columns of cut.
        function find_best_cut 
		(constant cut_address_widths: IntegerArray;
		    constant cut_data_widths: IntegerArray;
		    constant cut_row_heights: IntegerArray;
		    addr_width: in natural;  
		    data_width: in natural) return IntegerArray;

	function find_n_cols (constant cut_address_widths: IntegerArray;
		constant cut_data_widths: IntegerArray;
		constant cut_row_heights: IntegerArray;
		addr_width: natural;
		data_width: natural) return IntegerArray;

	--function Ceil_Log2(constant x : integer) return integer;
	function find_data_width (constant cut_data_widths: IntegerArray; 
		constant n_cols: Integerarray) return integer;
	function col_index (constant cut_data_widths: IntegerArray; 
		constant x: IntegerArray; index: integer) return integer;
	function MemDecoder(x: std_logic_vector) return std_logic_vector;
end package;

package body MemCutsPackage is

  -- Procedure: Min_array
  -- Description: Finds the minimum element (min) and it's position(index)
  -- 	in the given input array x, provided the element at the corresponding 
  -- 	position in the input array y is greater than 50.
  -- Inputs:
  -- 	x: array containing the number of replications of each cut
  --	y: array containing the utilization of each cut
  -- Outputs:
  -- 	min: minimum number of cuts having the cut utilization > 50%
  --	index: index of the minimum element in the input array x

  procedure Min_array(x: in IntegerArray;
		    y: in IntegerArray; 
		    min: out integer;
		    index: out integer ) is 
	alias lx:IntegerArray(1 to x'length) is x;
	alias ly:IntegerArray(1 to y'length) is y;
	variable min_var: integer;
	variable loc: integer;
  begin
	min_var := lx(1);
	loc := 1;
	for i in lx'length to 1 loop
		if (ly(i) > 50) then
			min_var := lx(i);
			loc := i;
		end if;
	end loop;
	
	for i in 1 to lx'length loop
		if (lx(i) < min_var) then
			if (ly(i) > 50) then
				min_var := lx(i);
				loc := i;
			end if;
		end if;
	end loop;

	min := min_var;
	index := loc;
  end Min_array; 
	    
  -- Procedure: opt_find
  -- Description: Covers the required MxN array with the smallest number 
  -- 	of column-replications subject to column utilization being at least 50%.
  -- Inputs:
  --	cut_address_widths: array of number of address lines of available cuts
  --	cut_data_widths: array of number of data lines of available cuts
  --	cut_row_heights: array of row heights of available cuts 
  -- 	addr_width: address width of the required MxN array
  -- 	data_width: data width of the required MxN array  
  -- Outputs:
  -- 	index: index of cut in 'cut_data_widths' using which minimum 
  -- 		column-replications are required to maximally cover N 
  -- 	n_cols: required number of column-replications of the optimal cut
  -- 	extra_cols: number of columns left after filling the N with optimal
  -- 		column-replications
	
  procedure opt_find (constant cut_address_widths: IntegerArray;
		constant cut_data_widths: IntegerArray;
		constant cut_row_heights: IntegerArray;
		addr_width: in natural;  
		data_width: in natural;
		index: out integer; 
		n_cols: out natural;
		extra_cols: out integer) is
	
	variable n_row_array, n_col_array, extra_col_array, n_cuts_array: IntegerArray(1 to cut_address_widths'length):= (others => 0);
	variable location, n_col: integer;
	variable Util_array: IntegerArray(1 to cut_address_widths'length);
  begin 
	for i in 1 to cut_address_widths'length loop

		if (data_width/cut_data_widths(i) = 0) then -- when data width is 
							    -- less than the cut width
			n_col_array(i) := 1;	
		-- when data width is integer multiples of cut width
		elsif (data_width/cut_data_widths(i) = 
			Ceiling (data_width, cut_data_widths(i))) then
			n_col_array(i) := data_width/cut_data_widths(i);		
		else
			n_col_array(i) := Ceiling(data_width, cut_data_widths(i))-1;
			extra_col_array(i) := data_width-n_col_array(i)*cut_data_widths(i);
		end if;

		n_row_array(i) := 2**(Maximum(0, addr_width-cut_address_widths(i)));
		Util_array(i) := 2**(addr_width)*data_width*100/
		(n_row_array(i)*cut_row_heights(i)*n_col_array(i)*cut_data_widths(i));	
		n_cuts_array(i) := n_row_array(i)*n_col_array(i);
	end loop;
	
	Min_array(n_cuts_array, Util_array, n_col, location);
	n_cols := n_col_array(location);
	index := location;	
	extra_cols := extra_col_array(location);
	
  end opt_find;
	
	-- return the cut that fills the maximum percentage of the
	-- area (with tie break advantage to row filling).
	-- returns a vector of length 3.
	--       index of cut (-1 if not found)
	--       addr_width of cut
        --       data_width of cut
	--       number of rows of cut
   function find_best_cut 
		(constant cut_address_widths: IntegerArray;
		    constant cut_data_widths: IntegerArray;
		    constant cut_row_heights: IntegerArray;
		    addr_width: in natural;  
		    data_width: in natural) return IntegerArray is
	variable a, r, s: natural;
	variable best_area, best_data_width, best_addr_width: natural;
	variable best_index: integer;
	variable ret_var: IntegerArray(1 to 5);
  begin

	s := ((2**addr_width) * data_width);
	ret_var := (others => 0);

	best_area := 0;
	best_data_width := 0;
 	best_addr_width := 0;
        best_index := -1;

        for  I in 1 to cut_address_widths'length loop
                a := (cut_row_heights(I) * cut_data_widths(I));
		if (a <= s) and  (cut_data_widths(I) <= data_width) and (cut_address_widths(I) <= addr_width)
			and ((a > best_area) or ((a = best_area) and (cut_data_widths(I) > best_data_width))) then
		   best_index := I;
		   best_area  := a;
                   best_data_width  := cut_data_widths(I);
		   best_addr_width := cut_address_widths(I);
		end if;
	end loop;

	ret_var(1) := best_index;
	if(best_index > 0) then
	   ret_var(2) := best_addr_width;
           ret_var(3) := best_data_width;
	   ret_var(4) := (2 ** (addr_width - best_addr_width));
	   ret_var(5) := (data_width/best_data_width);
        end if;

	return ret_var;
  end find_best_cut;

  -- function: find_n_cols
  -- Description: Finds the number of columns of each cut required to completely
  -- 		fill the data_width of the required MxN array
  -- Inputs:
  --	cut_address_widths: array of number of address lines of available cuts
  --	cut_data_widths: array of number of data lines of available cuts
  --	cut_row_heights: array of row heights of available cuts 
  -- 	addr_width: address width of the array to be build
  -- 	data_width: data width of the array to be build
  -- Output: 
  -- 	Array containing the required number of columns of availble cuts 
  
  function find_n_cols (constant cut_address_widths: IntegerArray;
		constant cut_data_widths: IntegerArray;
		constant cut_row_heights: IntegerArray;
		addr_width: natural;
		data_width: natural) return IntegerArray is

	variable n_col, additional_col: integer := 1;
	variable n_cols_array : IntegerArray(1 to cut_address_widths'length) := (others => 0);
	variable  empty_cols, index : integer := 1;
  begin
	empty_cols := data_width;
	while (additional_col /= 0) loop
		opt_find(cut_address_widths, cut_data_widths, cut_row_heights, 
		addr_width, empty_cols, index, n_col, additional_col);

		empty_cols := additional_col;
		n_cols_array(index) := n_cols_array(index) + n_col;
	end loop;
	
	return n_cols_array;
  end find_n_cols;

  -- function: Ceil_Log2
  -- Description: Calculates the ceiling of log to the base 2 of given integer x

  --function Ceil_Log2( constant x : integer) return integer is
	--variable ret_var : integer;
  --begin
    --ret_var := 0;
    --if(x > 1) then
      --while((2**ret_var) < x) loop
        --ret_var := ret_var + 1;
      --end loop;
    --end if;
    --return(ret_var);
  --end Ceil_Log2;


  -- function: find_data_width
  -- Description: Finds the resized data width of required memory cut
  -- Input:
  --	cut_data_widths: array of number of data lines of available cuts
  --	n_cols: array containing the number of columns of a available cuts
  --	   used to form the required MxN array
  -- Output:
  --	Sum of product of number of columns and cut data width of the
  -- 	available cuts

  function find_data_width (constant cut_data_widths: IntegerArray; 
	constant n_cols: Integerarray) return integer is 
	
	variable partial_prod: integer := 0;
  begin
	for i in 1 to cut_data_widths'length loop
		partial_prod := partial_prod + n_cols(i) * cut_data_widths(i);
	end loop;
	
	return(partial_prod);
  end function;


  -- function: col_index
  -- Description: Parts of N of MxN array are mapped to different cuts.
  -- 	To find out which part of N is mapped to a particular cut, index
  --	offset occured to due instantation of previous columns is to be known.
  -- 	This function returns the offset to be added to the resized_data's index 
  -- 	when generating a new column. 
  -- Inputs: 
  --	cut_data_widths: array of number of data lines of available cuts
  -- 	x: array containing the required number of columns of a available cuts  
  --	index: present index in the mem_gen instantiation loop

  function col_index (constant cut_data_widths: IntegerArray; 
	constant x: IntegerArray; index: integer) return integer is
	
	variable output: integer:=0;
  begin
		for i in 1 to index loop
			output := output + x(i)*cut_data_widths(i);
		end loop;
	
	return (output);		
  end function;
	
  -- function: MemDecoder
  -- Description: An n:2^n decoder  
  -- Input: n-bit vector x
  -- Output: 2^n-bit vector whose one of the bit = 0 that represents the given 
  -- input x, other output bits = 1

  function MemDecoder(x: std_logic_vector) return std_logic_vector is
	alias lx: std_logic_vector(x'length-1 downto 0) is x;
	variable ret_var: std_logic_vector((2**x'length)-1 downto 0);
	variable I : integer range 0 to (2**x'length)-1;
  begin
	ret_var := (others => '1');
	I := to_integer(to_unsigned(lx));
	ret_var(I) := '0';
	return(ret_var);
  end MemDecoder;

end package body;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.utilities.all;
--
-- dual port synchronous memory.. implemented with registers..
--
entity base_bank_dual_port_with_registers is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity base_bank_dual_port_with_registers;


architecture PlainRegisters of base_bank_dual_port_with_registers is
  type MemArray is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);
  signal mem_array : MemArray((2**g_addr_width)-1 downto 0) := (others => (others => '0'));
begin  -- PlainRegisters

  assert false report "DP MEMFF " & Convert_To_String ( g_data_width*(2**g_addr_width)) 
		severity note;
  --
  -- try to flag read/write clash!
  --
  process(clk, enable_0, enable_1, addrin_0, addrin_1) 
  begin
	if(clk'event and clk = '1') then
		if((enable_0 = '1') and (enable_1 = '1') and (addrin_0 = addrin_1) and
			(writebar_0 /= writebar_1)) then
			assert false report
				"Read and Write port clash in base_bank_dual_port " & name 
					severity error;
		end if;
	end if;
  end process; 

  -- read/write process
  process(clk, addrin_0,enable_0,writebar_0, addrin_1,enable_1,writebar_1)
  begin

    -- synch read-write memory
    if(clk'event and clk ='1') then

     if(reset = '1') then
	dataout_0 <= (others => '0');
	dataout_1 <= (others => '0');
     else
      	if(enable_0 = '1') then 
		if  (writebar_0 = '0') then
        		mem_array(To_Integer(unsigned(addrin_0))) <= datain_0;
		else
        		dataout_0 <= mem_array(To_Integer(unsigned(addrin_0)));
		end if;
      	end if;
      	if(enable_1 = '1') then
		if (writebar_1 = '0') then
        		mem_array(To_Integer(unsigned(addrin_1))) <= datain_1;
		else
        		dataout_1 <= mem_array(To_Integer(unsigned(addrin_1)));
		end if;
      	end if;
     end if;
    end if;
  end process;

end PlainRegisters;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.utilities.all;

-- memory implemented with registers..
entity base_bank_with_registers is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity base_bank_with_registers;


architecture PlainRegisters of base_bank_with_registers is
  type MemArray is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);
  signal mem_array : MemArray((2**g_addr_width)-1 downto 0) := (others => (others => '0'));
  signal read_data : std_logic_vector(g_data_width-1 downto 0);

begin  -- PlainRegisters

  assert false report "SP MEMFF " & Convert_To_String ( g_data_width*(2**g_addr_width)) 
		severity note;

  -- read/write process
  process(clk,addrin,enable,writebar)
  begin
    -- synch read-write memory
    if(clk'event and clk ='1') then
	if (reset = '1') then 
  		read_data <= (others => '0');
	elsif(enable = '1') then
		if(writebar = '0') then
        		mem_array(To_Integer(unsigned(addrin))) <= datain;
		else
  			read_data <= mem_array(To_Integer(unsigned(addrin)));
		end if;
	end if;
    end if;
  end process;
  dataout <= read_data;
end PlainRegisters;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;


-- a dummy ROM  which is never initialized.
-- any load to it returns 0.
entity dummy_read_only_memory_subsystem is
  generic(name: string;
	  num_loads             : natural := 5;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity dummy_read_only_memory_subsystem;


architecture Default_arch of dummy_read_only_memory_subsystem is
begin

     gen: for I in 0 to num_loads-1 generate
	lr_ack_out(I) <= lr_req_in(I);

	fsm: block
		signal busy : std_logic;
	begin
		lc_ack_out(I) <= busy;

		process(clock)
		begin
			if(clock'event and clock = '1') then
				if(reset = '1') then 
					busy <= '0';
				elsif (lr_req_in(I) = '1') then
					busy <= '1';
					lc_tag_out(((I+1)*tag_width)-1 downto (I*tag_width)) <= 
						lr_tag_in(((I+1)*tag_width)-1 downto (I*tag_width));
				elsif (lc_req_in(I) = '1') then
					busy <= '0';
				end if;
			end if;
		end process;
	end block;
     end generate gen;

end Default_arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

-- a dummy write-only memory (perfectly useless,
-- but plug-in for corner cases).
entity dummy_write_only_memory_subsystem is
  generic(name: string;
	  num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7);
  port(
    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity dummy_write_only_memory_subsystem;


-- architecture: synchronous R/W.
--               on destination conflict, writer with lowest index wins.
architecture Default_arch of dummy_write_only_memory_subsystem is
begin


     gen: for I in 0 to num_stores-1 generate
	sr_ack_out(I) <= sr_req_in(I);

	fsm: block
		signal busy : std_logic;
	begin
		sc_ack_out(I) <= busy;

		process(clock)
		begin
			if(clock'event and clock = '1') then
				if(reset = '1') then 
					busy <= '0';
				elsif (sr_req_in(I) = '1') then
					busy <= '1';
					sc_tag_out(((I+1)*tag_width)-1 downto I*tag_width) <= 
						sr_tag_in(((I+1)*tag_width)-1 downto I*tag_width);
				elsif (sc_req_in(I) = '1') then
					busy <= '0';
				end if;
			end if;
		end process;
	end block;
     end generate gen;

end Default_arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--
-- dual port synchronous memory.. implemented with registers..
--  with asynchronous read.
--
entity fifo_mem_synch_write_asynch_read is
   generic ( name: string; address_width: natural;  
			data_width : natural;
				mem_size: natural);
   port (
	 write_enable: in std_logic;
	 write_data: in std_logic_vector(data_width-1 downto 0);
	 write_address: in std_logic_vector(address_width-1 downto 0);
	 read_data: out std_logic_vector(data_width-1 downto 0);
	 read_address: in std_logic_vector(address_width-1 downto 0);
         clk: in std_logic);
end entity fifo_mem_synch_write_asynch_read;


architecture PlainRegisters of fifo_mem_synch_write_asynch_read is
  type MemArray is array (natural range <>) of std_logic_vector(data_width-1 downto 0);
  signal mem_array : MemArray(mem_size-1 downto 0);
begin  -- PlainRegisters

	process(clk, write_address, read_address, mem_array)
		variable wr_addr_var, rd_addr_var : integer;
		variable wr_ok: boolean;
	begin

		wr_addr_var := To_Integer(unsigned(write_address));
		wr_ok := (wr_addr_var < mem_size);

		if(clk'event and clk = '1') then

			if (wr_ok and (write_enable = '1')) then
        			mem_array(wr_addr_var) <= write_data;
			end if;

		end if;
	
		read_data <= mem_array(To_Integer(unsigned(read_address)));
	end process;

end PlainRegisters;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.mem_function_pack.all;
use ahir.mem_component_pack.all;

entity memory_bank_base is
   generic ( name: string;
	g_addr_width: natural; 
	g_data_width : natural;
        g_base_bank_addr_width: natural;
        g_base_bank_data_width: natural);
   port (data_in : in std_logic_vector(g_data_width-1 downto 0);
         data_out: out std_logic_vector(g_data_width-1 downto 0);
         addr_in: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         write_bar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity memory_bank_base;


architecture structural of memory_bank_base is
  constant bank_array_width : natural := Ceiling(g_data_width,g_base_bank_data_width);
  constant bank_array_height : natural := 2**(Maximum(0,g_addr_width-g_base_bank_addr_width));

  type BankArrayDataArray is array (0 to bank_array_height-1, 0 to bank_array_width -1) of std_logic_vector(g_base_bank_data_width-1 downto 0);
  signal data_in_array, data_out_array : BankArrayDataArray;
  

  type BankArrayControlArray is array (0 to bank_array_height-1, 0 to bank_array_width -1) of std_logic;
  signal enable_array,enable_array_reg: BankArrayControlArray;
  
  signal padded_data_in,padded_data_out : std_logic_vector(bank_array_width*g_base_bank_data_width -1 downto 0);
  signal base_addr_in : std_logic_vector(g_base_bank_addr_width -1 downto 0);
  
  signal write_bar_reg: std_logic;
begin  -- structural

   -- register write_bar_reg because memory read will finish after one clock.
    process(clk,reset)
    begin
        if(clk'event and clk = '1') then
		if(reset = '1') then
			write_bar_reg <= '0';
		else
			write_bar_reg <= write_bar;
		end if;
	end if;
    end process;

process(addr_in)
        constant l_index: natural := Minimum(g_addr_width-1, g_base_bank_addr_width-1);
    begin
        base_addr_in <= (others => '0');
        base_addr_in(l_index downto 0) <= addr_in(l_index downto 0);
    end process;
    
process(data_in)
    begin
        padded_data_in <= (others => '0');
        padded_data_in(g_data_width-1 downto 0) <= data_in;
    end process;
    
  data_out <= padded_data_out(g_data_width-1 downto 0);

  -- pack/unpack
  ColGen: for COL in 0 to bank_array_width-1 generate
    
    RowGen: for ROW in 0 to bank_array_height-1 generate
      process(addr_in, enable)
      begin
        enable_array(ROW,COL) <= '0';
        if(bank_array_height > 1) then
          if(enable = '1') then
            if(ROW = To_Integer(addr_in(g_addr_width - 1 downto g_base_bank_addr_width))) then
              enable_array(ROW,COL) <= '1';
            end if;
          end if;
        else
          enable_array(ROW,COL) <= enable;
        end if;
      end process;

      process(clk,reset)
      begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			enable_array_reg(ROW,COL) <= '0';
		else
			enable_array_reg(ROW,COL) <= enable_array(ROW,COL);
		end if;
	end if;
      end process;

      process(padded_data_in)
      begin
        data_in_array(ROW,COL) <= padded_data_in((COL+1)*g_base_bank_data_width - 1 downto COL*g_base_bank_data_width);
      end process;

      baseMem : base_bank generic map (
        name => name & "-baseMem", 
        g_addr_width => g_base_bank_addr_width,
        g_data_width => g_base_bank_data_width)
        port map (
          datain => data_in_array(ROW, COL),
          addrin => base_addr_in,
          enable => enable_array(ROW,COL),
          writebar => write_bar,
          dataout => data_out_array(ROW,COL),
          clk => clk,
          reset => reset);
      
    end generate RowGen;
    
    process(data_out_array,enable_array_reg, write_bar_reg)
    begin
      padded_data_out((COL+1)*g_base_bank_data_width -1 downto (COL*g_base_bank_data_width)) <= (others => '0');
      for ROW in 0 to bank_array_height-1 loop
	-- use delayed version of enable and write_bar to pass read data
        if(enable_array_reg(ROW,COL) = '1' and write_bar_reg = '1') then
          padded_data_out((COL+1)*g_base_bank_data_width -1 downto (COL*g_base_bank_data_width)) <= data_out_array(ROW,COL);
        end if;
      end loop;  -- ROW
    end process;
    
  end generate ColGen;

end structural;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.mem_function_pack.all;
use ahir.mem_component_pack.all;

entity memory_bank_revised is
   generic (
     name: string;
     g_addr_width: natural;
     g_data_width: natural;
     g_write_tag_width : natural;
     g_write_port_id_width : natural;
     g_read_tag_width : natural;
     g_read_port_id_width : natural;
     g_time_stamp_width: natural;
     g_base_bank_addr_width: natural;
     g_base_bank_data_width: natural
	);
   port (
     clk : in std_logic;
     reset: in std_logic;
     write_data     : in  std_logic_vector(g_data_width-1 downto 0);
     write_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     write_tag      : in std_logic_vector(g_write_tag_width-1 downto 0);
     write_time_stamp: in std_logic_vector(g_time_stamp_width-1 downto 0);
     write_tag_out  : out std_logic_vector(g_write_tag_width-1 downto 0);
     write_port_id      : in unsigned(g_write_port_id_width-1 downto 0);
     write_port_id_out  : out unsigned(g_write_port_id_width-1 downto 0);
     write_enable   : in std_logic;
     write_ack   : out std_logic;
     write_result_accept : in std_logic;
     write_result_ready : out std_logic;
     read_data     : out std_logic_vector(g_data_width-1 downto 0);
     read_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     read_tag      : in std_logic_vector(g_read_tag_width-1 downto 0);
     read_time_stamp: in std_logic_vector(g_time_stamp_width-1 downto 0);
     read_tag_out  : out std_logic_vector(g_read_tag_width-1 downto 0);
     read_port_id      : in unsigned(g_read_port_id_width-1 downto 0);
     read_port_id_out  : out unsigned(g_read_port_id_width-1 downto 0);
     read_enable   : in std_logic;
     read_ack      : out std_logic;
     read_result_accept: in std_logic;
     read_result_ready: out std_logic
     );
end entity memory_bank_revised;


architecture SimModel of memory_bank_revised is

  signal write_has_priority: std_logic;
  signal enable_base,enable_sig, write_enable_base, read_enable_base, read_enable_base_registered: std_logic;

  signal addr_base : std_logic_vector(g_addr_width-1 downto 0);
  signal read_data_base  : std_logic_vector(g_data_width-1 downto 0);
  signal read_data_base_reg  : std_logic_vector(g_data_width-1 downto 0);
  
  type FsmState is (IDLE, RDONE, WDONE);
  signal fsm_state : FsmState;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- behave

  Tstampgen: if g_time_stamp_width > 0 generate 
  
  tstamp_block: Block
  begin 
  	process(read_time_stamp,write_time_stamp, read_enable, write_enable)
  	begin
      	if(write_enable = '1' and read_enable = '1') then
		if(IsGreaterThan(write_time_stamp,read_time_stamp)) then
        		write_has_priority <=   '0';
		else
			write_has_priority <= '1';
		end if;
      	elsif(write_enable = '1') then
		write_has_priority <= '1';
      	elsif(read_enable = '1') then
		write_has_priority <= '0';
      	else
		write_has_priority <= '1';
      	end if;
  	end process;
   end block;
   end generate Tstampgen;

   NoTstampGen: if g_time_stamp_width <= 0 generate
        write_has_priority <= write_enable;
   end generate NoTstampGen;

  -- FSM
  process(clk, reset, fsm_state, 
		write_enable, write_addr, write_data, write_result_accept, write_has_priority,
		read_enable, read_addr, read_result_accept)
	variable next_state: FsmState;
	variable we_base, re_base: std_logic;
        variable wrr, rrr: std_logic;

	variable write_active, read_active: boolean;
  begin
	next_state := fsm_state;
	we_base := '0'; 
	re_base := '0';
	wrr	:= '0';
	rrr 	:= '0';

	write_active := ((((write_enable = '1') and (read_enable = '1')) and (write_has_priority = '1'))
				or
			 ((write_enable = '1') and (read_enable = '0')));
	read_active := ((((write_enable = '1') and (read_enable = '1')) and (write_has_priority = '0'))
				or
			 ((write_enable = '0') and (read_enable = '1')));

	case fsm_state is
		when IDLE =>
		        if(write_active) then
				we_base := '1';
				next_state := WDONE;
			elsif (read_active) then
				re_base := '1';
				next_state := RDONE;
			end if;
		when RDONE =>
			rrr := '1';
			if(read_result_accept = '1') then
		        	if(write_active) then
					we_base := '1';
					next_state := WDONE;
				elsif (read_active) then
					re_base := '1';
					next_state := RDONE;
				else
					next_state := IDLE;
				end if;
			end if;
		when WDONE =>
			wrr := '1';
			if(write_result_accept ='1') then
		        	if(write_active) then
					we_base := '1';
					next_state := WDONE;
				elsif (read_active) then
					re_base := '1';
					next_state := RDONE;
				else
					next_state := IDLE;
				end if;
			end if;
	end case;

	write_enable_base <= we_base;
	write_ack <= we_base;

	read_enable_base <= re_base;
	read_ack <= re_base;

	write_result_ready <= wrr;
	read_result_ready <= rrr;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			fsm_state <= IDLE;
			read_enable_base_registered <= '0';
		else
			fsm_state <= next_state;
			read_enable_base_registered <= re_base;
		end if;
	end if;
  end process;

  addr_base <= write_addr when write_enable_base = '1' else read_addr when read_enable_base = '1' else (others => '0');
  enable_sig <= write_enable_base or read_enable_base;
  
  memBase: memory_bank_base generic map(name => name & "-memBase", g_addr_width => g_addr_width,
                                        g_data_width => g_data_width,
					g_base_bank_addr_width => g_base_bank_addr_width,
					g_base_bank_data_width => g_base_bank_data_width)
    port map(data_in => write_data,
             addr_in => addr_base,
             data_out => read_data_base,
             enable => enable_sig,
             write_bar => read_enable_base,
             clk => clk,
             reset => reset);
 

  -- tag-out is updated in parallel with the
  -- memory access in memory_bank_base.
  process(clk)
  begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
		     read_tag_out <= (others => '0');
		     read_port_id_out <= (others => '0');

		     write_tag_out <= (others => '0');
		     write_port_id_out <= (others => '0');
		elsif(enable_sig = '1') then
			if(read_enable_base = '1') then
				read_tag_out <= read_tag;
				read_port_id_out <= read_port_id;
			else
				write_tag_out <= write_tag;
				write_port_id_out <= write_port_id;
			end if;
		end if;
	end if;
  end process;

  -- bypass register for read_data_base
  process(clk)
  begin
	if(clk'event and clk = '1') then
		if(read_enable_base_registered = '1') then 
			read_data_base_reg  <= read_data_base;
		end if;
	end if;
  end process;
  read_data <= read_data_base when (read_enable_base_registered = '1') else read_data_base_reg;

end SimModel;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.mem_function_pack.all;
use ahir.mem_component_pack.all;

entity memory_bank is
   generic (
     name: string;
     g_addr_width: natural;
     g_data_width: natural;
     g_write_tag_width : natural;
     g_read_tag_width : natural;
     g_time_stamp_width: natural;
     g_base_bank_addr_width: natural;
     g_base_bank_data_width: natural
	);
   port (
     clk : in std_logic;
     reset: in std_logic;
     write_data     : in  std_logic_vector(g_data_width-1 downto 0);
     write_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     write_tag      : in std_logic_vector(g_write_tag_width-1 downto 0);
     write_tag_out  : out std_logic_vector(g_write_tag_width-1 downto 0);
     write_enable   : in std_logic;
     write_ack   : out std_logic;
     write_result_accept : in std_logic;
     write_result_ready : out std_logic;
     read_data     : out std_logic_vector(g_data_width-1 downto 0);
     read_addr     : in std_logic_vector(g_addr_width-1 downto 0);
     read_tag      : in std_logic_vector(g_read_tag_width-1 downto 0);
     read_tag_out  : out std_logic_vector(g_read_tag_width-1 downto 0);
     read_enable   : in std_logic;
     read_ack      : out std_logic;
     read_result_accept: in std_logic;
     read_result_ready: out std_logic
     );
end entity memory_bank;


architecture SimModel of memory_bank is

  signal write_has_priority: std_logic;
  signal enable_base,enable_sig, write_enable_base, read_enable_base, read_enable_base_registered: std_logic;

  signal addr_base : std_logic_vector(g_addr_width-1 downto 0);
  signal read_data_base  : std_logic_vector(g_data_width-1 downto 0);
  signal read_data_base_reg  : std_logic_vector(g_data_width-1 downto 0);
  
  type FsmState is (IDLE, RDONE, WDONE);
  signal fsm_state : FsmState;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- behave

  Tstampgen: if g_time_stamp_width > 0 generate 
  
  tstamp_block: Block
  	signal read_time_stamp, write_time_stamp: std_logic_vector(g_time_stamp_width-1 downto 0);
  begin 
  	read_time_stamp <= read_tag(g_time_stamp_width-1 downto 0);
  	write_time_stamp <= write_tag(g_time_stamp_width-1 downto 0);

  	process(read_time_stamp,write_time_stamp, read_enable, write_enable)
  	begin
      	if(write_enable = '1' and read_enable = '1') then
		if(IsGreaterThan(write_time_stamp,read_time_stamp)) then
        		write_has_priority <=   '0';
		else
			write_has_priority <= '1';
		end if;
      	elsif(write_enable = '1') then
		write_has_priority <= '1';
      	elsif(read_enable = '1') then
		write_has_priority <= '0';
      	else
		write_has_priority <= '1';
      	end if;
  	end process;
   end block;
   end generate Tstampgen;

   NoTstampGen: if g_time_stamp_width <= 0 generate
        write_has_priority <= write_enable;
   end generate NoTstampGen;

  -- FSM
  process(clk, reset, fsm_state, 
		write_enable, write_addr, write_data, write_result_accept, write_has_priority,
		read_enable, read_addr, read_result_accept)
	variable next_state: FsmState;
	variable we_base, re_base: std_logic;
        variable wrr, rrr: std_logic;

	variable write_active, read_active: boolean;
  begin
	next_state := fsm_state;
	we_base := '0'; 
	re_base := '0';
	wrr	:= '0';
	rrr 	:= '0';

	write_active := ((((write_enable = '1') and (read_enable = '1')) and (write_has_priority = '1'))
				or
			 ((write_enable = '1') and (read_enable = '0')));
	read_active := ((((write_enable = '1') and (read_enable = '1')) and (write_has_priority = '0'))
				or
			 ((write_enable = '0') and (read_enable = '1')));

	case fsm_state is
		when IDLE =>
		        if(write_active) then
				we_base := '1';
				next_state := WDONE;
			elsif (read_active) then
				re_base := '1';
				next_state := RDONE;
			end if;
		when RDONE =>
			rrr := '1';
			if(read_result_accept = '1') then
		        	if(write_active) then
					we_base := '1';
					next_state := WDONE;
				elsif (read_active) then
					re_base := '1';
					next_state := RDONE;
				else
					next_state := IDLE;
				end if;
			end if;
		when WDONE =>
			wrr := '1';
			if(write_result_accept ='1') then
		        	if(write_active) then
					we_base := '1';
					next_state := WDONE;
				elsif (read_active) then
					re_base := '1';
					next_state := RDONE;
				else
					next_state := IDLE;
				end if;
			end if;
	end case;

	write_enable_base <= we_base;
	write_ack <= we_base;

	read_enable_base <= re_base;
	read_ack <= re_base;

	write_result_ready <= wrr;
	read_result_ready <= rrr;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			fsm_state <= IDLE;
			read_enable_base_registered <= '0';
		else
			fsm_state <= next_state;
			read_enable_base_registered <= re_base;
		end if;
	end if;
  end process;

  addr_base <= write_addr when write_enable_base = '1' else read_addr when read_enable_base = '1' else (others => '0');
  enable_sig <= write_enable_base or read_enable_base;
  
  memBase: memory_bank_base generic map(name => name & "-memBase", g_addr_width => g_addr_width,
                                        g_data_width => g_data_width,
					g_base_bank_addr_width => g_base_bank_addr_width,
					g_base_bank_data_width => g_base_bank_data_width)
    port map(data_in => write_data,
             addr_in => addr_base,
             data_out => read_data_base,
             enable => enable_sig,
             write_bar => read_enable_base,
             clk => clk,
             reset => reset);
 

  -- tag-out is updated in parallel with the
  -- memory access in memory_bank_base.
  process(clk)
  begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
		     read_tag_out <= (others => '0');
		     write_tag_out <= (others => '0');
		elsif(enable_sig = '1') then
			if(read_enable_base = '1') then
				read_tag_out <= read_tag;
			else
				write_tag_out <= write_tag;
			end if;
		end if;
	end if;
  end process;

  -- bypass register for read_data_base
  process(clk)
  begin
	if(clk'event and clk = '1') then
		if(read_enable_base_registered = '1') then 
			read_data_base_reg  <= read_data_base;
		end if;
	end if;
  end process;
  read_data <= read_data_base when (read_enable_base_registered = '1') else read_data_base_reg;

end SimModel;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

-- effectively a two entry queue.
-- used to break combinational paths
-- at the cost of a single cycle delay from input
-- to output.
entity mem_repeater is
    generic(name: string; g_data_width: integer := 32);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(g_data_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector(g_data_width-1 downto 0);
       req_out : out std_logic;
       ack_in: in std_logic);
end entity mem_repeater;

architecture behave of mem_repeater is
begin  -- SimModel

  bqueue: QueueBase
             generic map (name => name & ":bqueue", queue_depth => 2,  data_width => g_data_width,
				save_one_slot => false)
	     port map (clk => clk, reset => reset, 
       				data_in => data_in,
       				push_req => req_in,
       				push_ack => ack_out,
       				data_out => data_out,
       				pop_ack => req_out,
				pop_req => ack_in);
end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;
use ahir.mem_function_pack.all;

entity mem_shift_repeater is
    generic(name: string; g_data_width: integer := 32; g_number_of_stages: natural := 16);
    port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(g_data_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector(g_data_width-1 downto 0);
       req_out : out std_logic;
       ack_in: in std_logic);
end entity mem_shift_repeater;

architecture behave of mem_shift_repeater is

  type DataArray is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);
  signal idata : DataArray(0 to g_number_of_stages);
  signal ireq,iack : std_logic_vector(0 to g_number_of_stages);

begin  -- SimModel

  idata(0) <= data_in;
  ireq(0)  <= req_in;
  ack_out <= iack(0);

  data_out <= idata(g_number_of_stages);
  req_out <= ireq(g_number_of_stages);
  iack(g_number_of_stages) <= ack_in;

  ifGen: if g_number_of_stages > 0 generate

    RepGen: for I in 0 to g_number_of_stages-1 generate
      rptr : mem_repeater generic map (
	name => name & "-RepGen-rptr-" & Convert_Integer_To_String(I),
        g_data_width => g_data_width)
        port map (
          clk      => clk,
          reset    => reset,
          data_in  => idata(I),
          req_in   => ireq(I),
          ack_out  => iack(I),
          data_out => idata(I+1),
          req_out  => ireq(I+1),
          ack_in   => iack(I+1));
    end generate RepGen;
  end generate ifGen; 

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.utilities.all;

--
-- 1 read/1-write port synchronous memory.. implemented with registers..
--
entity register_file_1w_1r_port_with_registers  is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity register_file_1w_1r_port_with_registers ;


architecture PlainRegisters of register_file_1w_1r_port_with_registers  is
  type MemArray is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);
  signal mem_array : MemArray((2**g_addr_width)-1 downto 0) := (others => (others => '0'));
begin  -- PlainRegisters

  assert false report "1W1R MEMFF " & Convert_To_String ( g_data_width*(2**g_addr_width)) 
		severity note;

  -- read/write process
  process(clk, addrin_0,enable_0,addrin_1,enable_1)
  begin

    -- synch read-write memory
    if(clk'event and clk ='1') then

     if(reset = '1') then
	dataout_1 <= (others => '0');
     else
      	if(enable_0 = '1') then 
        	mem_array(To_Integer(unsigned(addrin_0))) <= datain_0;
      	end if;
      	if(enable_1 = '1') then
        	dataout_1 <= mem_array(To_Integer(unsigned(addrin_1)));
      	end if;
     end if;
    end if;

  end process;

end PlainRegisters;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.types.all;
use ahir.utilities.all;

package mem_ASIC_components is

  component DPRAM_32X8 is
   port(       QA,QB : out std_logic_vector(7 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(4 downto 0) := TieHighSlvConstant(5);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component DPRAM_256X32 is
   port(       QA,QB : out std_logic_vector(31 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(31 downto 0) := TieHighSlvConstant(32);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component DPRAM_2048X8 is
   port(       QA,QB : out std_logic_vector(7 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(10 downto 0) := TieHighSlvConstant(11);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component DPRAM_2048X36 is
   port(       QA,QB : out std_logic_vector(35 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(10 downto 0) := TieHighSlvConstant(11);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(35 downto 0) := TieHighSlvConstant(36);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component DPRAM_256X52 is
   port(       QA,QB : out std_logic_vector(51 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(51 downto 0) := TieHighSlvConstant(52);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component DPRAM_32X64 is
   port(       QA,QB : out std_logic_vector(63 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(4 downto 0) := TieHighSlvConstant(5);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(63 downto 0) := TieHighSlvConstant(64);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component DPRAM_32X4 is
   port(       QA,QB : out std_logic_vector(3 downto 0);
      AA,AB,AMA,AMB : in std_logic_vector(4 downto 0) := TieHighSlvConstant(5);
      DA,DB,DMA,DMB,BWEBA,BWEBB,BWEBMA,BWEBMB : in std_logic_vector(3 downto 0) := TieHighSlvConstant(4);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD, VG, VS  :   IN   std_logic := '1'; --- ????? 
      BIST  :   IN   std_logic := '1'; --- ????? 
      AWT:   IN   std_logic := '1'; --- ????? 
      WTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      RTSEL  :   IN   std_logic_vector(1 downto 0) := "11"; --- ????? 
      CEBA, CEBB :   IN   std_logic := '1';
      CEBMA, CEBMB :   IN   std_logic := '1';
      WEBA, WEBB :   IN   std_logic := '1';
      WEBMA, WEBMB :   IN   std_logic := '1';
      CLKA, CLKB, CLKM  :   IN   std_logic := '1');
  end component;
  component SRAM_64X4 is
   port(       Q : out std_logic_vector(3 downto 0);
      A, AM : in std_logic_vector(5 downto 0) := TieHighSlvConstant(6);
      D, DM, BWEB, BWEBM : in std_logic_vector(3 downto 0) := TieHighSlvConstant(4);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_64X32 is
   port(       Q : out std_logic_vector(31 downto 0);
      A, AM : in std_logic_vector(5 downto 0) := TieHighSlvConstant(6);
      D, DM, BWEB, BWEBM : in std_logic_vector(31 downto 0) := TieHighSlvConstant(32);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_256X8 is
   port(       Q : out std_logic_vector(7 downto 0);
      A, AM : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      D, DM, BWEB, BWEBM : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_256X32 is
   port(       Q : out std_logic_vector(31 downto 0);
      A, AM : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      D, DM, BWEB, BWEBM : in std_logic_vector(31 downto 0) := TieHighSlvConstant(32);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_8192X8 is
   port(       Q : out std_logic_vector(7 downto 0);
      A, AM : in std_logic_vector(12 downto 0) := TieHighSlvConstant(13);
      D, DM, BWEB, BWEBM : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_32X32 is
   port(       Q : out std_logic_vector(31 downto 0);
      A, AM : in std_logic_vector(4 downto 0) := TieHighSlvConstant(5);
      D, DM, BWEB, BWEBM : in std_logic_vector(31 downto 0) := TieHighSlvConstant(32);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_128X22 is
   port(       Q : out std_logic_vector(21 downto 0);
      A, AM : in std_logic_vector(6 downto 0) := TieHighSlvConstant(7);
      D, DM, BWEB, BWEBM : in std_logic_vector(21 downto 0) := TieHighSlvConstant(22);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_1024X8 is
   port(       Q : out std_logic_vector(7 downto 0);
      A, AM : in std_logic_vector(9 downto 0) := TieHighSlvConstant(10);
      D, DM, BWEB, BWEBM : in std_logic_vector(7 downto 0) := TieHighSlvConstant(8);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_1024X64 is
   port(       Q : out std_logic_vector(63 downto 0);
      A, AM : in std_logic_vector(9 downto 0) := TieHighSlvConstant(10);
      D, DM, BWEB, BWEBM : in std_logic_vector(63 downto 0) := TieHighSlvConstant(64);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_64X128 is
   port(       Q : out std_logic_vector(127 downto 0);
      A, AM : in std_logic_vector(5 downto 0) := TieHighSlvConstant(6);
      D, DM, BWEB, BWEBM : in std_logic_vector(127 downto 0) := TieHighSlvConstant(128);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_64X67 is
   port(       Q : out std_logic_vector(66 downto 0);
      A, AM : in std_logic_vector(5 downto 0) := TieHighSlvConstant(6);
      D, DM, BWEB, BWEBM : in std_logic_vector(66 downto 0) := TieHighSlvConstant(67);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_64X24 is
   port(       Q : out std_logic_vector(23 downto 0);
      A, AM : in std_logic_vector(5 downto 0) := TieHighSlvConstant(6);
      D, DM, BWEB, BWEBM : in std_logic_vector(23 downto 0) := TieHighSlvConstant(24);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
  component SRAM_64X90 is
   port(       Q : out std_logic_vector(89 downto 0);
      A, AM : in std_logic_vector(5 downto 0) := TieHighSlvConstant(6);
      D, DM, BWEB, BWEBM : in std_logic_vector(89 downto 0) := TieHighSlvConstant(90);
      SLP  :   IN   std_logic := '1'; --- ????? 
      SD   :   IN   std_logic := '1'; --- ????? 
      WEB  :   IN   std_logic;
      CEB  :   IN   std_logic;
      WEBM : in std_logic := '1'; --- ????? 
      CEBM : in std_logic := '1'; --- ????? 
      AWT  : in std_logic := '1'; --- ????? 
      BIST : in std_logic := '1'; --- ????? 
      CLK:   IN   std_logic);
  end component;
end package;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;
--use ahir.Utilities.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

package MemcutDescriptionPackage is
   constant spmem_cut_row_heights : IntegerArray(1 to 13) := (64, 64, 64, 64, 1024, 1024, 128, 32, 8192, 256, 256, 64, 64);
    constant spmem_cut_address_widths : IntegerArray(1 to 13) := (6, 6, 6, 6, 10, 10, 7, 5, 13, 8, 8, 6, 6);
    constant spmem_cut_data_widths : IntegerArray(1 to 13) := (90, 24, 67, 128, 64, 8, 22, 32, 8, 32, 8, 32, 4);
   constant dpmem_cut_row_heights : IntegerArray(1 to 7) := (32, 32, 256, 2048, 2048, 256, 32);
    constant dpmem_cut_address_widths : IntegerArray(1 to 7) := (5, 5, 8, 11, 11, 8, 5);
    constant dpmem_cut_data_widths : IntegerArray(1 to 7) := (4, 64, 52, 36, 8, 32, 8);
   constant register_file_1w_1r_cut_row_heights : IntegerArray(1 to 7) := (32, 32, 256, 2048, 2048, 256, 32);
    constant register_file_1w_1r_cut_address_widths : IntegerArray(1 to 7) := (5, 5, 8, 11, 11, 8, 5);
    constant register_file_1w_1r_cut_data_widths : IntegerArray(1 to 7) := (4, 64, 52, 36, 8, 32, 8);
end package;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_ASIC_components.all;
use ahir.types.all;
use ahir.utilities.all;

-- Entity to instantiate different available memory cuts based on the 
-- address_width and data_width generics passed.
entity dpmem_selector is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		WRITE_0_BAR : in std_logic;
		WRITE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAIN_1  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_0  : out std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK, RESET: in std_logic);
end entity dpmem_selector;

architecture StructGen of dpmem_selector is
	signal TIE_HIGH, TIE_LOW: std_logic;
        signal TIE_LOW_2, TIE_HIGH_2: std_logic_vector(1 downto 0);
        signal TIE_LOW_3: std_logic_vector(2 downto 0);
        signal TIE_LOW_4: std_logic_vector(3 downto 0);
begin
	TIE_HIGH <= '1';
	TIE_LOW <= '0';
	TIE_LOW_2 <= (others => '0');
	TIE_HIGH_2 <= (others => '1');
	TIE_LOW_3 <= (others => '0');
	TIE_LOW_4 <= (others => '0');
  DPRAM_32X8_gen: if (address_width = 5) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_32X8
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_32X8_gen;
  DPRAM_256X32_gen: if (address_width = 8) and (data_width = 32) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(31 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(31 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(7 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_256X32
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_256X32_gen;
  DPRAM_2048X8_gen: if (address_width = 11) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(10 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(10 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_2048X8
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_2048X8_gen;
  DPRAM_2048X36_gen: if (address_width = 11) and (data_width = 36) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(35 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(35 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(10 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(10 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_2048X36
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_2048X36_gen;
  DPRAM_256X52_gen: if (address_width = 8) and (data_width = 52) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(51 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(51 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(7 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_256X52
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_256X52_gen;
  DPRAM_32X64_gen: if (address_width = 5) and (data_width = 64) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(63 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(63 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_32X64
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_32X64_gen;
  DPRAM_32X4_gen: if (address_width = 5) and (data_width = 4) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(3 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(3 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_32X4
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => WRITE_0_BAR, WEBB => WRITE_1_BAR, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATAIN_1, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => DATAOUT_0, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_32X4_gen;
end StructGen;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_ASIC_components.all;

-- Entity to instantiate different available memory cuts based on the 
-- address_width and data_width generics passed.
entity register_file_1w_1r_selector is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK, RESET: in std_logic);
end entity register_file_1w_1r_selector;

architecture StructGen of register_file_1w_1r_selector is
	signal TIE_HIGH, TIE_LOW: std_logic;
        signal TIE_LOW_2, TIE_HIGH_2: std_logic_vector(1 downto 0);
        signal TIE_LOW_3: std_logic_vector(2 downto 0);
        signal TIE_LOW_4: std_logic_vector(3 downto 0);
begin
	TIE_HIGH <= '1';
	TIE_LOW <= '0';
        TIE_LOW_2 <= (others => '0');
        TIE_HIGH_2 <= (others => '1');
	TIE_LOW_3 <= (others => '0');
	TIE_LOW_4 <= (others => '0');
  DPRAM_32X8_gen: if (address_width = 5) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_32X8
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_32X8_gen;
  DPRAM_256X32_gen: if (address_width = 8) and (data_width = 32) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(31 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(31 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(7 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_256X32
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_256X32_gen;
  DPRAM_2048X8_gen: if (address_width = 11) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(10 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(10 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_2048X8
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_2048X8_gen;
  DPRAM_2048X36_gen: if (address_width = 11) and (data_width = 36) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(35 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(35 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(10 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(10 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_2048X36
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_2048X36_gen;
  DPRAM_256X52_gen: if (address_width = 8) and (data_width = 52) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(51 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(51 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(7 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_256X52
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_256X52_gen;
  DPRAM_32X64_gen: if (address_width = 5) and (data_width = 64) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(63 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(63 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_32X64
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_32X64_gen;
  DPRAM_32X4_gen: if (address_width = 5) and (data_width = 4) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(3 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(3 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: DPRAM_32X4
   port map (AA => ADDR_0, AB => ADDR_1, CLKA => CLK, CLKB => CLK, WEBA => ENABLE_0_BAR, WEBB => TIE_HIGH, CEBA => ENABLE_0_BAR, CEBB => ENABLE_1_BAR,  DA => DATAIN_0, DB => DATA_TIE_LOW, BWEBA => DATA_TIE_LOW, BWEBB => DATA_TIE_LOW, QA => OPEN, QB => DATAOUT_1,  SLP => TIE_LOW, SD => TIE_LOW, VG => TIE_LOW, VS => TIE_LOW, AWT => TIE_LOW, CEBMA => TIE_HIGH, CEBMB => TIE_HIGH, WEBMA => TIE_HIGH, WEBMB => TIE_HIGH,  BWEBMA => DATA_TIE_HIGH, BWEBMB => DATA_TIE_HIGH, AMA => ADDR_TIE_HIGH,  AMB => ADDR_TIE_HIGH,  DMA => DATA_TIE_HIGH,  DMB => DATA_TIE_HIGH, BIST => TIE_LOW,  WTSEL => TIE_LOW_2,  RTSEL => TIE_LOW_2);
         end block;
  end generate DPRAM_32X4_gen;
end StructGen;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_ASIC_components.all;
use ahir.types.all;
use ahir.utilities.all;

-- Entity to instantiate different available memory cuts based on the 
-- address_width and data_width generics passed.
entity spmem_selector is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR : in std_logic_vector(address_width-1 downto 0 );
		CLK : in std_logic;
	        RESET: in std_logic;
		WRITE_BAR: in std_logic;
		ENABLE_BAR: in std_logic;
		DATAIN  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT  : out std_logic_vector(data_width-1 downto 0));
end entity spmem_selector;

architecture StructGen of spmem_selector is

  signal TIE_HIGH, TIE_LOW: std_logic;
  signal TIE_LOW_2, TIE_HIGH_2: std_logic_vector(1 downto 0);
  signal TIE_LOW_3: std_logic_vector(2 downto 0);
  signal TIE_LOW_4: std_logic_vector(3 downto 0);

begin
  
  TIE_HIGH <= '1';
  TIE_LOW  <= '0';
  TIE_LOW_2 <= (others => '0');
  TIE_HIGH_2 <= (others => '1');
  TIE_LOW_3 <= (others => '0');
  TIE_LOW_4 <= (others => '0');
  SRAM_64X4_gen: if (address_width = 6) and (data_width = 4) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(3 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(3 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(5 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(5 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_64X4
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_64X4_gen;
  SRAM_64X32_gen: if (address_width = 6) and (data_width = 32) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(31 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(31 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(5 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(5 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_64X32
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_64X32_gen;
  SRAM_256X8_gen: if (address_width = 8) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(7 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_256X8
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_256X8_gen;
  SRAM_256X32_gen: if (address_width = 8) and (data_width = 32) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(31 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(31 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(7 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_256X32
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_256X32_gen;
  SRAM_8192X8_gen: if (address_width = 13) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(12 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(12 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_8192X8
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_8192X8_gen;
  SRAM_32X32_gen: if (address_width = 5) and (data_width = 32) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(31 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(31 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(4 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(4 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_32X32
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_32X32_gen;
  SRAM_128X22_gen: if (address_width = 7) and (data_width = 22) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(21 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(21 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(6 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(6 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_128X22
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_128X22_gen;
  SRAM_1024X8_gen: if (address_width = 10) and (data_width = 8) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(7 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(7 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(9 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(9 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_1024X8
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_1024X8_gen;
  SRAM_1024X64_gen: if (address_width = 10) and (data_width = 64) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(63 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(63 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(9 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(9 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_1024X64
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_1024X64_gen;
  SRAM_64X128_gen: if (address_width = 6) and (data_width = 128) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(127 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(127 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(5 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(5 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_64X128
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_64X128_gen;
  SRAM_64X67_gen: if (address_width = 6) and (data_width = 67) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(66 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(66 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(5 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(5 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_64X67
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_64X67_gen;
  SRAM_64X24_gen: if (address_width = 6) and (data_width = 24) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(23 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(23 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(5 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(5 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_64X24
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_64X24_gen;
  SRAM_64X90_gen: if (address_width = 6) and (data_width = 90) generate
     mc: block 
            signal DATA_TIE_LOW  : std_logic_vector(89 downto 0); 
            signal DATA_TIE_HIGH : std_logic_vector(89 downto 0); 
            signal ADDR_TIE_LOW  : std_logic_vector(5 downto 0); 
            signal ADDR_TIE_HIGH : std_logic_vector(5 downto 0); 
         begin 
              DATA_TIE_LOW <= (others => '0'); 
              DATA_TIE_HIGH <= (others => '1'); 
              ADDR_TIE_LOW <= (others => '0'); 
              ADDR_TIE_HIGH <= (others => '1'); 
               inst: SRAM_64X90
   port map ( A => ADDR,  CLK => CLK, WEB => WRITE_BAR, BWEB => DATA_TIE_LOW, CEB => ENABLE_BAR,  D => DATAIN, Q => DATAOUT,  SLP => TIE_LOW, SD => TIE_LOW, CEBM => TIE_HIGH, WEBM => TIE_HIGH, BWEBM => DATA_TIE_HIGH, AM => ADDR_TIE_HIGH, DM => DATA_TIE_HIGH, BIST  => TIE_LOW);
         end block;
  end generate SRAM_64X90_gen;
end StructGen;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--
-- dual port synchronous memory.
--   similar to a flip-flop as far as simultaneous read/write  is concerned
--   if both ports try to write to the same address, the second port (1) wins
--
entity base_bank_dual_port_for_vivado is
   generic ( name: string;  g_addr_width: natural := 10; g_data_width : natural := 16);
	port(
		clka : in std_logic;
		clkb : in std_logic;
		ena : in std_logic;
		enb : in std_logic;
		wea : in std_logic;
		web : in std_logic;
		addra : in std_logic_vector(g_addr_width-1 downto 0);
		addrb : in std_logic_vector(g_addr_width-1 downto 0);
		dia : in std_logic_vector(g_data_width-1 downto 0);
		dib : in std_logic_vector(g_data_width-1 downto 0);
		doa : out std_logic_vector(g_data_width-1 downto 0);
		dob : out std_logic_vector(g_data_width-1 downto 0)
		);
end entity base_bank_dual_port_for_vivado;


architecture XilinxBramInfer of base_bank_dual_port_for_vivado is
  type MemArray is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);
  shared variable mem_array : MemArray((2**g_addr_width)-1 downto 0) := (others => (others => '0'));
begin  -- XilinxBramInfer


 process(CLKA)	
	begin
	if CLKA'event and CLKA = '1' then
			if ENA = '1' then
					DOA <= mem_array(to_integer(unsigned(ADDRA)));
				if WEA = '1' then
					mem_array(to_integer(unsigned(ADDRA))) := DIA;
				end if;
			end if;
		end if;
	end process;

	process(CLKB)
	begin
		if CLKB'event and CLKB = '1' then
			if ENB = '1' then
				DOB <= mem_array(to_integer(unsigned(ADDRB)));
				if WEB = '1' then
					mem_array(to_integer(unsigned(ADDRB))) := DIB;
				end if;
			end if;
		end if;
	end process;
end XilinxBramInfer;


------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.

------------------------------------------------------------------------------------------------
-- modified base-bank dual-port implementation by Kalyani
-------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;

entity base_bank_dual_port_r_wrap is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity base_bank_dual_port_r_wrap;
architecture RecWrap of base_bank_dual_port_r_wrap is
begin
	rinst: base_bank_dual_port 
		generic map (name => name, g_addr_width => g_addr_width, g_data_width => g_data_width)
		port map (
				datain_0 => datain_0,
				dataout_0 => dataout_0,
				addrin_0 => addrin_0,
				enable_0 => enable_0,
				writebar_0 => writebar_0,
				datain_1 => datain_1,
				dataout_1 => dataout_1,
				addrin_1 => addrin_1,
				enable_1 => enable_1,
				writebar_1 => writebar_1,
				clk => clk , reset => reset
			);
end RecWrap;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

library ahir;
use ahir.Types.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.MemcutDescriptionPackage.all;
use ahir.mem_component_pack.all;

entity base_bank_dual_port is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity base_bank_dual_port;


architecture improved_struct of base_bank_dual_port is
  component base_bank_dual_port_r_wrap is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
   end component base_bank_dual_port_r_wrap;

	constant best_cut_info: IntegerArray(1 to 5) :=
			find_best_cut (dpmem_cut_address_widths, 
					dpmem_cut_data_widths,
					dpmem_cut_row_heights,
					g_addr_width, g_data_width);
	constant best_cut_address_width : integer := best_cut_info(2);
	constant best_cut_data_width    : integer := best_cut_info(3);
	constant best_cut_nrows         : integer := best_cut_info(4);
	constant best_cut_ncols         : integer := best_cut_info(5);
	constant use_side_strip: boolean :=
			(best_cut_info(1) > 0) and
					((best_cut_data_width*best_cut_ncols) < g_data_width);
begin
	noCutFound: if (best_cut_info(1) <= 0) generate
		regbb_inst: base_bank_dual_port_with_registers
				generic map (name => name & ":regs", g_addr_width => g_addr_width,
						g_data_width => g_data_width)
			        port map (
					datain_0 => datain_0, 
					dataout_0 => dataout_0, 
					addrin_0 => addrin_0,
					enable_0 => enable_0, 
					writebar_0 => writebar_0, 
					datain_1 => datain_1, 
					dataout_1 => dataout_1, 
					addrin_1 => addrin_1,
					enable_1 => enable_1, 
					writebar_1 => writebar_1, 
					clk => clk,
					reset => reset);
	end generate noCutFound;

	cutFound: if (best_cut_info(1) > 0) generate

           mb: block
		-- declare array access signals.
		constant array_addr_width : integer := g_addr_width;
		constant array_data_width : integer := best_cut_data_width*best_cut_ncols;

		signal array_datain_0: std_logic_vector(array_data_width-1 downto 0);
		signal array_dataout_0: std_logic_vector(array_data_width-1 downto 0);

		signal array_datain_1: std_logic_vector(array_data_width-1 downto 0);
		signal array_dataout_1: std_logic_vector(array_data_width-1 downto 0);

		signal latch_dataout_0, latch_dataout_1: std_logic;
		
		signal dataout_0_sig, dataout_1_sig, dataout_0_reg, dataout_1_reg:
			std_logic_vector(g_data_width-1 downto 0);
           begin

		array_datain_0 <= datain_0 (g_data_width-1 downto (g_data_width - array_data_width));
		dataout_0_sig (g_data_width-1 downto (g_data_width - array_data_width)) <= array_dataout_0;

		array_datain_1 <= datain_1 (g_data_width-1 downto (g_data_width - array_data_width));
		dataout_1_sig (g_data_width-1 downto (g_data_width - array_data_width)) <= array_dataout_1;


		-- selector array..
		arrayInst: dpmem_selector_array 
				generic map (name =>  name & ":marray",
						g_addr_width => array_addr_width,
						g_data_width => array_data_width,
						g_base_addr_width => best_cut_address_width,
						g_base_data_width => best_cut_data_width)
				port map (
					datain_0   =>  array_datain_0,
					dataout_0  =>  array_dataout_0,
					addrin_0   =>  addrin_0,
					enable_0   =>  enable_0,
				        writebar_0 =>  writebar_0,
					datain_1   =>  array_datain_1,
					dataout_1  =>  array_dataout_1,
					addrin_1   =>  addrin_1,
					enable_1   =>  enable_1,
				        writebar_1 =>  writebar_1,
					clk => clk,
					reset => reset);


		genSideStrip : if use_side_strip generate
		  sb: block
			signal sstrip_datain_0: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
			signal sstrip_datain_1: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
			signal sstrip_dataout_0: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
			signal sstrip_dataout_1: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
		  begin

			sstrip_datain_0 <= datain_0((g_data_width-array_data_width)-1 downto 0);
			dataout_0_sig((g_data_width-array_data_width)-1 downto 0) <= sstrip_dataout_0;

			sstrip_datain_1 <= datain_1((g_data_width-array_data_width)-1 downto 0);
			dataout_1_sig((g_data_width-array_data_width)-1 downto 0) <= sstrip_dataout_1;

			side_strip_inst: component base_bank_dual_port_r_wrap
				generic map (name => name & ":sstrip", 
						g_addr_width => g_addr_width,
						g_data_width => (g_data_width - array_data_width))
			        port map (
					datain_0 => sstrip_datain_0, 
					dataout_0 => sstrip_dataout_0, 
					addrin_0 => addrin_0,
					enable_0 => enable_0, 
					writebar_0 => writebar_0, 
					datain_1 => sstrip_datain_1, 
					dataout_1 => sstrip_dataout_1, 
					addrin_1 => addrin_1,
					enable_1 => enable_1, 
					writebar_1 => writebar_1, 
					clk => clk,
					reset => reset);
		   end block sb;
		end generate genSideStrip;

  	    	process(clk, reset)
  	    	begin
			if(clk'event and clk = '1') then
				if(reset = '1') then
					latch_dataout_0 <= '0';
					latch_dataout_1 <= '0';
				else
					latch_dataout_0 <= enable_0 and writebar_0;
					latch_dataout_1 <= enable_1 and writebar_1;
				end if;
			end if;
  	    	end process;
	
      	    	process (clk, latch_dataout_0, dataout_0_sig, latch_dataout_1, dataout_1_sig)
  	    	begin
			if(clk'event and clk = '1') then
				if(latch_dataout_0 = '1') then
					dataout_0_reg <= dataout_0_sig;
				end if;
				if(latch_dataout_1 = '1') then
					dataout_1_reg <= dataout_1_sig;
				end if;
			end if;
  	    	end process;
	
            	dataout_0 <= dataout_0_reg when (latch_dataout_0 = '0') else dataout_0_sig;
            	dataout_1 <= dataout_1_reg when (latch_dataout_1 = '0') else dataout_1_sig;
            
          end block mb;
	end generate cutFound;

end improved_struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.

------------------------------------------------------------------------------------------------
-- modified base-bank implementation by Kalyani
-------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;
entity base_bank_r_wrap  is
   generic ( name: string:="mem"; g_addr_width: natural := 5; 
	     g_data_width : natural := 20);
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity;

architecture WrapRec of base_bank_r_wrap is
begin
 ci: base_bank
	generic map (name => name, g_addr_width => g_addr_width, g_data_width => g_data_width)
	port map (
			datain => datain, dataout => dataout, addrin => addrin,
			enable => enable, writebar => writebar, clk => clk, reset => reset
		 );
end WrapRec;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

library ahir;
use ahir.Types.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.MemcutDescriptionPackage.all;
use ahir.mem_component_pack.all;

entity base_bank is
   generic ( name: string:="mem"; g_addr_width: natural := 5; 
	     g_data_width : natural := 20);
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity base_bank;


architecture improved_struct of base_bank is

   component base_bank_r_wrap  is
   generic ( name: string:="mem"; g_addr_width: natural := 5; 
	     g_data_width : natural := 20);
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
   end component;

	constant best_cut_info: IntegerArray(1 to 5) :=
			find_best_cut (spmem_cut_address_widths, 
					spmem_cut_data_widths,
					spmem_cut_row_heights,
					g_addr_width, g_data_width);
	constant best_cut_address_width : integer := best_cut_info(2);
	constant best_cut_data_width    : integer := best_cut_info(3);
	constant best_cut_nrows         : integer := best_cut_info(4);
	constant best_cut_ncols         : integer := best_cut_info(5);
	constant use_side_strip: boolean :=
			(best_cut_info(1) > 0) and
					((best_cut_data_width*best_cut_ncols) < g_data_width);
begin
	noCutFound: if (best_cut_info(1) <= 0) generate
		regbb_inst: base_bank_with_registers
				generic map (name => name & ":regs", g_addr_width => g_addr_width,
						g_data_width => g_data_width)
			        port map (
					datain => datain, dataout => dataout, addrin => addrin,
						enable => enable, writebar => writebar, clk => clk,
							reset => reset);
	end generate noCutFound;

	cutFound: if (best_cut_info(1) > 0) generate

           mb: block
		-- declare array access signals.
		constant array_addr_width : integer := g_addr_width;
		constant array_data_width : integer := best_cut_data_width*best_cut_ncols;

		signal array_datain: std_logic_vector(array_data_width-1 downto 0);
		signal array_dataout: std_logic_vector(array_data_width-1 downto 0);

		signal latch_dataout: std_logic;
		signal dataout_sig, dataout_reg: std_logic_vector(g_data_width-1 downto 0);	
           begin

		array_datain <= datain (g_data_width-1 downto (g_data_width - array_data_width));
		dataout_sig (g_data_width-1 downto (g_data_width - array_data_width)) <= array_dataout;

		-- selector array..
		arrayInst: spmem_selector_array 
				generic map (name =>  name & ":marray",
						g_addr_width => array_addr_width,
						g_data_width => array_data_width,
						g_base_addr_width => best_cut_address_width,
						g_base_data_width => best_cut_data_width)
				port map (
					datain   =>  array_datain,
					dataout  =>  array_dataout,
					addrin   =>  addrin,
					enable   =>  enable,
				        writebar =>  writebar,
					clk => clk,
					reset => reset);


		genSideStrip : if use_side_strip generate
		  sb: block
			signal sstrip_datain: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
			signal sstrip_dataout: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
		  begin

			sstrip_datain <= datain((g_data_width-array_data_width)-1 downto 0);
			dataout_sig ((g_data_width-array_data_width)-1 downto 0) <= sstrip_dataout;

			side_strip_inst: component base_bank_r_wrap
				generic map (name => name & ":sstrip", 
						g_addr_width => g_addr_width,
						g_data_width => (g_data_width - array_data_width))
			        port map (
					datain => sstrip_datain, 
					dataout => sstrip_dataout, 
					addrin => addrin,
					enable => enable, 
					writebar => writebar, 
					clk => clk,
					reset => reset);

		   end block sb;
		end generate genSideStrip;

  	    	process(clk, reset)
  	    	begin
			if(clk'event and clk = '1') then
				if(reset = '1') then
					latch_dataout <= '0';
				else
					latch_dataout <= enable and writebar;
				end if;
			end if;
  	    	end process;
	
      	    	process (clk, latch_dataout, dataout_sig)
  	    	begin
			if(clk'event and clk = '1') then
				if(latch_dataout = '1') then
					dataout_reg <= dataout_sig(dataout'length-1 downto 0);
				end if;
			end if;
  	    	end process;
	
            	dataout <= dataout_reg when (latch_dataout = '0') else dataout_sig;
            
          end block mb;
	end generate cutFound;

end improved_struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;

use ahir.MemcutDescriptionPackage.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.mem_component_pack.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

entity dpmem_column is
   generic (name: string:="dpmem_column"; 
	g_addr_width: natural := 2;
	g_base_bank_addr_width: natural:=4; 
	g_base_bank_data_width : natural := 4);
   port (datain_0 : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity dpmem_column;


architecture struct of dpmem_column is

  --finding the number of row-replications in the column being build
  constant n_rows: integer := 2**(Maximum(0, g_addr_width - g_base_bank_addr_width));
  type WordArray is array  ( natural range <> ) of std_logic_vector (g_base_bank_data_width-1 downto 0);

  --fixing the size of address to maximum of addr_width, cut_width
  constant resized_addr_width: integer := Maximum (g_addr_width, g_base_bank_addr_width);
  
  signal resized_addrin_0: std_logic_vector(resized_addr_width-1 downto 0);  
  signal resized_addrin_1: std_logic_vector(resized_addr_width-1 downto 0);  

begin

  process (addrin_0, addrin_1)
	begin 
		resized_addrin_0 <= (others => '0');
		resized_addrin_1 <= (others => '0');
		resized_addrin_0(addrin_0'length-1 downto 0) <= addrin_0;
		resized_addrin_1(addrin_1'length-1 downto 0) <= addrin_1;
  end process;
	
  rowgen_block : block
	  signal decoded_CSB_0, decoded_CSB_0_d: std_logic_vector(n_rows-1 downto 0):= (others=>'1');
	  signal decoded_CSB_1, decoded_CSB_1_d: std_logic_vector(n_rows-1 downto 0):= (others=>'1');
	  
  	   signal dataout_array_0 : WordArray(n_rows-1 downto 0);
  	   signal dataout_array_1 : WordArray(n_rows-1 downto 0);

	begin
	  process(enable_0, resized_addrin_0, clk, reset)
	  	variable decoded_CSB_0_var: 
			std_logic_vector(2**Maximum(0, g_addr_width-g_base_bank_addr_width)-1 downto 0):= 
								(others=>'1');
	    begin
		if (enable_0 = '1' and reset = '0') then
		  decoded_CSB_0_var := MemDecoder(resized_addrin_0(resized_addr_width-1
		  downto resized_addr_width - Ceil_log2(n_rows)));
		else 
		  decoded_CSB_0_var := (others=>'1');
		end if;
		
		decoded_CSB_0 <= decoded_CSB_0_var;
		if(clk'event and clk = '1') then
			decoded_CSB_0_d <= decoded_CSB_0_var;
	 	end if;

	  end process;
	  
	  process(enable_1, resized_addrin_1,  clk, reset)
	  	variable decoded_CSB_1_var: 
			std_logic_vector(2**Maximum(0, g_addr_width-g_base_bank_addr_width)-1 downto 0)
										:= (others=>'1');
	    begin
		if (enable_1 = '1' and reset = '0') then
		  decoded_CSB_1_var := MemDecoder(resized_addrin_1(resized_addr_width-1
		  downto resized_addr_width - Ceil_log2(n_rows)));
		else 
		  decoded_CSB_1_var := (others=>'1');
		end if;
		decoded_CSB_1 <= decoded_CSB_1_var;
		if(clk'event and clk = '1') then
			decoded_CSB_1_d <= decoded_CSB_1_var;
	 	end if;
	  end process;

	  row_gen: for j in 0 to n_rows-1 generate
		mem_inst: dpmem_selector generic map(address_width => g_base_bank_addr_width,
					data_width => g_base_bank_data_width )
		port map(ADDR_0 => resized_addrin_0 (g_base_bank_addr_width-1 downto 0),
			 ADDR_1 => resized_addrin_1 (g_base_bank_addr_width-1 downto 0),
			 ENABLE_0_BAR => decoded_CSB_0(j),
			 ENABLE_1_BAR => decoded_CSB_1(j),
			 WRITE_0_BAR  => writebar_0,
			 WRITE_1_BAR  => writebar_1,
			 DATAIN_0 => datain_0,
			 DATAIN_1 => datain_1,
			 DATAOUT_0 => dataout_array_0(j),
			 DATAOUT_1 => dataout_array_1(j),
			 CLK => clk, RESET => reset );
	  end generate row_gen;

	-- muxes.
          process(dataout_array_0, decoded_CSB_0_d)
		variable sel_data_var: std_logic_vector(g_base_bank_data_width-1 downto 0);
	  begin
		sel_data_var := (others => '0');
		for I in 0 to n_rows-1 loop
			if(decoded_CSB_0_d(I) = '0') then
				sel_data_var := dataout_array_0(I);
			end if;
		end loop;
		dataout_0 <= sel_data_var;
	  end process;
          process(dataout_array_1, decoded_CSB_1_d)
		variable sel_data_var: std_logic_vector(g_base_bank_data_width-1 downto 0);
	  begin
		sel_data_var := (others => '0');
		for I in 0 to n_rows-1 loop
			if(decoded_CSB_1_d(I) = '0') then
				sel_data_var := dataout_array_1(I);
			end if;
		end loop;
		dataout_1 <= sel_data_var;
	  end process;
  end block rowgen_block;
end struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
-------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.MemcutDescriptionPackage.all;
use ahir.mem_component_pack.all;

entity dpmem_selector_array is
   generic ( name: string:="mem";
		 g_addr_width: natural := 5; 
	      	 g_data_width : natural := 20;
		 g_base_addr_width: natural := 5; 
	      	 g_base_data_width : natural := 20
	   );
   port (datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_0: out std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
	 datain_1 : in std_logic_vector(g_data_width-1 downto 0);
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity;

architecture Struct of dpmem_selector_array is
	constant NCOLS : integer := (g_data_width/g_base_data_width);
begin
	assert((NCOLS*g_base_data_width) = g_data_width) report
		"In " & name & " g_data_width is not an exact multiple of g_base_data_width" 
			severity FAILURE;

	CGEN: for COL in 0 to NCOLS-1 generate
	     sel_inst: dpmem_column
		generic map (g_addr_width => g_addr_width,
				g_base_bank_addr_width => g_base_addr_width,
				g_base_bank_data_width => g_base_data_width)
			port map (
				datain_0  => datain_0(((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
				dataout_0 => dataout_0(((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
         			addrin_0 => addrin_0,
         			enable_0 => enable_0,
         			writebar_0 => writebar_0,
				datain_1  => datain_1(((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
				dataout_1 => dataout_1(((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
         			addrin_1 => addrin_1,
         			enable_1 => enable_1,
         			writebar_1 => writebar_1,
         			clk => clk,
         			reset => reset);
	end generate CGEN;
end Struct;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity spram_generic_reverse_wrapper is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR : in std_logic_vector(address_width-1 downto 0 );
		CLK : in std_logic;
		WRITE_BAR: in std_logic;
		ENABLE_BAR: in std_logic;
		DATAIN  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT  : out std_logic_vector(data_width-1 downto 0));
end entity spram_generic_reverse_wrapper;

architecture XilinxBramInfer of spram_generic_reverse_wrapper is
  type MemArray is array (natural range <>) of std_logic_vector(data_width-1 downto 0);
  signal mem_array : MemArray((2**address_width)-1 downto 0) := (others => (others => '0'));
begin  -- XilinxBramInfer

  -- read/write process
  process(CLK, ADDR, ENABLE_BAR, WRITE_BAR)
  begin

    -- synch read-write memory
    if(CLK'event and CLK ='1') then
      if(ENABLE_BAR = '0' and WRITE_BAR = '0') then
        mem_array(To_Integer(unsigned(ADDR))) <= DATAIN;
      end if;
    end if;
  end process;

  -- read data.
  process(clk) 
  begin
	if(clk'event and clk = '1') then
		if(ENABLE_BAR = '0') then
		 	DATAOUT  <= mem_array(To_Integer(unsigned(ADDR)));
		end if;
	end if;
  end process;

end XilinxBramInfer;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_ASIC_components.all;
use ahir.GlobalConstants.all;
use ahir.mem_component_pack.all;

-- Entity to instantiate different available memory cuts based on the 
-- address_width and data_width generics passed.
entity dpram_generic_reverse_wrapper is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		WRITE_0_BAR : in std_logic;
		WRITE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAIN_1  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_0  : out std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK: in std_logic);
end entity dpram_generic_reverse_wrapper;


architecture XilinxBramInfer of dpram_generic_reverse_wrapper is

  type MemArray is array (natural range <>) of std_logic_vector(data_width-1 downto 0);

begin  -- XilinxBramInfer
  genVivado: if global_use_vivado_bbank_dual_port generate
    gVblock: block
	signal ena, enb, wea, web: std_logic;
    begin
	ena <= not ENABLE_0_bAR;
	enb <= not ENABLE_1_bAR;
	wea <= not WRITE_0_BAR;
	web <= not WRITE_1_BAR;

	bbVivado: base_bank_dual_port_for_vivado
		generic map (name => "bbVivado", g_addr_width => address_Width, g_data_width => data_width)
		port map (
			clka => clk, 
			clkb => clk, 
			ena => ena,
			enb => enb,
			wea => wea,
			web => web,
			addra => ADDR_0,
			addrb => ADDR_1,
			dia => DATAIN_0,
			dib => DATAIN_1,
			doa => DATAOUT_0,
			dob => DATAOUT_1
		);
      end block;
  end generate genVivado;

  noGenVivado: if not global_use_vivado_bbank_dual_port generate
  bbNoGen: block
  	signal mem_array : MemArray((2**address_width)-1 downto 0) := (others => (others => '0'));
  begin
  -- read/write process
  process(CLK, ADDR_0, ENABLE_0_BAR, WRITE_0_BAR, ADDR_1, ENABLE_1_BAR, WRITE_1_BAR)
  begin


    -- synch read-write memory
    if(CLK'event and CLK ='1') then

      -- both ports write.. second one wins if writes
      -- are to the same address.
      if(ENABLE_0_BAR = '0' and WRITE_0_BAR = '0') then
        mem_array(To_Integer(unsigned(ADDR_0))) <= DATAIN_0;
      end if;
      if(ENABLE_1_BAR = '0' and WRITE_1_BAR = '0') then
        mem_array(To_Integer(unsigned(ADDR_1))) <= DATAIN_1;
      end if;
    end if;
  end process;
      	
  process(clk) 
  begin
	if(clk'event and clk = '1') then
		if(ENABLE_0_BAR = '0') then
  			DATAOUT_0 <= mem_array(To_Integer(unsigned(ADDR_0)));
		end if;
		if(ENABLE_1_BAR = '0') then
  			DATAOUT_1 <= mem_array(To_Integer(unsigned(ADDR_1)));
		end if;
	end if;
  end process;
  end block;
  end generate noGenVivado;
  
end XilinxBramInfer;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity register_file_1w_1r_generic_reverse_wrapper is
	generic(address_width: integer:=8; data_width: integer:=8);
	port (ADDR_0 : in std_logic_vector(address_width-1 downto 0 );
		ADDR_1 : in std_logic_vector(address_width-1 downto 0 );
		ENABLE_0_BAR : in std_logic;
		ENABLE_1_BAR : in std_logic;
		DATAIN_0  : in std_logic_vector(data_width-1 downto 0);
		DATAOUT_1  : out std_logic_vector(data_width-1 downto 0);
		CLK: in std_logic);
end entity;

architecture XilinxBramInfer of register_file_1w_1r_generic_reverse_wrapper is

  type MemArray is array (natural range <>) of std_logic_vector(data_width-1 downto 0);
  signal mem_array : MemArray((2**address_width)-1 downto 0) := (others => (others => '0'));

begin  -- XilinxBramInfer

  -- read/write process
  process(CLK, ADDR_0, ENABLE_0_BAR, ADDR_1, ENABLE_1_BAR)
  begin

    -- synch read-write memory
    if(CLK'event and CLK ='1') then

      -- port 0 writes.
      if(ENABLE_0_BAR = '0') then
        mem_array(To_Integer(unsigned(ADDR_0))) <= DATAIN_0;
      end if;
    end if;
  end process;
      	
  process(clk) 
  begin
	if(clk'event and clk = '1') then
		if(ENABLE_1_BAR = '0') then
  			DATAOUT_1 <= mem_array(To_Integer(unsigned(ADDR_1)));
		end if;
	end if;
  end process;

end XilinxBramInfer;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;

use ahir.MemcutDescriptionPackage.all;
use ahir.MemCutsPackage.all;
use ahir.mem_component_pack.all;
use ahir.mem_ASIC_components.all;
use ahir.MemcutDescriptionPackage.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

entity register_file_1w_1r_column is
   generic ( name: string:="register_file_1w_1r_column"; 
	g_addr_width: natural := 2;
	g_base_bank_addr_width: natural:=4; 
	g_base_bank_data_width : natural := 4);
   port (datain_0 : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         dataout_1: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity register_file_1w_1r_column;


architecture struct of register_file_1w_1r_column is

  --finding the number of row-replications in the column being build
  constant n_rows: integer := 2**(Maximum(0, g_addr_width - g_base_bank_addr_width));
  type WordArray is array  ( natural range <> ) of std_logic_vector (g_base_bank_data_width-1 downto 0);

  --fixing the size of address to maximum of addr_width, cut_width
  constant resized_addr_width: integer := Maximum (g_addr_width, g_base_bank_addr_width);
  
  signal resized_addrin_0: std_logic_vector(resized_addr_width-1 downto 0);  
  signal resized_addrin_1: std_logic_vector(resized_addr_width-1 downto 0);  

begin

  
  process (addrin_0, addrin_1)
	begin 
		resized_addrin_0 <= (others => '0');
		resized_addrin_1 <= (others => '0');
		resized_addrin_0(addrin_0'length-1 downto 0) <= addrin_0;
		resized_addrin_1(addrin_1'length-1 downto 0) <= addrin_1;
  end process;
	
  rowgen_block: block

	  signal decoded_CSB_0, decoded_CSB_0_d: std_logic_vector(n_rows-1 downto 0):= (others=>'1');
	  signal decoded_CSB_1, decoded_CSB_1_d: std_logic_vector(n_rows-1 downto 0):= (others=>'1');
	  
  	  signal dataout_array_0 : WordArray(n_rows-1 downto 0);
  	  signal dataout_array_1 : WordArray(n_rows-1 downto 0);

  begin
	  process(enable_0, resized_addrin_0, clk, reset)
	  	variable decoded_CSB_0_var: 
			std_logic_vector(2**Maximum(0, g_addr_width-g_base_bank_addr_width)-1 
										downto 0):= (others=>'1');
	  begin
		if (enable_0 = '1') then
		  decoded_CSB_0_var := MemDecoder(resized_addrin_0(resized_addr_width-1
		  					downto resized_addr_width - Ceil_log2(n_rows)));
		else 
		  decoded_CSB_0_var := (others=>'1');
		end if;
		
		decoded_CSB_0 <= decoded_CSB_0_var;

		if(clk'event and clk = '1') then
			decoded_CSB_0_d <= decoded_CSB_0_var;
		end if;
	  end process;
	  
	  process(enable_1, resized_addrin_1)
	  	variable decoded_CSB_1_var: 
			std_logic_vector(2**Maximum(0, g_addr_width-g_base_bank_addr_width)-1 downto 0)
							:= (others=>'1');
	    begin
		if (enable_1 = '1') then
		  decoded_CSB_1_var := MemDecoder(resized_addrin_1(resized_addr_width-1
		  downto resized_addr_width - Ceil_log2(n_rows)));
		else 
		  decoded_CSB_1_var := (others=>'1');
		end if;
		decoded_CSB_1 <= decoded_CSB_1_var;

		if(clk'event and clk = '1') then
			decoded_CSB_1_d <= decoded_CSB_1_var;
		end if;
	  end process;

	  row_gen: for j in 0 to n_rows-1 generate
		mem_inst: register_file_1w_1r_selector generic map(address_width => g_base_bank_addr_width,
					data_width => g_base_bank_data_width )
			port map(ADDR_0 => resized_addrin_0 (g_base_bank_addr_width-1 downto 0),
				 ENABLE_0_BAR => decoded_CSB_0(j),
				 ADDR_1 => resized_addrin_1 (g_base_bank_addr_width-1 downto 0),
				 ENABLE_1_BAR => decoded_CSB_1(j),
				 DATAIN_0  => datain_0,
				 DATAOUT_1 => dataout_array_1(j),
				 CLK     => clk, 
				 RESET   => reset);
	  end generate row_gen;

	-- mux.
          process(dataout_array_1, decoded_CSB_1_d)
		variable sel_data_var: std_logic_vector(g_base_bank_data_width-1 downto 0);
	  begin
		sel_data_var := (others => '0');
		for I in 0 to n_rows-1 loop
			if(decoded_CSB_1_d(I) = '0') then
				sel_data_var := dataout_array_1(I);
			end if;
		end loop;
		dataout_1 <= sel_data_var;
	  end process;
   end block;


end struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.mem_component_pack.all;

entity register_file_1w_1r_port_r_wrap is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 -- write port 0
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
	 -- read port 1
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
	
         clk: in std_logic;
         reset : in std_logic);
end entity register_file_1w_1r_port_r_wrap;

architecture RecWrap of register_file_1w_1r_port_r_wrap is
begin
	rinst: register_file_1w_1r_port
		generic map (name => name, g_addr_width => g_addr_width, g_data_width => g_data_width)
		port map (
				datain_0 => datain_0,
				addrin_0 => addrin_0,
				enable_0 => enable_0,
				dataout_1 => dataout_1,
				addrin_1 => addrin_1,
				enable_1 => enable_1,
				clk => clk, reset => reset
			);

end RecWrap;





library ahir;
use ahir.Utilities.all;
use ahir.GlobalConstants.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.GlobalConstants.all;
use ahir.mem_component_pack.all;
use ahir.MemCutsPackage.all;
use ahir.MemcutDescriptionPackage.all;
use ahir.mem_ASIC_components.all;
--
-- synchronous memory with 1 write and 1 read port.
--
entity register_file_1w_1r_port is
   generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   port (
	 -- write port 0
	 datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
	 -- read port 1
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
	
         clk: in std_logic;
         reset : in std_logic);
end entity register_file_1w_1r_port;


architecture improved_struct of register_file_1w_1r_port is
   component register_file_1w_1r_port_r_wrap is
   	generic ( name: string; g_addr_width: natural := 10; g_data_width : natural := 16);
   	port (
	 	-- write port 0
	 	datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         	addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         	enable_0: in std_logic;
	 	-- read port 1
         	dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         	addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         	enable_1: in std_logic;
		
         	clk: in std_logic;
         	reset : in std_logic);
   end component register_file_1w_1r_port_r_wrap;
	constant best_cut_info: IntegerArray(1 to 5) :=
			find_best_cut (register_file_1w_1r_cut_address_widths, 
					register_file_1w_1r_cut_data_widths,
					register_file_1w_1r_cut_row_heights,
					g_addr_width, g_data_width);
	constant best_cut_address_width : integer := best_cut_info(2);
	constant best_cut_data_width    : integer := best_cut_info(3);
	constant best_cut_nrows         : integer := best_cut_info(4);
	constant best_cut_ncols         : integer := best_cut_info(5);
	constant use_side_strip: boolean :=
			(best_cut_info(1) > 0) and
					((best_cut_data_width*best_cut_ncols) < g_data_width);
begin
	noCutFound: if (best_cut_info(1) <= 0) generate
		regbb_inst: register_file_1w_1r_port_with_registers
				generic map (name => name & ":regs", g_addr_width => g_addr_width,
						g_data_width => g_data_width)
			        port map (
					datain_0 => datain_0, 
					addrin_0 => addrin_0,
					enable_0 => enable_0, 
					dataout_1 => dataout_1, 
					addrin_1 => addrin_1,
					enable_1 => enable_1, 
					clk => clk,
					reset => reset);
	end generate noCutFound;

	cutFound: if (best_cut_info(1) > 0) generate

           mb: block
		-- declare array access signals.
		constant array_addr_width : integer := g_addr_width;
		constant array_data_width : integer := best_cut_data_width*best_cut_ncols;

		signal array_datain_0: std_logic_vector(array_data_width-1 downto 0);
		signal array_dataout_1: std_logic_vector(array_data_width-1 downto 0);

		signal latch_dataout_1: std_logic;
		
		signal dataout_1_sig, dataout_1_reg: std_logic_vector(g_data_width-1 downto 0);
           begin

		array_datain_0 <= datain_0(g_data_width-1 downto (g_data_width - array_data_width));
		dataout_1_sig (g_data_width-1 downto (g_data_width - array_data_width)) <= array_dataout_1;


		-- selector array..
		arrayInst: register_file_1w_1r_selector_array 
				generic map (name =>  name & ":marray",
						g_addr_width => array_addr_width,
						g_data_width => array_data_width,
						g_base_addr_width => best_cut_address_width,
						g_base_data_width => best_cut_data_width)
				port map (
					datain_0   =>  array_datain_0,
					addrin_0   =>  addrin_0,
					enable_0   =>  enable_0,
					dataout_1  =>  array_dataout_1,
					addrin_1   =>  addrin_1,
					enable_1   =>  enable_1,
					clk => clk,
					reset => reset);


		genSideStrip : if use_side_strip generate
		  sb: block
			signal sstrip_datain_0: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
			signal sstrip_dataout_1: std_logic_vector((g_data_width - array_data_width)-1 downto 0);
		  begin

			sstrip_datain_0 <= datain_0((g_data_width-array_data_width)-1 downto 0);
			dataout_1_sig((g_data_width-array_data_width)-1 downto 0) <= sstrip_dataout_1;

			side_strip_inst: component register_file_1w_1r_port_r_wrap
				generic map (name => name & ":sstrip", 
						g_addr_width => g_addr_width,
						g_data_width => (g_data_width - array_data_width))
			        port map (
					datain_0 => sstrip_datain_0, 
					addrin_0 => addrin_0,
					enable_0 => enable_0, 
					dataout_1 => sstrip_dataout_1, 
					addrin_1 => addrin_1,
					enable_1 => enable_1, 
					clk => clk,
					reset => reset);
		   end block sb;
		end generate genSideStrip;

  	    	process(clk, reset)
  	    	begin
			if(clk'event and clk = '1') then
				if(reset = '1') then
					latch_dataout_1 <= '0';
				else
					latch_dataout_1 <= enable_1;
				end if;
			end if;
  	    	end process;
	
      	    	process (clk, latch_dataout_1, dataout_1_sig)
  	    	begin
			if(clk'event and clk = '1') then
				if(latch_dataout_1 = '1') then
					dataout_1_reg <= dataout_1_sig;
				end if;
			end if;
  	    	end process;
	
            	dataout_1 <= dataout_1_reg when (latch_dataout_1 = '0') else dataout_1_sig;
            
          end block mb;
	end generate cutFound;

end improved_struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
-------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.MemcutDescriptionPackage.all;
use ahir.mem_component_pack.all;

entity register_file_1w_1r_selector_array is
   generic ( name: string:="mem";
		 g_addr_width: natural := 5; 
	      	 g_data_width : natural := 20;
		 g_base_addr_width: natural := 5; 
	      	 g_base_data_width : natural := 20
	   );
   port (datain_0 : in std_logic_vector(g_data_width-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         dataout_1: out std_logic_vector(g_data_width-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity;

architecture Struct of register_file_1w_1r_selector_array is
	constant NCOLS : integer := (g_data_width/g_base_data_width);
begin
	assert((NCOLS*g_base_data_width) = g_data_width) report
		"In " & name & " g_data_width is not an exact multiple of g_base_data_width" 
			severity FAILURE;

	CGEN: for COL in 0 to NCOLS-1 generate
	     sel_inst: register_file_1w_1r_column
		generic map (g_addr_width => g_addr_width,
				g_base_bank_addr_width => g_base_addr_width,
				g_base_bank_data_width => g_base_data_width)
			port map (
				datain_0  => datain_0(((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
         			addrin_0 => addrin_0,
         			enable_0 => enable_0,
				dataout_1 => dataout_1(((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
         			addrin_1 => addrin_1,
         			enable_1 => enable_1,
         			clk => clk,
         			reset => reset);
	end generate CGEN;
end Struct;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;	
use ahir.Types.all;	
use ahir.Subprograms.all;	
use ahir.mem_function_pack.all;
use ahir.memory_subsystem_package.all;

use ahir.MemcutDescriptionPackage.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.mem_component_pack.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

entity spmem_column is
   generic ( name: string:="spmem_column"; 
	g_addr_width: natural := 2;
	g_base_bank_addr_width: natural:=4; 
	g_base_bank_data_width : natural := 4);
   port (datain : in std_logic_vector(g_base_bank_data_width-1 downto 0);
         dataout: out std_logic_vector(g_base_bank_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity spmem_column;


architecture struct of spmem_column is

--finding the number of row-replications in the column being build
  constant n_rows: integer := 2**(Maximum(0, g_addr_width-g_base_bank_addr_width));

--fixing the size of address to maximum of addr_width, cut_width
  constant resized_addr_width: integer := Maximum(g_addr_width, g_base_bank_addr_width);
  signal resized_addrin: std_logic_vector(resized_addr_width-1 downto 0);  
  type WordArray is array  ( natural range <> ) of std_logic_vector (g_base_bank_data_width-1 downto 0);

begin
  process (addrin)
	begin 
		resized_addrin <= (others => '0');
		resized_addrin(addrin'length-1 downto 0) <= addrin;
  end process;
	
  rowgen_block: block
	  
  	   signal decoded_CSB, decoded_CSB_d: std_logic_vector(n_rows-1 downto 0):= (others=>'1');
  	   signal dataout_array : WordArray(n_rows-1 downto 0);

	  --chipselect is made low only when enable is high and reset is low.
	  --memory will not be read or written when enable is low.
	begin
	  process(resized_addrin, enable, clk)
	     variable decoded_CSB_var: std_logic_vector(2**Maximum(0, g_addr_width-g_base_bank_addr_width)-1 
							downto 0):= (others=>'1');
	    begin
		if (enable = '1') then
		  decoded_CSB_var := MemDecoder(resized_addrin(resized_addr_width-1
		  downto resized_addr_width-Ceil_log2(n_rows)));
		else 
		  decoded_CSB_var :=(others=>'1');
		end if;

		decoded_CSB <= decoded_CSB_var;
		if(clk'event and clk = '1') then
			decoded_CSB_d <= decoded_CSB_var;
		end if;
	  end process;
	  row_gen: for j in 0 to n_rows-1 generate
		mem_inst: spmem_selector generic map(address_width => g_base_bank_addr_width,
					data_width => g_base_bank_data_width )
			port map(ADDR => resized_addrin(g_base_bank_addr_width-1 downto 0),
				 CLK => clk,
				 RESET => reset,
				 WRITE_BAR => writebar,
				 ENABLE_BAR => decoded_CSB(j),
				 DATAIN => datain,
				 DATAOUT => dataout_array(j));
	  end generate row_gen;

  	  -- mux.
          process(dataout_array, decoded_CSB_d)
		variable sel_data_var: std_logic_vector(g_base_bank_data_width-1 downto 0);
	  begin
		sel_data_var := (others => '0');
		for I in 0 to n_rows-1 loop
			if(decoded_CSB_d(I) = '0') then
				sel_data_var := dataout_array(I);
			end if;
		end loop;
		dataout <= sel_data_var;
	  end process;
   end block;
  
end struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
-------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.MemCutsPackage.all;
use ahir.mem_ASIC_components.all;
use ahir.MemcutDescriptionPackage.all;
use ahir.mem_component_pack.all;

entity spmem_selector_array is
   generic ( name: string:="mem";
		 g_addr_width: natural := 5; 
	      	 g_data_width : natural := 20;
		 g_base_addr_width: natural := 5; 
	      	 g_base_data_width : natural := 20
	   );
   port (datain : in std_logic_vector(g_data_width-1 downto 0);
         dataout: out std_logic_vector(g_data_width-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity;

architecture Struct of spmem_selector_array is
	constant NCOLS : integer := (g_data_width/g_base_data_width);
begin
	assert((NCOLS*g_base_data_width) = g_data_width) report
		"In " & name & " g_data_width is not an exact multiple of g_base_data_width" 
			severity FAILURE;

	CGEN: for COL in 0 to NCOLS-1 generate
	     sel_inst: spmem_column
		generic map (g_addr_width => g_addr_width,
				g_base_bank_addr_width => g_base_addr_width,
				g_base_bank_data_width => g_base_data_width)
			port map (
				datain  => datain (((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
				dataout => dataout (((COL+1)*g_base_data_width)-1 downto (COL*g_base_data_width)),
				addrin => addrin,
				enable  => enable,
				writebar => writebar,
				clk => clk, reset => reset);
	end generate CGEN;
end Struct;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;

entity combinational_merge is
  generic (
    name: string;
    g_data_width       : natural;
    g_number_of_inputs: natural;
    g_time_stamp_width : natural);
  port(
    in_data: in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    in_tstamp: in std_logic_vector((g_number_of_inputs*g_time_stamp_width)-1 downto 0);
    out_data: out std_logic_vector(g_data_width-1 downto 0);
    out_tstamp: out std_logic_vector(g_time_stamp_width-1 downto 0);
    in_req: in std_logic_vector(g_number_of_inputs-1 downto 0);
    in_ack: out std_logic_vector(g_number_of_inputs-1 downto 0);
    out_req: out std_logic;
    out_ack: in std_logic);
end combinational_merge;

architecture combinational_merge of combinational_merge is

  signal sel_vector : std_logic_vector(g_number_of_inputs-1 downto 0);
  
begin  -- combinational_merge

  process(in_tstamp,in_data,in_req)
    variable best_tstamp_var : std_logic_vector(1 to g_time_stamp_width);
    variable best_data : std_logic_vector(1 to g_data_width);
    variable sel_var : std_logic_vector(g_number_of_inputs-1 downto 0);
    variable vflag : std_logic;
  begin
    Select_Best_Index(in_tstamp,in_data, in_req,best_tstamp_var,best_data,sel_var,vflag);
    if(vflag = '1') then
      out_tstamp <= best_tstamp_var;
      out_data <= best_data;
      sel_vector <= sel_var;
      out_req <= '1';
    else
      out_tstamp <= (others => '0');
      out_data <= (others => '0');
      sel_vector <= (others => '0');
      out_req <= '0';
    end if;
  end process;
  
  AckGen: for I in 0 to g_number_of_inputs-1 generate
    in_ack(I) <= '1' when (sel_vector(I) = '1'  and out_ack = '1' and in_req(I) = '1') else '0';
  end generate AckGen;
  
end combinational_merge;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity combinational_merge_with_repeater is
  generic (
    name: string;
    g_data_width       : natural;
    g_number_of_inputs: natural;
    g_time_stamp_width : natural);
  port(
    clk : in std_logic;
    reset : in std_logic;
    in_data: in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    in_tstamp: in std_logic_vector((g_number_of_inputs*g_time_stamp_width)-1 downto 0);
    out_data: out std_logic_vector(g_data_width-1 downto 0);
    out_tstamp: out std_logic_vector(g_time_stamp_width-1 downto 0);
    in_req: in std_logic_vector(g_number_of_inputs-1 downto 0);
    in_ack: out std_logic_vector(g_number_of_inputs-1 downto 0);
    out_req: out std_logic;
    out_ack: in std_logic);
end combinational_merge_with_repeater;

architecture Struct of combinational_merge_with_repeater is

  signal sel_vector : std_logic_vector(g_number_of_inputs-1 downto 0);

  signal rep_data_in : std_logic_vector(g_data_width-1 downto 0);
  signal rep_req_in, rep_ack_out: std_logic;
  
begin  

   cmerge: combinational_merge 
		generic map (name => name & "-cmerge", g_data_width => g_data_width,
			 g_number_of_inputs => g_number_of_inputs,
			 g_time_stamp_width => g_time_stamp_width)
		port map(in_data => in_data,
			 in_tstamp => in_tstamp,
			 out_data => rep_data_in,
			 out_tstamp => open,
			 in_req => in_req,
			 in_ack => in_ack,
			 out_req => rep_req_in,
			 out_ack => rep_ack_out);

    -- instantiate repeater only if the number of inputs is > 1.
    moreThanOneInputGen: if (g_number_of_inputs > 1) generate
    rptr:  mem_repeater generic map (name => name & "-rptr", g_data_width => g_data_width)
		port map(clk => clk, reset => reset,
			 data_in => rep_data_in,
			 req_in => rep_req_in,
			 ack_out => rep_ack_out,
			 data_out => out_data,
			 req_out => out_req,
			 ack_in => out_ack);	
    end generate moreThanOneInputGen;

    OneInputGen: if (g_number_of_inputs = 1) generate
         out_data <= rep_data_in;
         out_req  <= rep_req_in;
         rep_ack_out <= out_ack;
    end generate OneInputGen;
  
end Struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity demerge_tree is
  generic (
    name: string;
    g_demux_degree: natural := 10;
    g_number_of_outputs: natural := 5;
    g_data_width: natural := 8;
    g_id_width: natural := 3;
    g_stage_id: natural := 0
    );       

  port (
    demerge_data_out : out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
    demerge_ready_out  : out std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_accept_in   : in std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_data_in: in std_logic_vector(g_data_width-1 downto 0);
    demerge_ack_out : out std_logic;
    demerge_req_in  : in std_logic;
    demerge_sel_in: in std_logic_vector(g_id_width-1 downto 0);
    clock: in std_logic;
    reset: in std_logic);
end demerge_tree;

-- a much simpler architecture, which is likely to be equally
-- effective.
architecture Simple of demerge_tree is
  constant inserted_delay  : integer := Maximum(1,Ceil_Log2(g_number_of_outputs/g_demux_degree));
begin  -- Simple

  demux : mem_demux generic map (
    name => name & "-demux",
    g_data_width        => g_data_width,
    g_id_width          => g_id_width,
    g_number_of_outputs => g_number_of_outputs,
    g_delay_count => inserted_delay)
    port map (
      data_in  => demerge_data_in,
      sel_in   => demerge_sel_in,
      req_in   => demerge_req_in,
      ack_out  => demerge_ack_out,
      data_out => demerge_data_out,
      req_out  => demerge_ready_out,
      ack_in   => demerge_accept_in,
      clk      => clock,
      reset    => reset);
end Simple;




------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity demerge_tree_wrap is
  generic (
    name: string;
    g_demux_degree: natural;
    g_number_of_outputs: natural;
    g_data_width: natural;
    g_id_width: natural;
    g_stage_id: natural
    );       

  port (
    demerge_data_out : out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
    demerge_ready_out  : out std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_accept_in   : in std_logic_vector(g_number_of_outputs-1 downto 0);
    demerge_data_in: in std_logic_vector(g_data_width-1 downto 0);
    demerge_ack_out : out std_logic;
    demerge_req_in  : in std_logic;
    demerge_sel_in: in std_logic_vector(g_id_width-1 downto 0);
    clock: in std_logic;
    reset: in std_logic);
  
end demerge_tree_wrap;



architecture wrapper of demerge_tree_wrap is
begin
      
      demTree: component demerge_tree
        generic map (
          name => name & "-demTree", 
          g_data_width => g_data_width,
          g_id_width   => g_id_width,
          g_number_of_outputs => g_number_of_outputs,
          g_stage_id => g_stage_id,
          g_demux_degree => g_demux_degree)
        port map (
          demerge_data_out => demerge_data_out,
          demerge_ready_out => demerge_ready_out,
          demerge_accept_in => demerge_accept_in,
          demerge_data_in   => demerge_data_in,
          demerge_req_in  => demerge_req_in,
          demerge_ack_out => demerge_ack_out,
          demerge_sel_in  => demerge_sel_in,
          clock => clock,
          reset => reset);
end wrapper;




------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity mem_demux is
  generic ( name: string;
	    g_data_width: natural := 10;
            g_id_width : natural := 3;
            g_number_of_outputs: natural := 8;
	    g_delay_count: natural := 1);
  port(data_in: in std_logic_vector(g_data_width-1 downto 0);  -- data & id & time-stamp
       sel_in : in std_logic_vector(g_id_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0 );
       req_out: out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clk: in std_logic;
       reset: in std_logic);
end entity;

architecture behave of mem_demux is
  type SigArrayType is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);

  signal data_out_sig,repeater_out_sig : SigArrayType(g_number_of_outputs-1 downto 0);
  signal req_out_sig, ack_in_sig : std_logic_vector(g_number_of_outputs-1 downto 0);

begin  -- behave

 -- demux is required only if there is more than one output...
 MoreThanOneOutputGen:  if (g_number_of_outputs > 1) generate

  process(ack_in_sig)
    variable ack_out_var : std_logic;
  begin
    ack_out_var := '0';
    for I in 0 to g_number_of_outputs-1 loop
      ack_out_var := ack_out_var or ack_in_sig(I);
    end loop;  -- I
    ack_out <= ack_out_var;
  end process;
    
  gen: for I in 0 to g_number_of_outputs-1 generate

    data_out_sig(I) <= data_in;
    
    process(data_in, sel_in, req_in)
      variable port_index : natural;
    begin
      port_index := To_Integer(sel_in);
      req_out_sig(I) <= '0';
      if(req_in = '1' and port_index = I) then
        req_out_sig(I) <= req_in;
      end if;
    end process;
      
    Repeater : mem_shift_repeater generic map(name => name & "-Repeater", g_data_width => g_data_width, g_number_of_stages => g_delay_count)
    port map (
      clk      => clk,
      reset    => reset,
      data_in  => data_out_sig(I),
      req_in   => req_out_sig(I),
      ack_out  => ack_in_sig(I),
      data_out => repeater_out_sig(I),
      req_out  => req_out(I),
      ack_in   => ack_in(I));

    data_out((I+1)*g_data_width -1 downto I*g_data_width) <= repeater_out_sig(I);

  end generate gen;
 end generate MoreThanOneOutputGen;

 OnlyOneOutputGen: if (g_number_of_outputs = 1) generate

      data_out <= data_in;
      ack_out <= ack_in(0);
      req_out(0) <= req_in;

 end generate OnlyOneOutputGen;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

-- memory subsystem guarantees that accesses to the same location
-- will take place in the order of the time-stamp assigned to each
-- access (tie breaks will be random). Time-stamp is set at the
-- point of acceptance of an access request.

entity memory_subsystem_core is
  generic(name: string;
	  num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          time_stamp_width      : natural := 11;
          number_of_banks       : natural := 1;
          mux_degree            : natural := 10;
          demux_degree          : natural := 10;
	  base_bank_addr_width  : natural := 8;
	  base_bank_data_width  : natural := 8);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    -- time-stamp for request: will be used for all ordering inside
    -- the subsystem
    lr_time_stamp_in   : in  std_logic_vector((num_loads*time_stamp_width)-1 downto 0);
    
    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    -- time-stamp for request: will be used for all ordering inside
    -- the subsystem
    sr_time_stamp_in   : in  std_logic_vector((num_stores*time_stamp_width)-1 downto 0);
    
    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity memory_subsystem_core;


-- simplified logic.  Use one memory bank only..
architecture pipelined of memory_subsystem_core is

  	constant c_load_port_id_width : natural := Maximum(1,Ceil_Log2(num_loads));
  	constant c_store_port_id_width : natural := Maximum(1,Ceil_Log2(num_stores));

	signal lc_ack_out_sig : std_logic_vector(num_loads-1 downto 0);
	signal sc_ack_out_sig : std_logic_vector(num_stores-1 downto 0);

	signal load_request_selected: std_logic;
	signal load_request_accepted: std_logic;
	signal load_request_address: std_logic_vector(addr_width-1 downto 0);
	signal load_request_id, load_complete_id: unsigned(c_load_port_id_width-1 downto 0);
	signal load_request_tag: std_logic_vector((tag_width-1) downto 0);
	signal load_request_time_stamp: std_logic_vector((time_stamp_width-1) downto 0);

	signal load_request_selected_repeated: std_logic;
	signal load_request_accepted_repeated: std_logic;
	signal load_request_address_repeated: std_logic_vector(addr_width-1 downto 0);
	signal load_request_id_repeated : unsigned(c_load_port_id_width-1 downto 0);
	signal load_request_tag_repeated: std_logic_vector((tag_width-1) downto 0);
	signal load_request_time_stamp_repeated: std_logic_vector((time_stamp_width-1) downto 0);

	signal load_complete_data: std_logic_vector(data_width-1 downto 0);
	signal load_complete_ready: std_logic;
	signal load_complete_accept: std_logic;
	signal load_complete_tag: std_logic_vector((tag_width-1) downto 0);

	signal store_request_selected: std_logic;
	signal store_request_accepted: std_logic;
	signal store_request_address: std_logic_vector(addr_width-1 downto 0);
	signal store_request_data: std_logic_vector(data_width-1 downto 0);
	signal store_request_id, store_complete_id: unsigned(c_store_port_id_width-1 downto 0);
	signal store_request_tag: std_logic_vector((tag_width-1) downto 0);
	signal store_request_time_stamp: std_logic_vector((time_stamp_width-1) downto 0);

	signal store_request_selected_repeated: std_logic;
	signal store_request_accepted_repeated: std_logic;
	signal store_request_address_repeated: std_logic_vector(addr_width-1 downto 0);
	signal store_request_data_repeated: std_logic_vector(data_width-1 downto 0);
	signal store_request_id_repeated : unsigned(c_store_port_id_width-1 downto 0);
	signal store_request_tag_repeated: std_logic_vector((tag_width-1) downto 0);
	signal store_request_time_stamp_repeated: std_logic_vector((time_stamp_width-1) downto 0);

	signal store_complete_ready: std_logic;
	signal store_complete_accept: std_logic;
	signal store_complete_tag: std_logic_vector((tag_width-1) downto 0);


	signal store_complete_accept_array: std_logic_vector(num_stores-1 downto 0);
	signal load_complete_accept_array: std_logic_vector(num_loads-1 downto 0);

	signal lrr_data_in, lrr_data_out : 
		std_logic_vector((time_stamp_width + c_load_port_id_width + addr_width + tag_width)-1
					downto 0);
	signal srr_data_in, srr_data_out : 
		std_logic_vector(((time_stamp_width + c_store_port_id_width + addr_width + data_width + 
						tag_width)-1) downto 0);

begin

  -----------------------------------------------------------------------------
  -- stage 1: choose a load and store request with lowest time-stamp.  The request could be
  --          a read or a write.  
  -----------------------------------------------------------------------------
  process(lr_req_in, lr_time_stamp_in, lr_addr_in, lr_tag_in)
	variable load_request_selected_var: std_logic;
	variable load_request_address_var: std_logic_vector(addr_width-1 downto 0);
	variable load_request_id_var: unsigned(c_load_port_id_width-1 downto 0);
	variable load_request_tag_var: std_logic_vector((tag_width-1) downto 0);

	variable smallest_time_stamp_var: std_logic_vector(time_stamp_width-1 downto 0);
	variable curr_time_stamp_var: std_logic_vector(time_stamp_width-1 downto 0);
	variable none_valid_so_far: std_logic;



  begin
	none_valid_so_far := '1';

	load_request_selected_var := '0';
	load_request_address_var := (others => '0');
	load_request_id_var := (others => '0');
	load_request_tag_var := (others => '0');
	smallest_time_stamp_var := (others => '0');

	for I in  0 to num_loads-1 loop
		if(lr_req_in(I) = '1') then
			curr_time_stamp_var := 
				lr_time_stamp_in (((I+1)*time_stamp_width)-1 downto
								I*time_stamp_width);
			if ((none_valid_so_far = '1') or 
				IsGreaterThan(smallest_time_stamp_var,curr_time_stamp_var)) then
				none_valid_so_far := '0';
				smallest_time_stamp_var := curr_time_stamp_var;
				load_request_id_var := to_unsigned(I,c_load_port_id_width);
				load_request_selected_var := '1';
				load_request_address_var := 
					lr_addr_in(((I+1)*addr_width)-1 downto I*addr_width);
				load_request_tag_var := 
					lr_tag_in(((I+1)*tag_width)-1 downto I*tag_width);
			end if;
		end if;
	end loop;


	load_request_selected <= load_request_selected_var;
	load_request_id <= load_request_id_var;
	load_request_address <= load_request_address_var;
	load_request_tag <= load_request_tag_var;
	load_request_time_stamp <= smallest_time_stamp_var;

  end process;

  lrr_data_in <= load_request_time_stamp & to_slv(load_request_id) & 
					load_request_address & load_request_tag;

  load_request_time_stamp_repeated <= 
		lrr_data_out((time_stamp_width+c_load_port_id_width+addr_width+tag_width)-1 downto 
							(c_load_port_id_width+addr_width+tag_width));
  load_request_id_repeated <= to_unsigned(lrr_data_out((c_load_port_id_width+addr_width+tag_width)-1 
							downto (addr_width+tag_width)));
  load_request_address_repeated <= lrr_data_out((addr_width+tag_width)-1 downto tag_width);
  load_request_tag_repeated <= lrr_data_out(tag_width-1 downto 0);
  lrr : QueueBase
		generic map (name => name & ":lrr", 
				queue_depth => 2,
				data_width => (time_stamp_width + c_load_port_id_width + 
								addr_width + tag_width))
		port map (clk => clock, reset => reset,
				data_in => lrr_data_in,
				data_out => lrr_data_out,
				push_req =>  load_request_selected,
				push_ack =>  load_request_accepted,
				pop_req  =>  load_request_accepted_repeated,
				pop_ack  =>  load_request_selected_repeated);	

  process(sr_req_in, sr_time_stamp_in, sr_addr_in, sr_data_in, sr_tag_in)
	variable store_request_selected_var: std_logic;
	variable store_request_address_var: std_logic_vector(addr_width-1 downto 0);
	variable store_request_data_var: std_logic_vector(data_width-1 downto 0);
	variable store_request_id_var: unsigned(c_store_port_id_width-1 downto 0);
	variable store_request_tag_var: std_logic_vector((tag_width-1) downto 0);
	variable smallest_time_stamp_var: std_logic_vector(time_stamp_width-1 downto 0);
	variable curr_time_stamp_var: std_logic_vector(time_stamp_width-1 downto 0);
	variable none_valid_so_far: std_logic;

  begin
	none_valid_so_far := '1';

	store_request_selected_var := '0';
	store_request_address_var := (others => '0');
	store_request_data_var := (others => '0');
	store_request_id_var := (others => '0');
	store_request_tag_var := (others => '0');
	smallest_time_stamp_var := (others => '0');

	for J in  0 to num_stores-1 loop
		if(sr_req_in(J) = '1') then
			curr_time_stamp_var := 
				sr_time_stamp_in (((J+1)*time_stamp_width)-1 downto
								J*time_stamp_width);
			if((none_valid_so_far = '1') or
				IsGreaterThan(smallest_time_stamp_var,
							curr_time_stamp_var)) then
				none_valid_so_far := '0';
				smallest_time_stamp_var := curr_time_stamp_var;
				store_request_id_var := to_unsigned(J, c_store_port_id_width);
				store_request_selected_var := '1';
				store_request_address_var := 
					sr_addr_in(((J+1)*addr_width)-1 downto J*addr_width);
				store_request_data_var := 
					sr_data_in(((J+1)*data_width)-1 downto J*data_width);
				store_request_tag_var := 
						sr_tag_in(((J+1)*tag_width)-1 downto J*tag_width);
			end if;
		end if;
	end loop;
	
	store_request_selected <= store_request_selected_var;
	store_request_id <= store_request_id_var;
	store_request_address <= store_request_address_var;
	store_request_data <= store_request_data_var;
	store_request_tag <= store_request_tag_var;
	store_request_time_stamp <= smallest_time_stamp_var;
  end process;

  srr_data_in <= store_request_time_stamp & 
			to_slv(store_request_id) &  
			store_request_address & store_request_data & store_request_tag;
  store_request_time_stamp_repeated <= 
			srr_data_out((time_stamp_width + c_store_port_id_width + 
							addr_width+data_width+tag_width)-1 downto 
					(c_store_port_id_width + addr_width+data_width + tag_width));
  store_request_id_repeated <= to_unsigned(srr_data_out((c_store_port_id_width + 
							addr_width+data_width+tag_width)-1 downto 
							(addr_width+data_width + tag_width)));
  store_request_address_repeated <= srr_data_out((addr_width+data_width+tag_width)-1 downto 
							(data_width + tag_width));
  store_request_data_repeated <= srr_data_out((data_width+tag_width)-1 downto tag_width);
  store_request_tag_repeated  <= srr_data_out(tag_width-1 downto 0);

  srr : QueueBase
		generic map (name => name & ":srr", 
				queue_depth => 2,
				data_width => (time_stamp_width + c_store_port_id_width +
						addr_width + data_width + tag_width))
		port map (clk => clock, reset => reset,
				data_in => srr_data_in,
				data_out => srr_data_out,
				push_req =>  store_request_selected,
				push_ack =>  store_request_accepted,
				pop_req  =>  store_request_accepted_repeated,
				pop_ack  =>  store_request_selected_repeated);	

  loadReqAcceptGen: for L in 0 to num_loads-1 generate
	lr_ack_out(L) <= '1' when ((load_request_selected = '1')  and 
						(load_request_accepted = '1')
					and (load_request_id = to_unsigned(L, c_load_port_id_width))) else '0';
  end generate loadReqAcceptGen;

  storeReqAcceptGen: for S in 0 to num_stores-1 generate
	sr_ack_out(S) <= '1' when ((store_request_selected = '1')  and 
						(store_request_accepted = '1')
					and (store_request_id = to_unsigned(S,c_store_port_id_width))) else '0';
  end generate storeReqAcceptGen;

  -----------------------------------------------------------------------------
  -- stage 2: memory access through memory bank.
  -----------------------------------------------------------------------------
  DebugGen: if (global_debug_flag) generate
      process(clock)
      begin
	if(clock'event and clock='1') then
		if(reset = '0') then
			if((store_request_selected_repeated = '1') and
				(store_request_accepted_repeated = '1'))  then
				assert false report
				"MS:" & name & "STORE TS=" & 
					Convert_Integer_To_String(To_Integer(store_request_time_stamp_repeated)) & 
		" ADDR=" & Convert_To_String(store_request_address_repeated) & 
		" DATA="  & Convert_To_String(store_request_data_repeated) 
				severity note;
			end if;
			if((load_request_selected_repeated = '1') and
				(load_request_accepted_repeated = '1'))  then
				assert false report
				"MS:" & name & "LOAD  TS=" & 
					Convert_To_String(load_request_time_stamp_repeated) & 
		" ADDR=" & Convert_Integer_To_String(To_Integer(load_request_address_repeated)) 
				severity note;
			end if;
		end if;
	end if;
      end process;
  end generate DebugGen;

  mb: memory_bank_revised
	generic map (name => name & ":memory_bank",
			g_addr_width => addr_width,
			g_data_width => data_width,
			g_write_tag_width => tag_width,
			g_read_tag_width => tag_width,
			g_read_port_id_width => c_load_port_id_width,
			g_write_port_id_width => c_store_port_id_width,
			g_time_stamp_width => time_stamp_width,
     			g_base_bank_addr_width => addr_width,
     			g_base_bank_data_width => data_width)
	port map ( clk => clock, reset => reset,
			write_data => store_request_data_repeated,
			write_addr => store_request_address_repeated,
			write_port_id => store_request_id_repeated,
			write_port_id_out => store_complete_id,
			write_tag  => store_request_tag_repeated,
			write_time_stamp => store_request_time_stamp_repeated,
			write_tag_out => store_complete_tag,
			write_enable => store_request_selected_repeated,
			write_ack => store_request_accepted_repeated,
			write_result_ready => store_complete_ready,
			write_result_accept => store_complete_accept,
			read_data => load_complete_data,
			read_addr => load_request_address_repeated,
			read_tag =>  load_request_tag_repeated,
			read_time_stamp => load_request_time_stamp_repeated,
			read_tag_out => load_complete_tag,
			read_port_id => load_request_id_repeated,
			read_port_id_out => load_complete_id,
			read_enable => load_request_selected_repeated,
			read_ack => load_request_accepted_repeated,
			read_result_ready => load_complete_ready,
			read_result_accept => load_complete_accept);
			

  -----------------------------------------------------------------------------
  -- stage 3:  write to appropriate destination.
  -----------------------------------------------------------------------------
  load_complete_accept <= OrReduce(load_complete_accept_array);
  loadCompleteAcceptGen: for CL in 0 to num_loads-1 generate
    llogic: block
	signal pop_req,pop_ack,push_req,push_ack: std_logic;
	signal rdata_in, rdata_out: std_logic_vector((data_width+tag_width)-1 downto 0);
    begin
	lnr: NullRepeater  -- a place-holder
		generic map (name => name & ":lfrr",
				data_width => (data_width + tag_width))
		port map (clk => clock, reset => reset,
				data_in => rdata_in,
				data_out => rdata_out,
				push_req => push_req,
				push_ack => push_ack,
				pop_req => pop_req,
				pop_ack => pop_ack);
				
	
	rdata_in <= load_complete_data & load_complete_tag;
	push_req <= '1' when ((load_complete_ready = '1') 
					and (load_complete_id = to_unsigned(CL,c_load_port_id_width)))
						else '0';
	load_complete_accept_array(CL) <= push_ack when 
				(load_complete_id = to_unsigned(CL,c_load_port_id_width)) else '0';

	pop_req <= lc_req_in(CL);
	lc_ack_out(CL) <= pop_ack;

	lc_data_out(((CL+1)*data_width)-1 downto CL*data_width) 
		<= rdata_out((data_width + tag_width)-1 downto tag_width);
	lc_tag_out(((CL+1)*tag_width)-1 downto CL*tag_width) <= rdata_out(tag_width-1 downto 0);
     end block;
  end generate loadCompleteAcceptGen;

  store_complete_accept <= OrReduce(store_complete_accept_array);
  storeCompleteAcceptGen: for CS in 0 to num_stores-1 generate
    slogic: block
	signal pop_req,pop_ack,push_req,push_ack: std_logic;
	signal rdata_in, rdata_out: std_logic_vector(tag_width-1 downto 0);
    begin
	snr: NullRepeater 
		generic map (name => name & ":sfrr",
				data_width => tag_width)
		port map (clk => clock, reset => reset,
				data_in => rdata_in,
				data_out => rdata_out,
				push_req => push_req,
				push_ack => push_ack,
				pop_req => pop_req,
				pop_ack => pop_ack);

	rdata_in <= store_complete_tag;
	push_req <= '1' when ((store_complete_ready = '1') 
					and (store_complete_id = to_unsigned(CS, c_store_port_id_width)))
					 else '0';
	store_complete_accept_array(CS) <= push_ack when 
				(store_complete_id = to_unsigned(CS, c_store_port_id_width)) else '0';

	pop_req <= sc_req_in(CS);
	sc_ack_out(CS) <= pop_ack;

	sc_tag_out(((CS+1)*tag_width)-1 downto CS*tag_width) <= rdata_out;

     end block;
  end generate storeCompleteAcceptGen;

end pipelined;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

-- memory subsystem guarantees that accesses to the same location
-- will take place in the order of the time-stamp assigned to each
-- access (tie breaks will be random). Time-stamp is set at the
-- point of acceptance of an access request.

entity memory_subsystem is
  generic(name: string;
	  num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          number_of_banks       : natural := 1;
          mux_degree            : natural := 10;
          demux_degree          : natural := 10;
	  base_bank_addr_width  : natural := 8;
	  base_bank_data_width  : natural := 8);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity memory_subsystem;


architecture bufwrap of memory_subsystem is

  constant time_stamp_width : natural := 2 + Ceil_Log2(num_loads + num_stores);   --  two msb bits for identification
  
  signal lr_addr_in_core :std_logic_vector((num_loads*addr_width)-1 downto 0);
  signal lr_req_in_core  :std_logic_vector(num_loads-1 downto 0);
  signal lr_ack_out_core :std_logic_vector(num_loads-1 downto 0);
  signal lr_tag_in_core :std_logic_vector((num_loads*tag_width)-1 downto 0);
  signal lr_time_stamp_in_core :std_logic_vector((num_loads*time_stamp_width)-1 downto 0);  

  signal sr_addr_in_core :std_logic_vector((num_stores*addr_width)-1 downto 0);
  signal sr_data_in_core :std_logic_vector((num_stores*data_width)-1 downto 0);
  signal sr_req_in_core  : std_logic_vector(num_stores-1 downto 0);
  signal sr_ack_out_core : std_logic_vector(num_stores-1 downto 0);
  signal sr_tag_in_core :std_logic_vector((num_stores*tag_width)-1 downto 0);
  signal sr_time_stamp_in_core :std_logic_vector((num_stores*time_stamp_width)-1 downto 0);
  

  type LoadRepeaterData is array (natural range <> ) of std_logic_vector(time_stamp_width+addr_width+tag_width - 1 downto 0);
  type StoreRepeaterData is array (natural range <> ) of std_logic_vector(time_stamp_width+data_width+addr_width+tag_width - 1 downto 0);
  signal load_repeater_data_in, load_repeater_data_out: LoadRepeaterData(0 to num_loads-1);
  signal store_repeater_data_in, store_repeater_data_out: StoreRepeaterData(0 to num_stores-1);

  signal raw_time_stamp: std_logic_vector(time_stamp_width-1 downto 0);

begin

  -----------------------------------------------------------------------------
  -- time-stamp generation
  -----------------------------------------------------------------------------

  process(clock,reset)
  begin

    if clock'event and clock = '1' then
      if(reset = '1') then
        raw_time_stamp <= (others => '0');
      else
        raw_time_stamp <= IncrementSLV(raw_time_stamp);
      end if;
    end if;
  end process;

  -- instantiate repeaters for each load and store input
  LoadRepGen: for LOAD in 0 to num_loads-1 generate

    load_repeater_data_in(LOAD) <= raw_time_stamp &
                                   lr_addr_in((LOAD+1)*addr_width-1 downto LOAD*addr_width) &
                                   lr_tag_in((LOAD+1)*tag_width - 1 downto LOAD*tag_width);

    lr_time_stamp_in_core((LOAD+1)*time_stamp_width -1 downto LOAD*time_stamp_width) <=
      load_repeater_data_out(LOAD)(time_stamp_width+addr_width+tag_width-1 downto addr_width+tag_width);
    
    lr_addr_in_core((LOAD+1)*addr_width -1 downto LOAD*addr_width) <=
      load_repeater_data_out(LOAD)(addr_width+tag_width-1 downto tag_width);
    lr_tag_in_core((LOAD+1)*tag_width-1 downto LOAD*tag_width) <= load_repeater_data_out(LOAD)(tag_width-1 downto 0);
    
    Rptr : mem_shift_repeater generic map (
      name => name & "-load-mem-shift-repeater-" & Convert_Integer_To_String(LOAD),
      g_data_width => time_stamp_width+ addr_width + tag_width,
	g_number_of_stages => 0)
      port map (
        clk      => clock,
        reset    => reset,
        data_in  => load_repeater_data_in(LOAD),
        req_in   => lr_req_in(LOAD),
        ack_out  => lr_ack_out(LOAD),
        data_out => load_repeater_data_out(LOAD),
        req_out  => lr_req_in_core(LOAD),
        ack_in   => lr_ack_out_core(LOAD));
    
  end generate LoadRepGen;


  StoreRepGen: for STORE in 0 to num_stores-1 generate
    store_repeater_data_in(STORE) <= raw_time_stamp &
                                     sr_data_in((STORE+1)*data_width-1 downto STORE*data_width) &
                                     sr_addr_in((STORE+1)*addr_width-1 downto STORE*addr_width) &
                                     sr_tag_in((STORE+1)*tag_width - 1 downto STORE*tag_width);

    sr_time_stamp_in_core((STORE+1)*time_stamp_width -1 downto STORE*time_stamp_width) <=
      store_repeater_data_out(STORE)(time_stamp_width+data_width+addr_width+tag_width-1 downto data_width+addr_width+tag_width);
    sr_data_in_core((STORE+1)*data_width -1 downto STORE*data_width) <=
          store_repeater_data_out(STORE)(data_width+addr_width+tag_width-1 downto addr_width+tag_width);
    sr_addr_in_core((STORE+1)*addr_width -1 downto STORE*addr_width) <=
      store_repeater_data_out(STORE)(addr_width+tag_width-1 downto tag_width);
    sr_tag_in_core((STORE+1)*tag_width-1 downto STORE*tag_width) <= store_repeater_data_out(STORE)(tag_width-1 downto 0);
    
    Rptr : mem_shift_repeater generic map (
      name => name & "-store-mem-shift-repeater-" & Convert_Integer_To_String(STORE),
      g_data_width => time_stamp_width+data_width + addr_width + tag_width,
      g_number_of_stages => 0)
      port map (
        clk      => clock,
        reset    => reset,
        data_in  => store_repeater_data_in(STORE),
        req_in   => sr_req_in(STORE),
        ack_out  => sr_ack_out(STORE),
        data_out => store_repeater_data_out(STORE),
        req_out  => sr_req_in_core(STORE),
        ack_in   => sr_ack_out_core(STORE));
    
  end generate StoreRepGen;

  core: memory_subsystem_core
    generic map (
      name => name & "-core",
      num_loads            => num_loads,
      num_stores           => num_stores,
      addr_width           => addr_width,
      data_width           => data_width,
      tag_width            => tag_width,
      time_stamp_width     => time_stamp_width,
      number_of_banks      => number_of_banks,
      mux_degree           => mux_degree,
      demux_degree         => demux_degree,
      base_bank_addr_width => base_bank_addr_width,
      base_bank_data_width => base_bank_data_width)
    port map (
      lr_addr_in  => lr_addr_in_core,
      lr_req_in   => lr_req_in_core,
      lr_ack_out  => lr_ack_out_core,
      lr_tag_in   => lr_tag_in_core,
      lr_time_stamp_in => lr_time_stamp_in_core,
      lc_data_out => lc_data_out,
      lc_req_in   => lc_req_in,
      lc_ack_out  => lc_ack_out,
      lc_tag_out  => lc_tag_out,
      sr_addr_in  => sr_addr_in_core,
      sr_data_in  => sr_data_in_core,
      sr_req_in   => sr_req_in_core,
      sr_ack_out  => sr_ack_out_core,
      sr_tag_in   => sr_tag_in_core,
      sr_time_stamp_in => sr_time_stamp_in_core,      
      sc_ack_out  => sc_ack_out,
      sc_req_in   => sc_req_in,
      sc_tag_out  => sc_tag_out,
      clock       => clock,
      reset       => reset);    
end bufwrap;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;
-- TODO: some bug here.

entity merge_box_with_repeater is 
  generic (name: string;
	   g_data_width: natural := 10;
           g_number_of_inputs: natural := 8;
           g_number_of_outputs: natural := 1;
           g_time_stamp_width : natural := 3;   -- width of timestamp
           g_tag_width : natural := 3;  -- width of tag
           g_pipeline_flag: integer := 1     -- if 0, dont add pipe-line stage
           );            

  port(data_left: in  std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
       req_in : in std_logic_vector(g_number_of_inputs-1 downto 0);
       ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
       data_right: out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
       req_out : out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clock: in std_logic;
       reset: in std_logic);

end merge_box_with_repeater;

architecture behave of merge_box_with_repeater is

  constant c_actual_data_width  : natural := g_data_width - g_time_stamp_width;
  constant c_num_inputs_per_tree : natural := Ceiling(g_number_of_inputs,g_number_of_outputs);
  constant c_residual_num_inputs_per_tree : natural := (g_number_of_inputs - ((g_number_of_outputs-1)*c_num_inputs_per_tree));
  
  signal in_data : std_logic_vector((c_actual_data_width*g_number_of_inputs)-1 downto 0);
  signal in_tstamp : std_logic_vector((g_time_stamp_width*g_number_of_inputs)-1 downto 0);
  signal in_req,in_ack : std_logic_vector(g_number_of_inputs-1 downto 0);
  signal out_req,out_ack : std_logic_vector(g_number_of_outputs-1 downto 0);
  signal out_data : std_logic_vector((g_number_of_outputs*c_actual_data_width)-1 downto 0);
  signal out_tstamp : std_logic_vector((g_number_of_outputs*g_time_stamp_width)-1 downto 0);
  
  signal repeater_in, repeater_out : std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0);
  signal repeater_in_req,repeater_in_ack,repeater_out_req,repeater_out_ack : std_logic_vector(g_number_of_outputs-1 downto 0);

  function RepeaterShiftDelay (constant x : integer)
    return integer is
    variable ret_var :integer;
  begin
    ret_var := 0;
    if(x > 0) then
      ret_var := 1;
    end if;
    return(ret_var);
  end RepeaterShiftDelay;
  constant shift_delay : integer := RepeaterShiftDelay(g_pipeline_flag);
  
begin  -- behave

  assert g_number_of_inputs > 0 and g_number_of_outputs > 0 report "at least one i/p and o/p needed in merge-box with repeater" severity error;
  
  -- unpack input-side signals.
  genIn: for I in 0 to g_number_of_inputs-1 generate
    in_data((c_actual_data_width*(I+1))-1 downto (c_actual_data_width*I)) <=
      data_left((g_data_width*(I+1) -1) downto ((g_data_width*(I+1))-c_actual_data_width));
    in_tstamp((g_time_stamp_width*(I+1))-1 downto (g_time_stamp_width*I)) <=
      data_left(((g_data_width*(I+1) - c_actual_data_width) - 1) downto (g_data_width*I));
    in_req(I) <= req_in(I);
    ack_out(I) <= in_ack(I);
  end generate genIn;

  -- unpack output side signals.
  genOut: for I in 0 to g_number_of_outputs-1 generate
    repeater_in((g_data_width)*(I+1)-1 downto ((g_data_width)*I))
      <= out_data((c_actual_data_width*(I+1))-1 downto (c_actual_data_width*I)) &
           out_tstamp((g_time_stamp_width*(I+1))-1 downto (g_time_stamp_width*I));

    repeater_in_req(I) <= out_req(I);
    out_ack(I) <= repeater_in_ack(I);
    
    data_right((g_data_width*(I+1))-1 downto (g_data_width*I)) <=
          repeater_out((g_data_width)*(I+1)-1 downto ((g_data_width)*I));
    req_out(I) <= repeater_out_req(I);
    repeater_out_ack(I) <= ack_in(I);
  end generate genOut;

  -- now instantiate the comb.merge block followed by the
  -- repeater.
  ifgen: if g_number_of_outputs > 1 generate
    
    genLogic: for J in 0 to g_number_of_outputs-2 generate

      cmerge: combinational_merge
        generic map(name => name & "-cmerge" & Convert_Integer_To_String(J), 
		    g_data_width        => c_actual_data_width,
                    g_number_of_inputs  => c_num_inputs_per_tree,
                    g_time_stamp_width  => g_time_stamp_width)
        port map(in_data    => in_data    (((J+1)*c_num_inputs_per_tree*c_actual_data_width)-1
                                           downto
                                           (J*c_num_inputs_per_tree*c_actual_data_width)),
                 in_tstamp  => in_tstamp  (((J+1)*c_num_inputs_per_tree*g_time_stamp_width)-1
                                           downto
                                           (J*c_num_inputs_per_tree*g_time_stamp_width)),
                 out_data   => out_data   ((J+1)*(c_actual_data_width)-1 downto (J*c_actual_data_width)),
                 out_tstamp => out_tstamp ((J+1)*(g_time_stamp_width)-1 downto (J*g_time_stamp_width)),
                 in_req     => in_req     (((J+1)*c_num_inputs_per_tree)-1 downto (J*c_num_inputs_per_tree)),
                 in_ack     => in_ack     (((J+1)*c_num_inputs_per_tree)-1 downto (J*c_num_inputs_per_tree)),
                 out_req    => out_req    (J),
                 out_ack    => out_ack    (J));

      Rptr: mem_shift_repeater generic map(name => name & "-Rptr",
						g_data_width => g_data_width, g_number_of_stages => shift_delay)
        port map(clk      => clock,
                 reset    => reset,
                 data_in  => repeater_in      ((J+1)*(g_data_width) -1 downto (J*(g_data_width))),
                 req_in   => repeater_in_req  (J),
                 ack_out  => repeater_in_ack  (J),
                 data_out => repeater_out     ((J+1)*(g_data_width) -1 downto (J*(g_data_width))),
                 req_out  => repeater_out_req (J),
                 ack_in   => repeater_out_ack (J));
      
    end generate genLogic;
  end generate ifgen;


  -- residual block
  cmerge: combinational_merge
    generic map(name => name & "-residual-cmerge", g_data_width        => c_actual_data_width,
                g_number_of_inputs  => c_residual_num_inputs_per_tree,
                g_time_stamp_width  => g_time_stamp_width)
    port map(in_data    => in_data    ((g_number_of_inputs*c_actual_data_width-1) downto
                                       ((g_number_of_inputs*c_actual_data_width) -
                                        (c_residual_num_inputs_per_tree*c_actual_data_width))),
             in_tstamp  => in_tstamp  ((g_number_of_inputs*g_time_stamp_width-1) downto
                                       ((g_number_of_inputs*g_time_stamp_width) -
                                        (c_residual_num_inputs_per_tree*g_time_stamp_width))),
             out_data   => out_data   ((g_number_of_outputs)*(c_actual_data_width)-1 downto
                                       ((g_number_of_outputs-1)*c_actual_data_width)),
             out_tstamp => out_tstamp ((g_number_of_outputs)*(g_time_stamp_width)-1 downto
                                       ((g_number_of_outputs-1)*g_time_stamp_width)),
             in_req     => in_req     (g_number_of_inputs-1 downto
                                       (g_number_of_inputs - c_residual_num_inputs_per_tree)),
             in_ack     => in_ack     (g_number_of_inputs-1 downto
                                       (g_number_of_inputs - c_residual_num_inputs_per_tree)),
             out_req    => out_req    (g_number_of_outputs-1),
             out_ack    => out_ack    (g_number_of_outputs-1));

  -- residual repeater
  Rptr: mem_shift_repeater generic map(name => name & "-residual-Rptr", g_data_width => g_data_width, g_number_of_stages => shift_delay)
    port map(clk      => clock,
             reset    => reset,
             data_in  => repeater_in      ((g_number_of_outputs)*(g_data_width) -1 downto ((g_number_of_outputs-1)*(g_data_width))),
             req_in   => repeater_in_req  (g_number_of_outputs-1),
             ack_out  => repeater_in_ack  (g_number_of_outputs-1),
             data_out => repeater_out     ((g_number_of_outputs)*(g_data_width) -1 downto ((g_number_of_outputs-1)*(g_data_width))),
             req_out  => repeater_out_req (g_number_of_outputs-1),
             ack_in   => repeater_out_ack (g_number_of_outputs-1));

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity merge_tree is
  generic (
    name: string;
    g_number_of_inputs: natural;          
    g_data_width: natural;          -- total width of data
                                        -- (= actual-data & timestamp)
    g_time_stamp_width : natural ;   -- width of timestamp
    g_tag_width : natural;          -- width of tag
    g_mux_degree :natural;         -- max-indegree of each pipeline-stage
    g_num_stages: natural ;
    g_port_id_width: natural
    );       

  port (
    merge_data_in : in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    merge_req_in  : in std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_data_out: out std_logic_vector(g_data_width-1 downto 0);
    merge_req_out : out std_logic;
    merge_ack_in  : in std_logic;
    clock: in std_logic;
    reset: in std_logic);
  
end merge_tree;


architecture pipelined of merge_tree is
  constant c_number_of_stages : integer := Maximum(1,Ceil_Log(g_number_of_inputs, g_mux_degree));
  constant c_residual_num_stages : integer := Maximum(0,g_num_stages - c_number_of_stages);
  constant c_total_intermediate_width : natural := Total_Intermediate_Width(g_number_of_inputs,g_mux_degree);

  -- intermediate signals used to cross levels.
  signal intermediate_vector : std_logic_vector(0 to ((g_data_width)*c_total_intermediate_width)-1);  
  signal intermediate_req_vector : std_logic_vector(0 to (c_total_intermediate_width)-1);
  signal intermediate_ack_vector : std_logic_vector(0 to (c_total_intermediate_width)-1);

begin  -- behave
  assert g_num_stages >= c_number_of_stages report "requested number of stages should be >= number of stages implied by mux-degree" severity error;
  assert Stage_Width(c_number_of_stages,g_mux_degree, g_number_of_inputs) = 1 report "last stage should have one input!" severity error;
  
  intermediate_vector(
    Left_Index(0,g_mux_degree,g_number_of_inputs)*g_data_width to
    ((Right_Index(0,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1)
    <= merge_data_in;

  intermediate_req_vector(
    Left_Index(0,g_mux_degree,g_number_of_inputs) to
    Right_Index(0,g_mux_degree,g_number_of_inputs))
    <= merge_req_in;

  merge_ack_out <=
    intermediate_ack_vector(
      Left_Index(0,g_mux_degree,g_number_of_inputs) to
      Right_Index(0,g_mux_degree,g_number_of_inputs));

  PipelineGen:  for LEVEL  in 0 to c_number_of_stages-1  generate

    -- mbox with repeater has multiple outputs, with tree driving
    -- each output and repeater present at each output.
    mBoxPipeStage : merge_box_with_repeater generic map (
      name => name & "-mBoxPipeState-" & Convert_To_String(LEVEL),
      g_data_width => g_data_width,
      g_number_of_inputs => Stage_Width(LEVEL,g_mux_degree,g_number_of_inputs),
      g_number_of_outputs => Stage_Width(LEVEL+1,g_mux_degree,g_number_of_inputs),
      g_time_stamp_width => g_time_stamp_width,
      g_tag_width => g_tag_width,
      g_pipeline_flag => c_number_of_stages-1 )
      port map ( data_left =>
                 intermediate_vector(
                   Left_Index(LEVEL,g_mux_degree,g_number_of_inputs)*g_data_width to
                   ((Right_Index(LEVEL,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1),
                 req_in =>
                 intermediate_req_vector(
                   Left_Index(LEVEL,g_mux_degree,g_number_of_inputs) to
                   Right_Index(LEVEL,g_mux_degree,g_number_of_inputs)),
                 ack_out =>
                   intermediate_ack_vector(
                     Left_Index(LEVEL,g_mux_degree,g_number_of_inputs) to
                     Right_Index(LEVEL,g_mux_degree,g_number_of_inputs)),
                 data_right =>
                 intermediate_vector(
                   Left_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)*g_data_width to
                   ((Right_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1),
                 req_out =>
                 intermediate_req_vector(
                   Left_Index(LEVEL+1,g_mux_degree,g_number_of_inputs) to
                   Right_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)),
                 ack_in =>
                   intermediate_ack_vector(
                     Left_Index(LEVEL+1,g_mux_degree,g_number_of_inputs) to
                     Right_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)),
                 clock => clock,
                 reset => reset);
                   
  end generate;  -- PipelineGen

  -- to the right (pad the required number of shifts)
  finalRptr : mem_shift_repeater generic map (
    name => name & "-finalRptr",
    g_data_width => g_data_width,
    g_number_of_stages => c_residual_num_stages)
    port map (
      clk     => clock,
      reset   => reset,
      data_in => intermediate_vector(
        Left_Index(c_number_of_stages,g_mux_degree,g_number_of_inputs)*g_data_width to
        ((Right_Index(c_number_of_stages,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1),
      req_in => intermediate_req_vector(Left_Index(c_number_of_stages,g_mux_degree, g_number_of_inputs)),
      ack_out =>   intermediate_ack_vector(Left_Index(c_number_of_stages,g_mux_degree, g_number_of_inputs)),
      data_out => merge_data_out,
      req_out => merge_req_out,
      ack_in => merge_ack_in);
end pipelined;

architecture combinational_arch of merge_tree is
  constant actual_data_width : natural := g_data_width - (g_time_stamp_width);
  signal data_sig : std_logic_vector(g_number_of_inputs*actual_data_width-1 downto 0);

  signal out_data_sig : std_logic_vector(actual_data_width-1 downto 0);
  signal out_tstamp_sig : std_logic_vector(g_time_stamp_width-1 downto 0);
  signal tstamp_sig : std_logic_vector(g_number_of_inputs*g_time_stamp_width -1  downto 0);
  
begin  
  assert g_data_width > g_time_stamp_width report "data width smaller than time-stamp in merge?" severity error;
  packGen: for P in 0 to g_number_of_inputs-1 generate
    data_sig((P+1)*actual_data_width-1 downto P*actual_data_width) <=
      merge_data_in((P+1)*g_data_width-1 downto (P+1)*g_data_width - (actual_data_width));
    tstamp_sig((P+1)*g_time_stamp_width-1 downto P*g_time_stamp_width) <=
      merge_data_in((P*g_data_width)+g_time_stamp_width-1 downto P*g_data_width);
  end generate packGen;

  cMerge : combinational_merge generic map (
    name => name & ":cMerge:", 
    g_data_width       => actual_data_width,
    g_number_of_inputs => g_number_of_inputs,
    g_time_stamp_width => g_time_stamp_width)
    port map (
      in_data    => data_sig,
      out_data   => out_data_sig,
      in_tstamp  => tstamp_sig,
      out_tstamp => out_tstamp_sig,
      in_req     => merge_req_in,
      in_ack     => merge_ack_out,
      out_req    => merge_req_out,
      out_ack    => merge_ack_in);

  merge_data_out <= out_data_sig & out_tstamp_sig;
end combinational_arch;
  
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

-- memory subsystem guarantees that accesses to the same location
-- will take place in the order of the time-stamp assigned to each
-- access (tie breaks will be random). Time-stamp is set at the
-- point of acceptance of an access request.

entity ordered_memory_subsystem is
  generic(name: string;
	  num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          time_stamp_width      : natural := 0;
          number_of_banks       : natural := 1;
          mux_degree            : natural := 10;
          demux_degree          : natural := 10;
	  base_bank_addr_width  : natural := 8;
	  base_bank_data_width  : natural := 8);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag + timestamp: tag will be returned on completion..
    lr_tag_in: in std_logic_vector((num_loads*(tag_width+time_stamp_width))-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*(tag_width+time_stamp_width))-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity ordered_memory_subsystem;


architecture bufwrap of ordered_memory_subsystem is

  
  signal lr_addr_in_core :std_logic_vector((num_loads*addr_width)-1 downto 0);
  signal lr_req_in_core  :std_logic_vector(num_loads-1 downto 0);
  signal lr_ack_out_core :std_logic_vector(num_loads-1 downto 0);
  signal lr_tag_in_core :std_logic_vector((num_loads*tag_width)-1 downto 0);
  signal lr_time_stamp_in_core :std_logic_vector((num_loads*time_stamp_width)-1 downto 0);  

  signal sr_addr_in_core :std_logic_vector((num_stores*addr_width)-1 downto 0);
  signal sr_data_in_core :std_logic_vector((num_stores*data_width)-1 downto 0);
  signal sr_req_in_core  : std_logic_vector(num_stores-1 downto 0);
  signal sr_ack_out_core : std_logic_vector(num_stores-1 downto 0);
  signal sr_tag_in_core :std_logic_vector((num_stores*tag_width)-1 downto 0);
  signal sr_time_stamp_in_core :std_logic_vector((num_stores*time_stamp_width)-1 downto 0);
  

  type LoadRepeaterData is array (natural range <> ) of std_logic_vector(time_stamp_width+addr_width+tag_width - 1 downto 0);
  type StoreRepeaterData is array (natural range <> ) of std_logic_vector(time_stamp_width+data_width+addr_width+tag_width - 1 downto 0);
  signal load_repeater_data_in, load_repeater_data_out: LoadRepeaterData(0 to num_loads-1);
  signal store_repeater_data_in, store_repeater_data_out: StoreRepeaterData(0 to num_stores-1);

  signal raw_time_stamp: std_logic_vector(time_stamp_width-1 downto 0);

begin


  ifMoreThanOneLoad: if num_loads > 1 generate
  -- instantiate repeaters for each load and store input
  LoadRepGen: for LOAD in 0 to num_loads-1 generate


    load_repeater_data_in(LOAD) <= lr_addr_in((LOAD+1)*addr_width-1 downto LOAD*addr_width) &
                                   lr_tag_in((LOAD+1)*(tag_width+time_stamp_width) - 1 downto 
					LOAD*(tag_width+time_stamp_width));

    lr_time_stamp_in_core((LOAD+1)*time_stamp_width -1 downto LOAD*time_stamp_width) <=
      load_repeater_data_out(LOAD)(time_stamp_width-1 downto 0);
    
    lr_addr_in_core((LOAD+1)*addr_width -1 downto LOAD*addr_width) <=
      load_repeater_data_out(LOAD)(addr_width+tag_width+time_stamp_width-1 downto tag_width+time_stamp_width);
    lr_tag_in_core((LOAD+1)*tag_width-1 downto LOAD*tag_width) <= load_repeater_data_out(LOAD)(tag_width+time_stamp_width-1 downto time_stamp_width);
    
    Rptr : mem_shift_repeater generic map (
      name => name & "-load-Rptr-" & Convert_Integer_To_String(LOAD),
      g_data_width => time_stamp_width+ addr_width + tag_width,
	g_number_of_stages => 1)
      port map (
        clk      => clock,
        reset    => reset,
        data_in  => load_repeater_data_in(LOAD),
        req_in   => lr_req_in(LOAD),
        ack_out  => lr_ack_out(LOAD),
        data_out => load_repeater_data_out(LOAD),
        req_out  => lr_req_in_core(LOAD),
        ack_in   => lr_ack_out_core(LOAD));
    
  end generate LoadRepGen;
  end generate ifMoreThanOneLoad;

  onlyOneLoad: if num_loads = 1 generate
      lr_tag_in_core <= lr_tag_in((tag_width+time_stamp_width) - 1 downto  time_stamp_width);
      lr_time_stamp_in_core <= lr_tag_in(time_stamp_width - 1 downto  0);
      lr_req_in_core <= lr_req_in;
      lr_addr_in_core <= lr_addr_in;

      lr_ack_out  <= lr_ack_out_core;
  end generate onlyOneLoad;


  ifMoreThanOneStore: if num_stores > 1 generate
  StoreRepGen: for STORE in 0 to num_stores-1 generate
    store_repeater_data_in(STORE) <= sr_data_in((STORE+1)*data_width-1 downto STORE*data_width) &
                                     sr_addr_in((STORE+1)*addr_width-1 downto STORE*addr_width) &
                                     sr_tag_in((STORE+1)*(tag_width+time_stamp_width) - 1 downto 
						STORE*(tag_width+time_stamp_width));

    sr_time_stamp_in_core((STORE+1)*time_stamp_width -1 downto STORE*time_stamp_width) <=
      store_repeater_data_out(STORE)(time_stamp_width-1 downto 0);
    sr_data_in_core((STORE+1)*data_width -1 downto STORE*data_width) <=
          store_repeater_data_out(STORE)(data_width+addr_width+tag_width+time_stamp_width-1 downto addr_width+tag_width+time_stamp_width);
    sr_addr_in_core((STORE+1)*addr_width -1 downto STORE*addr_width) <=
      store_repeater_data_out(STORE)(addr_width+tag_width+time_stamp_width-1 downto tag_width+time_stamp_width);
    sr_tag_in_core((STORE+1)*tag_width-1 downto STORE*tag_width) <= store_repeater_data_out(STORE)(tag_width+time_stamp_width-1 downto time_stamp_width);
    
    Rptr : mem_shift_repeater generic map (
      name => name & "-store-Rptr-" & Convert_Integer_To_String(STORE),
      g_data_width => time_stamp_width+data_width + addr_width + tag_width,
      g_number_of_stages => 1)
      port map (
        clk      => clock,
        reset    => reset,
        data_in  => store_repeater_data_in(STORE),
        req_in   => sr_req_in(STORE),
        ack_out  => sr_ack_out(STORE),
        data_out => store_repeater_data_out(STORE),
        req_out  => sr_req_in_core(STORE),
        ack_in   => sr_ack_out_core(STORE));
    
  end generate StoreRepGen;
  end generate ifMoreThanOneStore;

  onlyOneStore: if num_stores = 1 generate

      sr_tag_in_core <= sr_tag_in((tag_width+time_stamp_width) - 1 downto  time_stamp_width);
      sr_time_stamp_in_core <= sr_tag_in(time_stamp_width - 1 downto  0);
      sr_req_in_core  <= sr_req_in;
      sr_addr_in_core <= sr_addr_in;
      sr_data_in_core <= sr_data_in;

      sr_ack_out  <= sr_ack_out_core;
  end generate onlyOneStore;

  nonTrivGen: if (num_loads > 0) and (num_stores > 0) generate
  core: memory_subsystem_core
    generic map (
      name => name & "-core",
      num_loads            => num_loads,
      num_stores           => num_stores,
      addr_width           => addr_width,
      data_width           => data_width,
      tag_width            => tag_width,
      time_stamp_width     => time_stamp_width,
      number_of_banks      => number_of_banks,
      mux_degree           => mux_degree,
      demux_degree         => demux_degree,
      base_bank_addr_width => base_bank_addr_width,
      base_bank_data_width => base_bank_data_width)
    port map (
      lr_addr_in  => lr_addr_in_core,
      lr_req_in   => lr_req_in_core,
      lr_ack_out  => lr_ack_out_core,
      lr_tag_in   => lr_tag_in_core,
      lr_time_stamp_in => lr_time_stamp_in_core,
      lc_data_out => lc_data_out,
      lc_req_in   => lc_req_in,
      lc_ack_out  => lc_ack_out,
      lc_tag_out  => lc_tag_out,
      sr_addr_in  => sr_addr_in_core,
      sr_data_in  => sr_data_in_core,
      sr_req_in   => sr_req_in_core,
      sr_ack_out  => sr_ack_out_core,
      sr_tag_in   => sr_tag_in_core,
      sr_time_stamp_in => sr_time_stamp_in_core,      
      sc_ack_out  => sc_ack_out,
      sc_req_in   => sc_req_in,
      sc_tag_out  => sc_tag_out,
      clock       => clock,
      reset       => reset);    
   end generate nonTrivGen;
end bufwrap;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.types.all;
use ahir.utilities.all;
use ahir.subprograms.all;

entity CombinationalMux is
  generic (
    name : string;
    g_data_width       : integer := 32;
    g_number_of_inputs: integer := 2);
  port(
    in_data: in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    out_data: out std_logic_vector(g_data_width-1 downto 0);
    in_req: in std_logic_vector(g_number_of_inputs-1 downto 0);
    in_ack: out std_logic_vector(g_number_of_inputs-1 downto 0);
    out_req: out std_logic;
    out_ack: in std_logic);
end CombinationalMux;

architecture combinational_merge of CombinationalMux is

  signal sel_vector : std_logic_vector(g_number_of_inputs-1 downto 0);
  
begin  -- combinational_merge

  sel_vector <= PriorityEncode(in_req);
  out_req <= OrReduce(in_req);
  in_ack <= sel_vector when out_ack = '1' else (others => '0');



  process(sel_vector,in_data)
  begin
    out_data <= (others => '0');
    for I in 0 to g_number_of_inputs-1 loop
	if(sel_vector(I) = '1') then
	 	out_data <= in_data((g_data_width*(I+1))-1 downto (g_data_width*I));
		exit;
	end if;
    end loop;
  end process;
	   
  
  AckGen: for I in 0 to g_number_of_inputs-1 generate
    in_ack(I) <= '1' when (sel_vector(I) = '1'  and out_ack = '1' and in_req(I) = '1') else '0';
  end generate AckGen;
  
end combinational_merge;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity PipelinedDemux is
  generic ( name: string;
	    g_data_width: natural := 10;
            g_destination_id_width : natural := 3;
            g_number_of_outputs: natural := 8);
  port(data_in: in std_logic_vector(g_data_width-1 downto 0);  -- data & destination-id 
       sel_in : in std_logic_vector(g_destination_id_width-1 downto 0);
       req_in: in std_logic;
       ack_out : out std_logic;
       data_out: out std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0 );
       req_out: out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clk: in std_logic;
       reset: in std_logic);
end entity;

architecture behave of PipelinedDemux is
  type SigArrayType is array (natural range <>) of std_logic_vector(g_data_width-1 downto 0);

  signal data_out_sig,repeater_out_sig : SigArrayType(g_number_of_outputs-1 downto 0);
  signal req_out_sig, ack_in_sig : std_logic_vector(g_number_of_outputs-1 downto 0);
  signal conditioned_ack_in_sig: std_logic_vector(g_number_of_outputs-1 downto 0);

begin  -- behave

  
  conditioned_ack_in_sig <= ack_in_sig and req_out_sig;
  ack_out <= OrReduce(conditioned_ack_in_sig);
    
  gen: for I in 0 to g_number_of_outputs-1 generate

    data_out_sig(I) <= data_in;
    
    process(data_in, sel_in, req_in)
      variable port_index : natural;
    begin
      port_index := To_Integer(sel_in);
      req_out_sig(I) <= '0';
      if(req_in = '1' and port_index = I) then
        req_out_sig(I) <= req_in;
      end if;
    end process;
      
    Repeater : QueueBase generic map(
      				name => name & "-Repeater-" & Convert_Integer_To_String(I),
				queue_depth => 2, data_width => g_data_width)
    port map (
      clk      => clk,
      reset    => reset,
      data_in  => data_out_sig(I),
      push_req  => req_out_sig(I),
      push_ack  => ack_in_sig(I),
      data_out => repeater_out_sig(I),
      pop_ack  => req_out(I),
      pop_Req   => ack_in(I));

    data_out((I+1)*g_data_width -1 downto I*g_data_width) <= repeater_out_sig(I);
  end generate gen;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;
use ahir.BaseComponents.all;

entity PipelinedMuxStage is 
  generic (name: string;
	   g_data_width: integer := 10;
           g_number_of_inputs: integer := 8;
           g_number_of_outputs: integer := 1;
           g_tag_width : integer := 3  -- width of tag
           );            

  port(data_left: in  std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
       req_in : in std_logic_vector(g_number_of_inputs-1 downto 0);
       ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
       data_right: out std_logic_vector((g_data_width*g_number_of_outputs)-1 downto 0);
       req_out : out std_logic_vector(g_number_of_outputs-1 downto 0);
       ack_in : in std_logic_vector(g_number_of_outputs-1 downto 0);
       clock: in std_logic;
       reset: in std_logic);

end PipelinedMuxStage;

architecture behave of PipelinedMuxStage is

  constant c_num_inputs_per_tree : integer := Ceiling(g_number_of_inputs,g_number_of_outputs);
  constant c_residual_num_inputs_per_tree : integer := (g_number_of_inputs - ((g_number_of_outputs-1)*c_num_inputs_per_tree));
  
  signal in_data : std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
  signal in_req,in_ack : std_logic_vector(g_number_of_inputs-1 downto 0);
  signal out_req,out_ack : std_logic_vector(g_number_of_outputs-1 downto 0);
  signal out_data : std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0);
  
  signal repeater_in, repeater_out : std_logic_vector((g_number_of_outputs*g_data_width)-1 downto 0);
  signal repeater_in_req,repeater_in_ack,repeater_out_req,repeater_out_ack : std_logic_vector(g_number_of_outputs-1 downto 0);

  
begin  -- behave

  assert g_number_of_inputs > 0 and g_number_of_outputs > 0 report "at least one i/p and o/p needed in merge-box with repeater" severity error;
  
  -- unpack input-side signals.
  genIn: for I in 0 to g_number_of_inputs-1 generate
    in_data((g_data_width*(I+1))-1 downto (g_data_width*I)) <=
      data_left((g_data_width*(I+1) -1) downto (g_data_width*I));
    in_req(I) <= req_in(I);
    ack_out(I) <= in_ack(I);
  end generate genIn;

  -- unpack output side signals.
  genOut: for I in 0 to g_number_of_outputs-1 generate
    repeater_in((g_data_width)*(I+1)-1 downto ((g_data_width)*I))
      <= out_data((g_data_width*(I+1))-1 downto (g_data_width*I));
    repeater_in_req(I) <= out_req(I);
    out_ack(I) <= repeater_in_ack(I);
    
    data_right((g_data_width*(I+1))-1 downto (g_data_width*I)) <=
          repeater_out((g_data_width)*(I+1)-1 downto ((g_data_width)*I));
    req_out(I) <= repeater_out_req(I);
    repeater_out_ack(I) <= ack_in(I);
  end generate genOut;

  -- now instantiate the comb.merge block followed by the
  -- repeater.
  ifgen: if g_number_of_outputs > 1 generate
    
    genLogic: for J in 0 to g_number_of_outputs-2 generate

      cmerge: CombinationalMux
        generic map(name => name & "-cmerge-" & Convert_Integer_To_String(J), 
		    g_data_width        => g_data_width,
                    g_number_of_inputs  => c_num_inputs_per_tree)
        port map(in_data    => in_data    (((J+1)*c_num_inputs_per_tree*g_data_width)-1
                                           downto
                                           (J*c_num_inputs_per_tree*g_data_width)),
                 out_data   => out_data   ((J+1)*(g_data_width)-1 downto (J*g_data_width)),
                 in_req     => in_req     (((J+1)*c_num_inputs_per_tree)-1 downto (J*c_num_inputs_per_tree)),
                 in_ack     => in_ack     (((J+1)*c_num_inputs_per_tree)-1 downto (J*c_num_inputs_per_tree)),
                 out_req    => out_req    (J),
                 out_ack    => out_ack    (J));

      Rptr: QueueBase generic map(name => name & "-Rptr-" & Convert_Integer_To_String(J),
		  			queue_depth => 2, data_width => g_data_width)
        port map(clk      => clock,
                 reset    => reset,
                 data_in  => repeater_in      ((J+1)*(g_data_width) -1 downto (J*(g_data_width))),
                 push_req   => repeater_in_req  (J),
                 push_ack  => repeater_in_ack  (J),
                 data_out => repeater_out     ((J+1)*(g_data_width) -1 downto (J*(g_data_width))),
                 pop_ack  => repeater_out_req (J),
                 pop_req   => repeater_out_ack (J));
      
    end generate genLogic;
  end generate ifgen;


  -- residual block
  cmerge: CombinationalMux
    generic map(name => name & "-cmerge-residual",
		g_data_width        => g_data_width,
                g_number_of_inputs  => c_residual_num_inputs_per_tree)
    port map(in_data    => in_data    ((g_number_of_inputs*g_data_width-1) downto
                                       ((g_number_of_inputs*g_data_width) -
                                        (c_residual_num_inputs_per_tree*g_data_width))),
             out_data   => out_data   ((g_number_of_outputs)*(g_data_width)-1 downto
                                       ((g_number_of_outputs-1)*g_data_width)),
             in_req     => in_req     (g_number_of_inputs-1 downto
                                       (g_number_of_inputs - c_residual_num_inputs_per_tree)),
             in_ack     => in_ack     (g_number_of_inputs-1 downto
                                       (g_number_of_inputs - c_residual_num_inputs_per_tree)),
             out_req    => out_req    (g_number_of_outputs-1),
             out_ack    => out_ack    (g_number_of_outputs-1));

  -- residual repeater
  Rptr: QueueBase generic map(name => name & "-Rptr-residual",
				queue_depth => 2, data_width => g_data_width)
    port map(clk      => clock,
             reset    => reset,
             data_in  => repeater_in      ((g_number_of_outputs)*(g_data_width) -1 downto ((g_number_of_outputs-1)*(g_data_width))),
             push_req   => repeater_in_req  (g_number_of_outputs-1),
             push_ack  => repeater_in_ack  (g_number_of_outputs-1),
             data_out => repeater_out     ((g_number_of_outputs)*(g_data_width) -1 downto ((g_number_of_outputs-1)*(g_data_width))),
             pop_ack  => repeater_out_req (g_number_of_outputs-1),
             pop_req   => repeater_out_ack (g_number_of_outputs-1));

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;


library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

entity PipelinedMux is
  generic (
    name : string;
    g_number_of_inputs: natural;          
    g_data_width: natural;          -- total width of data
                                        -- (= actual-data & tag & port_id)
    g_mux_degree :natural;         -- max-indegree of each pipeline-stage
    g_port_id_width: natural
    );       

  port (
    merge_data_in : in std_logic_vector((g_data_width*g_number_of_inputs)-1 downto 0);
    merge_req_in  : in std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_ack_out : out std_logic_vector(g_number_of_inputs-1 downto 0);
    merge_data_out: out std_logic_vector(g_data_width-1 downto 0);
    merge_req_out : out std_logic;
    merge_ack_in  : in std_logic;
    clock: in std_logic;
    reset: in std_logic);
  
end PipelinedMux;


architecture pipelined of PipelinedMux is
  constant c_number_of_stages : integer := Maximum(1,Ceil_Log(g_number_of_inputs, g_mux_degree));
  constant c_total_intermediate_width : natural := Total_Intermediate_Width(g_number_of_inputs,g_mux_degree);

  -- intermediate signals used to cross levels.
  signal intermediate_vector : std_logic_vector(0 to ((g_data_width)*c_total_intermediate_width)-1);  
  signal intermediate_req_vector : std_logic_vector(0 to (c_total_intermediate_width)-1);
  signal intermediate_ack_vector : std_logic_vector(0 to (c_total_intermediate_width)-1);

begin  -- behave

  assert Stage_Width(c_number_of_stages,g_mux_degree, g_number_of_inputs) = 1 report "last stage should have one input!" severity error;
  
  intermediate_vector(
    Left_Index(0,g_mux_degree,g_number_of_inputs)*g_data_width to
    ((Right_Index(0,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1)
    <= merge_data_in;

  intermediate_req_vector(
    Left_Index(0,g_mux_degree,g_number_of_inputs) to
    Right_Index(0,g_mux_degree,g_number_of_inputs))
    <= merge_req_in;

  merge_ack_out <=
    intermediate_ack_vector(
      Left_Index(0,g_mux_degree,g_number_of_inputs) to
      Right_Index(0,g_mux_degree,g_number_of_inputs));

  PipelineGen:  for LEVEL  in 0 to c_number_of_stages-1  generate

    -- Each stage has multiple inputs and multiple outputs..
    mBoxPipeStage : PipelinedMuxStage generic map (
      name => name & "-mBoxPipeState-" & Convert_Integer_To_String(LEVEL),
      g_data_width => g_data_width,
      g_number_of_inputs => Stage_Width(LEVEL,g_mux_degree,g_number_of_inputs),
      g_number_of_outputs => Stage_Width(LEVEL+1,g_mux_degree,g_number_of_inputs))
      port map ( data_left =>
                 intermediate_vector(
                   Left_Index(LEVEL,g_mux_degree,g_number_of_inputs)*g_data_width to
                   ((Right_Index(LEVEL,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1),
                 req_in =>
                 intermediate_req_vector(
                   Left_Index(LEVEL,g_mux_degree,g_number_of_inputs) to
                   Right_Index(LEVEL,g_mux_degree,g_number_of_inputs)),
                 ack_out =>
                   intermediate_ack_vector(
                     Left_Index(LEVEL,g_mux_degree,g_number_of_inputs) to
                     Right_Index(LEVEL,g_mux_degree,g_number_of_inputs)),
                 data_right =>
                 intermediate_vector(
                   Left_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)*g_data_width to
                   ((Right_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1),
                 req_out =>
                 intermediate_req_vector(
                   Left_Index(LEVEL+1,g_mux_degree,g_number_of_inputs) to
                   Right_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)),
                 ack_in =>
                   intermediate_ack_vector(
                     Left_Index(LEVEL+1,g_mux_degree,g_number_of_inputs) to
                     Right_Index(LEVEL+1,g_mux_degree,g_number_of_inputs)),
                 clock => clock,
                 reset => reset);
                   
  end generate;  -- PipelineGen

  -- to the right (pad the required number of shifts)
  merge_data_out <= intermediate_vector(
        Left_Index(c_number_of_stages,g_mux_degree,g_number_of_inputs)*g_data_width to
        ((Right_Index(c_number_of_stages,g_mux_degree,g_number_of_inputs)+1)*g_data_width)-1);
  merge_req_out <= 
	intermediate_req_vector(Left_Index(c_number_of_stages,g_mux_degree, g_number_of_inputs));
  intermediate_ack_vector(Left_Index(c_number_of_stages,g_mux_degree, g_number_of_inputs)) 
	<= merge_ack_in;


end pipelined;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

-------------------------------------------------------------------------------
-- a simplified version of the memory subsystem to be used
-- when the number of storage locations is small..
--
-- this is equivalent to a num_loads read-port, num_stores write_port
-- register bank.
-------------------------------------------------------------------------------

entity register_bank is
  generic(name: string;
	  num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          num_registers         : natural := 1);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity register_bank;


-- architecture: synchronous R/W.
--               on destination conflict, writer with lowest index wins.
architecture Default_arch of register_bank is
  type DataArray is array (natural range <>) of std_logic_vector(data_width-1 downto 0);
  type AddrArray is array (natural range <>) of std_logic_vector(addr_width-1 downto 0);

  signal register_array : DataArray(num_registers-1 downto 0) := (others => (others => '0'));

  signal lr_ack_flag: std_logic_vector(num_loads-1 downto 0);
  signal sr_ack_flag : std_logic_vector(num_stores-1 downto 0);
  
  signal lc_ack_flag : std_logic_vector(num_loads-1 downto 0);
  signal sc_ack_flag : std_logic_vector(num_stores-1 downto 0);

  signal lc_data_out_sig : std_logic_vector((num_loads*data_width)-1 downto 0);
  signal sc_tag_out_sig : std_logic_vector((num_stores*tag_width)-1 downto 0);
  signal lc_tag_out_sig : std_logic_vector((num_loads*tag_width)-1 downto 0);

  constant zero_addr : std_logic_vector(addr_width-1 downto 0) := (others => '0');
                                                                 
    
begin

  assert(2**addr_width >= num_registers) report "not enough address bits" severity failure;


  -- the read process. fully parallel reads.
  ReadGen: for R in 0 to num_loads-1 generate

    process(clock,lr_req_in,lc_ack_flag,reset,lr_addr_in)
      variable ack_var : std_logic;
      variable index : integer;
                                 
    begin
      ack_var := '0';
      index := 0;
      
      if(lr_req_in(R) = '1') then
        index := To_Integer(lr_addr_in(((R+1)*addr_width)-1 downto R*addr_width));
      end if;
      
      if(lr_req_in(R) = '1' and lc_ack_flag(R) = '0') then
        ack_var := '1';
      end if;
      
      lr_ack_out(R) <= ack_var;
      
      if(clock'event and clock = '1') then
        if(ack_var = '1') then
          assert (index < num_registers) report "index overflow." severity error;
          assert (index >= 0) report "index underflow" severity error;
          
          lc_data_out_sig(((R+1)*data_width)-1 downto R*data_width) <= register_array(index);
          lc_tag_out_sig(((R+1)*tag_width)-1 downto R*tag_width) <=
            lr_tag_in(((R+1)*tag_width)-1 downto R*tag_width);
          
        end if;
        
        if(reset = '1') then
          lc_ack_flag(R) <= '0';
        else
          if(ack_var = '1') then
            lc_ack_flag(R) <= '1';
          elsif lc_ack_flag(R) = '1' and lc_req_in(R) = '1' then
            lc_ack_flag(R) <= '0';
          end if;
        end if;
      end if;
    end process;
    
  end generate ReadGen;
  
  -- the write process
  -- for each register. loop across those who want to write in
  -- and find the lowest index which wins.
  process(clock,
	  reset,
          sr_req_in,
          sr_addr_in,
          sr_data_in,
          sr_tag_in,
          sc_req_in,
          sc_ack_flag,
	  sc_tag_out_sig,
          register_array)
    
    variable sc_ack_set, sc_ack_clear: std_logic_vector(num_stores-1 downto 0);
    variable sr_pending : std_logic_vector(num_registers-1 downto 0);
    
    variable sc_tag_out_var : std_logic_vector((num_stores*tag_width)-1 downto 0);
    variable register_array_var : DataArray(num_registers-1 downto 0);
    
  begin


    sc_ack_set := (others => '0');
    sc_ack_clear := (others => '0');
    sr_pending := (others => '0');

    sc_tag_out_var := sc_tag_out_sig;

    register_array_var := register_array;
    
    
    if(reset = '1') then
      sc_ack_clear := (others => '1');
    end if;
      
    -- for each register.
    for REG  in 0 to num_registers-1 loop
      
      -- writes: for each reg, lowest index succeeds.
      for W in 0 to num_stores-1 loop
        
        -- if W is a store request to this register
        -- and no j
        if(sr_pending(REG) = '0' and
           sr_req_in(W) = '1' and
           sc_ack_flag(W) = '0' and 
           (sr_addr_in(((W+1)*addr_width)-1 downto W*addr_width) = Natural_To_SLV(REG,addr_width)))
        then
          sr_pending(REG) := '1';
          sc_ack_set(W) := '1';
          register_array_var(REG) := sr_data_in(((W+1)*data_width)-1 downto W*data_width);
          sc_tag_out_var(((W+1)*tag_width)-1 downto W*tag_width) :=
            sr_tag_in(((W+1)*tag_width)-1 downto W*tag_width);
          
          exit;
        end if;
      end loop;  -- W
    end loop;  -- REG
    
    -- output latches and registers
    if(clock'event and clock = '1') then
      register_array <= register_array_var;
      sc_tag_out_sig <= sc_tag_out_var;
    end if;
  
    -- lc/sc ack clears.
    if(clock'event and clock = '1') then                
      for W in 0 to num_stores-1 loop
        
        -- if ack and req are both asserted, clear
        -- it unless asked to set it.
        if(sc_ack_flag(W) = '1' and sc_req_in(W) = '1') then
          sc_ack_clear(W) := '1';
        end if;
        
        -- set dominant!
        if(sc_ack_set(W) = '1') then
          sc_ack_flag(W) <= '1';
        elsif (sc_ack_clear(W) = '1') then
          sc_ack_flag(W) <= '0';
        end if;
      end loop;
    end if;      

    sr_ack_out <= sc_ack_set;
  end process;

  sc_ack_out <= sc_ack_flag;
  lc_ack_out <= lc_ack_flag;
  lc_data_out <= lc_data_out_sig;
  lc_tag_out <= lc_tag_out_sig;
  sc_tag_out <= sc_tag_out_sig;
  
end Default_arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_function_pack.all;
use ahir.merge_functions.all;
use ahir.mem_component_pack.all;

-- memory subsystem guarantees that accesses to the same location
-- will take place in the order of the time-stamp assigned to each
-- access (tie breaks will be random). Time-stamp is set at the
-- point of acceptance of an access request.

entity UnorderedMemorySubsystem is
  generic(name: string;
	  num_loads             : natural := 5;
          num_stores            : natural := 10;
          addr_width            : natural := 9;
          data_width            : natural := 5;
          tag_width             : natural := 7;
          -- number_of_banks       : natural := 1; (will always be 1 in this memory)
          mux_degree            : natural := 10;
          demux_degree          : natural := 10;
	  base_bank_addr_width  : natural := 8;
	  base_bank_data_width  : natural := 8);
  port(
    ------------------------------------------------------------------------------
    -- load request ports
    ------------------------------------------------------------------------------
    lr_addr_in : in std_logic_vector((num_loads*addr_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on load request.
    lr_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lr_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag for request, will be returned on completion.
    lr_tag_in : in std_logic_vector((num_loads*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- load complete ports
    ---------------------------------------------------------------------------
    lc_data_out : out std_logic_vector((num_loads*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, user should latch data_out.
    lc_req_in  : in  std_logic_vector(num_loads-1 downto 0);
    lc_ack_out : out std_logic_vector(num_loads-1 downto 0);

    -- tag of completed request.
    lc_tag_out : out std_logic_vector((num_loads*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- store request ports
    ------------------------------------------------------------------------------
    sr_addr_in : in std_logic_vector((num_stores*addr_width)-1 downto 0);
    sr_data_in : in std_logic_vector((num_stores*data_width)-1 downto 0);

    -- req/ack pair:
    -- when both are asserted, time-stamp is set on store request.
    sr_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sr_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag for request, will be returned on completion.
    sr_tag_in : in std_logic_vector((num_stores*tag_width)-1 downto 0);

    ---------------------------------------------------------------------------
    -- store complete ports
    ---------------------------------------------------------------------------
    -- req/ack pair:
    -- when both are asserted, user assumes that store is done.
    sc_req_in  : in  std_logic_vector(num_stores-1 downto 0);
    sc_ack_out : out std_logic_vector(num_stores-1 downto 0);

    -- tag of completed request.
    sc_tag_out : out std_logic_vector((num_stores*tag_width)-1 downto 0);

    ------------------------------------------------------------------------------
    -- clock, reset
    ------------------------------------------------------------------------------
    clock : in std_logic;  -- only rising edge is used to trigger activity.
    reset : in std_logic               -- active high.
    );
end entity UnorderedMemorySubsystem;


architecture struct of UnorderedMemorySubsystem is

  
  constant c_load_port_id_width : natural := Maximum(1,Ceil_Log2(num_loads));
  constant c_store_port_id_width : natural := Maximum(1,Ceil_Log2(num_stores));

  type LoadPortIdArray is array (natural range <>) of std_logic_vector(c_load_port_id_width-1 downto 0);
  type StorePortIdArray is array (natural range <>) of std_logic_vector(c_store_port_id_width-1 downto 0);
  
  function StorePortIdGen (
    constant x : natural;
    constant width : natural
    )
    return StorePortIdArray
  is
    variable ret_var : StorePortIdArray(0 to x-1);
    variable curr_value : std_logic_vector(width-1 downto 0);
  begin
    curr_value := (others => '0');
    ret_var := (others => (others => '0'));
    for I  in 0 to x-1 loop
      ret_var(I) := curr_value;
      curr_value := IncrementSLV(curr_value);
    end loop;  -- I
    return(ret_var);
  end function StorePortIdGen;

  function LoadPortIdGen (
    constant x : natural;
    constant width : natural
    )
    return LoadPortIdArray
  is
    variable ret_var : LoadPortIdArray(0 to x-1);
    variable curr_value : std_logic_vector(width-1 downto 0);
  begin
    curr_value := (others => '0');
    ret_var := (others => (others => '0'));
    for I  in 0 to x-1 loop
      ret_var(I) := curr_value;
      curr_value := IncrementSLV(curr_value);
    end loop;  -- I
    return(ret_var);
  end function LoadPortIdGen;

  constant c_load_port_id_array : LoadPortIdArray(0 to num_loads-1) := LoadPortIdGen(num_loads, c_load_port_id_width);
  signal s_load_port_id_array: LoadPortIdArray(0 to num_loads-1);
  constant c_store_port_id_array : StorePortIdArray(0 to num_stores-1) := StorePortIdGen(num_stores, c_store_port_id_width);
  signal s_store_port_id_array: StorePortIdArray(0 to num_stores-1) ;

  constant rd_mux_data_width: integer :=  (addr_width + tag_width + c_load_port_id_width );
  constant wr_mux_data_width: integer :=  (addr_width + data_width + tag_width + c_store_port_id_width);

  signal rd_mux_data_in : std_logic_vector((num_loads*rd_mux_data_width)-1 downto 0);
  signal rd_mux_data_out : std_logic_vector(rd_mux_data_width-1 downto 0);
  signal rd_mux_out_req : std_logic;
  signal rd_mux_out_ack : std_logic;

  signal wr_mux_data_in : std_logic_vector((num_stores*wr_mux_data_width)-1 downto 0);
  signal wr_mux_data_out : std_logic_vector(wr_mux_data_width-1 downto 0);
  signal wr_mux_out_req : std_logic;
  signal wr_mux_out_ack : std_logic;

  signal rd_demux_sel_in  : std_logic_vector(c_load_port_id_width-1 downto 0);
  signal rd_demux_data_in : std_logic_vector(data_width+tag_width-1 downto 0);
  signal rd_demux_data_out : std_logic_vector((num_loads*(data_width+tag_width))-1 downto 0);
  signal rd_demux_in_req, rd_demux_in_ack : std_logic;
  signal rd_demux_out_req, rd_demux_out_ack : std_logic_vector(num_loads-1 downto 0);

  signal wr_demux_sel_in : std_logic_vector(c_store_port_id_width-1 downto 0);
  signal wr_demux_data_in : std_logic_vector(tag_width-1 downto 0);
  signal wr_demux_data_out : std_logic_vector((num_stores*tag_width)-1 downto 0);
  signal wr_demux_in_req, wr_demux_in_ack : std_logic;
  signal wr_demux_out_req, wr_demux_out_ack : std_logic_vector(num_stores-1 downto 0);

  signal mem_bank_write_data     : std_logic_vector(data_width-1 downto 0);
  signal mem_bank_write_addr     : std_logic_vector(addr_width-1 downto 0);
  signal mem_bank_write_tag, mem_bank_write_tag_out : 
	std_logic_vector(tag_width+c_store_port_id_width-1 downto 0);
  signal mem_bank_write_enable   : std_logic;
  signal mem_bank_write_ack   : std_logic;
  signal mem_bank_write_result_accept : std_logic;
  signal mem_bank_write_result_ready : std_logic;
  signal mem_bank_read_data     : std_logic_vector(data_width-1 downto 0);
  signal mem_bank_read_addr     : std_logic_vector(addr_width-1 downto 0);
  signal mem_bank_read_tag,mem_bank_read_tag_out  : std_logic_vector((c_load_port_id_width+tag_width)-1 downto 0);
  signal mem_bank_read_enable   : std_logic;
  signal mem_bank_read_ack      : std_logic;
  signal mem_bank_read_result_accept: std_logic;
  signal mem_bank_read_result_ready: std_logic;

begin

   s_load_port_id_array <= c_load_port_id_array;
   s_store_port_id_array <= c_store_port_id_array;

   -- read mux data aggregation
   process(lr_addr_in, lr_tag_in)
   begin
	for I in 0 to num_loads-1 loop
		rd_mux_data_in((rd_mux_data_width*(I+1))-1 downto rd_mux_data_width*I)
			<= lr_addr_in((addr_width*(I+1))-1 downto addr_width*I) &
				lr_tag_in((tag_width*(I+1))-1 downto tag_width*I) &
				   c_load_port_id_array(I); 
	end loop;
   end process;

  
   -- read mux data aggregation
   process(sr_addr_in,sr_data_in, sr_tag_in)
   begin
	for I in 0 to num_stores-1 loop
		wr_mux_data_in((wr_mux_data_width*(I+1))-1 downto wr_mux_data_width*I)
			<= sr_addr_in((addr_width*(I+1))-1 downto addr_width*I) & 
			     sr_data_in((data_width*(I+1))-1 downto data_width*I) & 
				sr_tag_in((tag_width*(I+1))-1 downto tag_width*I) &
				 c_store_port_id_array(I); 
	end loop;
   end process;
 
   -- Readmux instantiation.
   rmux: PipelinedMux generic map(name => name & "-rmux", g_number_of_inputs => num_loads,
				g_data_width => rd_mux_data_width,
			        g_mux_degree => mux_degree,
				g_port_id_width => c_load_port_id_width)
		port map(merge_data_in => rd_mux_data_in,
			  merge_req_in => lr_req_in,
			  merge_ack_out => lr_ack_out,
			  merge_data_out => rd_mux_data_out,
			  merge_req_out => rd_mux_out_req,
			  merge_ack_in => rd_mux_out_ack,
		          clock => clock,
			  reset => reset);	

    -- connect rmux to memory bank
    mem_bank_read_addr <= rd_mux_data_out(rd_mux_data_width-1 downto (rd_mux_data_width-addr_width));
    mem_bank_read_tag <= rd_mux_data_out((rd_mux_data_width-addr_width)-1 downto 0); -- tag & port-id
    mem_bank_read_enable <= rd_mux_out_req;
    rd_mux_out_ack <= mem_bank_read_ack;
    
				
   -- Writemux instantiation.
   wmux: PipelinedMux generic map(name => name & "-wmux", g_number_of_inputs => num_stores,
				g_data_width => wr_mux_data_width,
			        g_mux_degree => mux_degree,
				g_port_id_width => c_store_port_id_width)
		port map(merge_data_in => wr_mux_data_in,
			  merge_req_in => sr_req_in,
			  merge_ack_out => sr_ack_out,
			  merge_data_out => wr_mux_data_out,
			  merge_req_out => wr_mux_out_req,
			  merge_ack_in => wr_mux_out_ack,
		          clock => clock,
			  reset => reset);	

    -- connect to memory bank.
    mem_bank_write_addr <= wr_mux_data_out(wr_mux_data_width-1 downto (wr_mux_data_width-addr_width));
    mem_bank_write_data <= wr_mux_data_out((wr_mux_data_width-addr_width)-1 downto 
	((wr_mux_data_width-addr_width)-data_width));
    mem_bank_write_tag <= wr_mux_data_out((wr_mux_data_width-(data_width+addr_width))-1 downto 0);
    mem_bank_write_enable <= wr_mux_out_req;
    wr_mux_out_ack <= mem_bank_write_ack;


    -- the memory bank..
    mbank: memory_bank generic map(name => name & "-mbank", 
				   g_addr_width => addr_width,
				   g_data_width => data_width,
				   g_write_tag_width => (tag_width + c_store_port_id_width),
				   g_read_tag_width => (tag_width + c_load_port_id_width),
				   g_time_stamp_width => 0,  -- no time-stamp.
				   g_base_bank_addr_width => base_bank_addr_width,
			           g_base_bank_data_width => base_bank_data_width)
		port map(clk => clock,
			 reset => reset,
			 write_data => mem_bank_write_data,
			 write_addr => mem_bank_write_addr,
			 write_tag => mem_bank_write_tag,
			 write_tag_out => mem_bank_write_tag_out,
			 write_enable => mem_bank_write_enable,
			 write_ack => mem_bank_write_ack,
			 write_result_ready => mem_bank_write_result_ready,
			 write_result_accept => mem_bank_write_result_accept,
			 read_data => mem_bank_read_data,
			 read_addr => mem_bank_read_addr,
			 read_tag => mem_bank_read_tag,
			 read_tag_out => mem_bank_read_tag_out,
			 read_enable => mem_bank_read_enable,
			 read_ack => mem_bank_read_ack,
			 read_result_ready => mem_bank_read_result_ready,
			 read_result_accept => mem_bank_read_result_accept);
			

    -- memory bank to read-demux
    rd_demux_sel_in  <= mem_bank_read_tag_out(c_load_port_id_width-1 downto 0);
    rd_demux_data_in <= mem_bank_read_data & mem_bank_read_tag_out((tag_width+c_load_port_id_width)-1 downto c_load_port_id_width);
    rd_demux_in_req <= mem_bank_read_result_ready;
    mem_bank_read_result_accept <= rd_demux_in_ack;
 
    rd_demux: PipelinedDemux generic map (name => name & "-rd_demux",
					g_data_width => data_width+tag_width,
				       g_destination_id_width => c_load_port_id_width,
				       g_number_of_outputs => num_loads)
		port map(data_in => rd_demux_data_in,
			 sel_in => rd_demux_sel_in,
			 req_in => rd_demux_in_req,
			 ack_out => rd_demux_in_ack,
			 data_out => rd_demux_data_out,
			 req_out => rd_demux_out_req,
			 ack_in => rd_demux_out_ack,
			 clk => clock,
			 reset => reset);

    process(rd_demux_data_out)
    begin
       for I in 0 to num_loads-1 loop
	 lc_data_out(((I+1)*data_width)-1 downto I*data_width) 
		<= rd_demux_data_out(((I+1)*(data_width+tag_width))-1 downto (I*(data_width+tag_width))+tag_width);
	 lc_tag_out(((I+1)*tag_width)-1 downto I*tag_width) 
		<= rd_demux_data_out((I*(data_width+tag_width))+tag_width-1 downto (I*(data_width+tag_width)));
       end loop;
    end process;

    rd_demux_out_ack <= lc_req_in;
    lc_ack_out <= rd_demux_out_req;
					 
    -- memory bank to write-demux
    wr_demux_sel_in <= mem_bank_write_tag_out(c_store_port_id_width-1 downto 0);
    wr_demux_data_in <= mem_bank_write_tag_out(tag_width+c_store_port_id_width-1 downto c_store_port_id_width);
    wr_demux_in_req <= mem_bank_write_result_ready;
    mem_bank_write_result_accept <= wr_demux_in_ack;
    
    wr_demux: PipelinedDemux generic map (name => name & "-wr_demux",
					g_data_width => tag_width,
				       g_destination_id_width => c_store_port_id_width,
				       g_number_of_outputs => num_stores)
		port map(data_in => wr_demux_data_in,
			 sel_in => wr_demux_sel_in,
			 req_in => wr_demux_in_req,
			 ack_out => wr_demux_in_ack,
			 data_out => wr_demux_data_out,
			 req_out => wr_demux_out_req,
			 ack_in => wr_demux_out_ack,
			 clk => clock,
			 reset => reset);

    sc_tag_out <= wr_demux_data_out;
    wr_demux_out_ack <= sc_req_in;
    sc_ack_out <= wr_demux_out_req;

end struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- author: Madhav Desai
--
-- limit the number of pending requests
-- to at most num_slots.
--
--  That is, forward req -> regulated-req
--  only if the numer of pending req's which
--  have not been acked is less than num_slots.
--
library ieee;
use ieee.std_logic_1164.all;


-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;
entity access_regulator_base is
  generic (name : string;  num_slots: integer := 1);
  port (
    -- the req-ack pair being regulated.
    req   : in Boolean;
    ack   : out Boolean;
    -- the regulated versions of req/ack
    regulated_req : out Boolean;
    regulated_ack : in Boolean;
    -- transitions on the next two will
    -- open up a slot.
    release_req   : in Boolean;
    release_ack   : in Boolean; -- this is superfluous..
    clk   : in  std_logic;
    reset : in  std_logic);

end access_regulator_base;

architecture default_arch of access_regulator_base is
  
   signal req_place_preds, req_place_succs : BooleanArray(0 downto 0);
   signal req_place_token : Boolean;

   signal release_req_place_preds, release_ack_place_preds: BooleanArray(0 downto 0);
   signal release_req_place_succs, release_ack_place_succs: BooleanArray(0 downto 0);
   signal release_req_place_token, release_ack_place_token: boolean;
   
   signal regulated_req_join_preds: BooleanArray(2 downto 0);
   signal regulated_req_token: Boolean; 
  
   signal regulated_req_join: boolean;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- default_arch

   req_place_preds(0) <= req;
   reqPlace: place_with_bypass 
	generic map(capacity => 1, marking => 0, name => name & ":req_place:")
	port map(preds => req_place_preds, 
			succs => req_place_succs, 
			token => req_place_token,
				clk => clk, reset => reset);


   -- the next two places manage the slots
   -- note that the capacity must be num_slots+1, because
   -- a release requests may arrive earlier than the 
   -- unregulated request.  However at most one release-request
   -- can arrive before the first request (because of the way the
   -- CP is constructed).
   release_req_place_preds(0) <= release_req;
   releaseReqPlace: place 
	generic map(capacity => num_slots+1, marking => num_slots, name => name & ":release_req_place:")
	port map(preds => release_req_place_preds, 
			succs => release_req_place_succs, 
			token => release_req_place_token,
			clk => clk, reset => reset);


   -- the join fires when all places have tokens. 
   regulated_req_join <= release_req_place_token and req_place_token;
   release_req_place_succs(0) <= regulated_req_join;
   req_place_succs(0) <= regulated_req_join;


   -- the req that goes out.
   -- the req goes out only if a token is present in the req-place, the release-req-place
   -- and the release-ack place.
   regulated_req <= regulated_req_join;

   -- ack from RHS is forwarded to the left.
   ack <= regulated_ack;
   
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- author: Madhav Desai.

library ahir;
use ahir.Types.all;
use ahir.Utilities.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;


entity access_regulator is
  generic (name: string; num_reqs : integer := 1; num_slots: integer := 1);
  port (
    -- the req-ack pair being regulated.
    req   : in BooleanArray(num_reqs-1 downto 0);
    ack   : out BooleanArray(num_reqs-1 downto 0);
    -- the regulated versions of req/ack
    regulated_req : out BooleanArray(num_reqs-1 downto 0);
    regulated_ack : in BooleanArray(num_reqs-1 downto 0);
    -- transitions on the next two will
    -- open up a slot.
    release_req   : in BooleanArray(num_reqs-1 downto 0);
    release_ack   : in BooleanArray(num_reqs-1 downto 0);
    clk   : in  std_logic;
    reset : in  std_logic);

end access_regulator;

architecture default_arch of access_regulator is


begin  -- default_arch
   gen: for I in 0 to num_reqs-1 generate
	aR: access_regulator_base generic map(name => name & "(" & Convert_To_String(I) & ")", num_slots => num_slots)
		port map(req => req(I),
			 ack => ack(I),
			 regulated_req => regulated_req(I),
			 regulated_ack => regulated_ack(I),
			 release_req => release_req(I),
			 release_ack => release_ack(I),
			 clk => clk, 
			 reset => reset);
   end generate gen;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- on reset, trigger an AHIR module, and keep
-- retriggering it..
entity auto_run is
  generic (
    use_delay : boolean := true);
  port (clk   : in  std_logic;
    	reset : in  std_logic;
	start_req: out std_logic;
        start_ack: in std_logic;
        fin_req: out std_logic;
        fin_ack: in std_logic);
end auto_run;

architecture default_arch of auto_run is

begin  

  process(clk)
  begin
    if(clk'event and clk = '1') then
	if(reset = '1') then
		start_req <= '0';
 		fin_req <= '0';
	else
		start_req <= '1';
		fin_req <= '1';
	end if;
    end if;
  end process;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- conditional-fork.
--    forward in-transition to out-transitions if triggers are enabled.
-- written by Madhav P. Desai, December 2015.
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.Utilities.all;

-- for a transition on in-transition, produce a transition on an out-transitions 
-- if the trigger is enabled (disable all triggers when the out-transition is fired).
entity conditional_fork is
       generic (place_capacity: integer := 1; 
			ntriggers: integer; name : string);
       port (triggers: in BooleanArray(0 to ntriggers-1);
			in_transition: in Boolean;
			out_transitions: out BooleanArray(0 to ntriggers-1);
			clk: in std_logic; reset: in std_logic);
end entity conditional_fork;

architecture Basic of conditional_fork is
    signal trig_places, trig_clears: BooleanArray(0 to ntriggers-1);
    signal in_trans_place, in_trans_clear: Boolean;
begin
    TrigPlaces: for I in 0 to (ntriggers-1) generate
	placeBlock: block
	  signal place_pred, place_succ: BooleanArray(0 downto 0);
        begin
	  place_pred(0) <= triggers(I);
	  place_succ(0) <= trig_clears(I);

          -- a bypass place: in order to speed up loop turnaround times.
	  pI: place_with_bypass generic map(capacity => place_capacity, marking => 0,
		     name => name & ":trigplaces:" & Convert_To_String(I))
		  port map(preds => place_pred,succs =>place_succ,token => trig_places(I),clk => clk, reset => reset);
        end block;
    end generate TrigPlaces;

    inTransPlaceBlock: block
      signal place_pred, place_succ: BooleanArray(0 downto 0);
    begin
      place_pred(0) <= in_transition;
      place_succ(0) <= in_trans_clear;

      -- a bypass place: in order to speed up loop turnaround times.
      pI: place_with_bypass generic map(capacity => place_capacity, marking => 0,
		     name => name & ":inTransPlace:")
		  port map(preds => place_pred, succs => place_succ,token => in_trans_place, clk => clk, reset => reset);
    end block;

    cGen: for I in 0 to ntriggers-1 generate
	trig_clears(I) <= in_trans_place and trig_places(I);
	out_transitions(I) <= trig_clears(I);
    end generate cGen;
  
     -- clear in-transition when any of the trigs are cleared.
     in_trans_clear <= OrReduce(trig_clears);

end Basic;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
entity control_delay_element is
  generic (name: string; delay_value: integer := 0);
  port (
    req   : in Boolean;
    ack   : out Boolean;
    clk   : in  std_logic;
    reset : in  std_logic);

end control_delay_element;

architecture default_arch of control_delay_element is
  
-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- default_arch

  ZeroDelay: if (delay_value <= 0) generate
    ack <= req;
  end generate ZeroDelay;

  UnitDelay: if (delay_value = 1) generate

	process(clk)
        begin
		if(clk'event and clk = '1') then 
			if(reset = '1') then
				ack <= false;
			else	
				ack <= req;
			end if;
		end if;
	end process;

  end generate UnitDelay;


  DelayGTOne: if (delay_value > 1) generate

   ShiftReg: block
	signal sr_state: BooleanArray(0 to delay_value-1);
   begin
 	process(clk)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				sr_state <= (others => false);
			else
				sr_state(0) <= req;
				for I in 1 to delay_value-1 loop
					sr_state(I) <= sr_state(I-1);
				end loop;
			end if;
		end if;
	end process;
	ack <= sr_state(delay_value-1);
   end block;
  end generate DelayGTOne;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;

use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.utilities.all;

entity generic_join is
  generic(number_of_predecessors: integer; name: string; place_capacities: IntegerArray; place_markings: IntegerArray; place_delays: IntegerArray);
  port ( preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end generic_join;

architecture default_arch of generic_join is
  signal symbol_out_sig : BooleanArray(0 downto 0);
  signal place_sigs: BooleanArray(1 to preds'length);
  constant pmarkings : IntegerArray(1 to preds'length) := place_markings;
  constant pcapacities: IntegerArray(1 to preds'length) := place_capacities;
  constant pdelays: IntegerArray(1 to preds'length) := place_delays;
  alias ppreds : BooleanArray(1 to preds'length) is preds;
begin  -- default_arch

  assert ((preds'length = place_capacities'length) and (place_capacities'length = place_delays'length)
		and (place_delays'length = place_markings'length) )
	report "Mismatch in lengths of marking/capacity arrays." severity failure;
  
  placegen: for I in 1 to number_of_predecessors generate
    placeBlock: block
	signal place_pred: BooleanArray(0 downto 0);
    begin
      dly: control_delay_element generic map(name => name & "-placegen-dly-" & Convert_To_String(I), delay_value => pdelays(I))
                   port map(req => ppreds(I), ack => place_pred(0), clk => clk, reset => reset);
      pI: place_with_bypass
        generic map(capacity => pcapacities(I),
                    marking => pmarkings(I),
                    name => name & "-placegen-pI-" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
    end block;
  end generate placegen;

  -- The transition is enabled only when all preds are true.
  symbol_out_sig(0) <= AndReduce(place_sigs);
  symbol_out <= symbol_out_sig(0);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;

entity join2 is
  generic(bypass : boolean := true; name : string);
  port ( pred0, pred1      : in   Boolean;
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end join2;

architecture default_arch of join2 is
  signal preds: BooleanArray(1 downto 0);
begin  -- default_arch

  preds <= pred0 & pred1;
  baseJoin : join
    generic map(number_of_predecessors => 2, bypass => bypass, name => name & ":base")
    port map (preds => preds,
              symbol_out => symbol_out,
              clk => clk,
              reset => reset);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;

entity join3 is
  generic(bypass : boolean := true; name: string);
  port ( pred0, pred1, pred2      : in   Boolean;
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end join3;

architecture default_arch of join3 is
  signal preds: BooleanArray(2 downto 0);
begin  -- default_arch

  preds <= pred0 & pred1 & pred2;
  baseJoin : join
    generic map(number_of_predecessors => 3, bypass => bypass, name => name & ":base")
    port map (preds => preds,
              symbol_out => symbol_out,
              clk => clk,
              reset => reset);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.utilities.all;

entity join is
  generic (number_of_predecessors: integer; place_capacity : integer := 1;bypass: boolean := true; name : string );
  port ( preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end join;

architecture default_arch of join is
  signal symbol_out_sig : BooleanArray(0 downto 0);
  signal place_sigs: BooleanArray(preds'range);
  constant H: integer := preds'high;
  constant L: integer := preds'low;

begin  -- default_arch
  
  placegen: for I in H downto L generate
    placeBlock: block
	signal place_pred: BooleanArray(0 downto 0);
    begin
	place_pred(0) <= preds(I);

      bypassgen: if bypass generate
	pI: place_with_bypass
		generic map(capacity => place_capacity, 
				marking => 0,
				name => name & ":" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
      end generate bypassgen;

      nobypassgen: if (not bypass) generate
	pI: place
		generic map(capacity => place_capacity, 
				marking => 0,
				name => name & ":" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
      end generate nobypassgen;

    end block;
  end generate placegen;
  -- The transition is enabled only when all preds are true.
  
  symbol_out_sig(0) <= AndReduce(place_sigs);
  symbol_out <= symbol_out_sig(0);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.utilities.all;

entity join_with_input is
  generic (number_of_predecessors: integer; place_capacity : integer := 1; bypass : boolean := true; name : string);
  port ( preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
    	symbol_in  : in   boolean;
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end join_with_input;

architecture default_arch of join_with_input is
  signal symbol_out_sig : BooleanArray(0 downto 0);
  signal place_sigs: BooleanArray(preds'range);
  signal inp_place_sig: Boolean;
  constant H: integer := number_of_predecessors-1;
  constant L: integer := 0;
begin  -- default_arch
  
  Byp: if bypass generate 
    placegen: for I in H downto L generate
      placeBlock: block
	  signal place_pred: BooleanArray(0 downto 0);
      begin
	  place_pred(0) <= preds(I);
	  pI: place_with_bypass generic map(capacity => place_capacity, marking => 0,
				   name => name & ":" & Convert_To_String(I) )
		  port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
      end block;
    end generate placegen;
    
    inplaceBlock: block
	  signal place_pred: BooleanArray(0 downto 0);
    begin
	  place_pred(0) <= symbol_in;
	  pI: place_with_bypass generic map(capacity => place_capacity, marking => 0,
				   name => name & ":inputplace")
		  port map(place_pred,symbol_out_sig,inp_place_sig,clk,reset);
    end block;
  end generate Byp;

  NoByp: if (not bypass) generate 
    placegen: for I in H downto L generate
      placeBlock: block
	  signal place_pred: BooleanArray(0 downto 0);
      begin
	  place_pred(0) <= preds(I);
	  pI: place generic map(capacity => place_capacity, marking => 0,
				   name => name & ":" & Convert_To_String(I) )
		  port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
      end block;
    end generate placegen;
    
    inplaceBlock: block
	  signal place_pred: BooleanArray(0 downto 0);
    begin
	  -- note: input transitions are always bypassed, because they
	  --       always come with a delay (no need to incur an additional delay for them).
	  place_pred(0) <= symbol_in;
	  pI: place_with_bypass generic map(capacity => place_capacity, marking => 0,
				   name => name & ":inputplace")
		  port map(place_pred,symbol_out_sig,inp_place_sig,clk,reset);
    end block;
  end generate NoByp;


  -- The transition is enabled only when all preds are true.
  symbol_out_sig(0) <= inp_place_sig and AndReduce(place_sigs);
  symbol_out <= symbol_out_sig(0);
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.BaseComponents.all;
-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##


-- on reset, trigger an AHIR module, and keep
-- retriggering it..
-- TODO: add a single cycle delay in lreq -> preq
-- path and also in the pack -> lack path in order
-- to control the clock period...
entity level_to_pulse is
  generic (name: string; forward_delay: integer; backward_delay: integer);
  port (clk   : in  std_logic;
    	reset : in  std_logic;
        lreq: in std_logic;
        lack: out std_logic;
        preq: out boolean;
        pack: in boolean);
end level_to_pulse;

architecture default_arch of level_to_pulse is
  type L2PState is (idle,waiting);
  signal l2p_state : L2PState;
  signal pack_sig, preq_sig: boolean;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

  process(clk,reset,lreq, pack_sig, l2p_state)
    variable nstate : L2PState;
    variable lack_v : std_logic;
    variable preq_v : boolean;
    
  begin
    lack_v := '0';
    preq_v := false;
    nstate := l2p_state;
    if(l2p_state = idle) then
      if(lreq ='1') then
        preq_v := true;
        if(pack_sig) then
          lack_v := '1';
        else
          nstate := waiting;
        end if;
      end if;
    else
      if(pack_sig) then
        lack_v := '1';
        nstate := idle;
      end if;
    end if;

    lack     <= lack_v;
    preq_sig <= preq_v;
    
    if(reset = '1') then
      nstate := idle;
    end if;

    if(clk'event and clk = '1') then
      l2p_state <= nstate;
    end if;
    
  end process;

  fDelay: control_delay_element generic map(name => name & "-fDelay", delay_value => forward_delay)
	port map(req => preq_sig, ack => preq, clk => clk, reset => reset);

  bDelay: control_delay_element generic map(name => name & "-bDelay", delay_value => backward_delay)
	port map(req => pack, ack => pack_sig, clk => clk, reset => reset);

  
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- loop-terminator element for use in pipelined loops.
-- written by Madhav P. Desai, December 2012.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.utilities.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity loop_terminator is
  
  generic (name: string; max_iterations_in_flight : integer := 4);
  port(loop_body_exit: in boolean;
       loop_continue: in boolean;
       loop_terminate: in boolean;
       loop_back: out boolean;
       loop_exit: out boolean;
       clk: in std_logic;
       reset: in std_logic);

end loop_terminator;

--
-- Let M = max iterations in flight.
--
-- initialize the counter (at reset) to M-1.
--
-- Anytime you see loop-body-exit, increment the
-- counter
--
-- if lc has arrived, and if the counter is > 0,
-- then emit loop-back, and decrement the counter.
--
-- if lt has arrived, wait until the counter reaches M
-- and then emit loop-exit, resetting the counter to M-1.
--
architecture Behave of loop_terminator is

  type FSMState is (idle, pending_continue, pending_exit);

  signal fsm_state : FSMState;
  signal available_iterations : unsigned ((Ceil_Log2(max_iterations_in_flight+1) - 1) downto 0);

  signal lc_place_preds, lc_place_succs : BooleanArray(0 downto 0);
  signal clear_lc_place, lc_place_token : boolean;

  signal lt_place_preds, lt_place_succs : BooleanArray(0 downto 0);
  signal clear_lt_place, lt_place_token: boolean;

  signal lbe_place_preds, lbe_place_succs : BooleanArray(0 downto 0);
  signal clear_lbe_place, lbe_place_token: boolean;  
  
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  -- places to remember loop-continue, loop-terminate, loop-body-exit

  -- critical place: make it a bypass place in order to
  -- speed up loop turnaround times.  The clock period
  -- will not be an issue since the branch ack is 
  -- registered.
  lc_place : place_with_bypass generic map (
    capacity => 1,
    marking  => 0,
    name => "loop_terminator:lc_place")
    port map (
      preds => lc_place_preds,
      succs => lc_place_succs,
      token => lc_place_token,
      clk   => clk,
      reset => reset);
  lc_place_preds(0) <= loop_continue;
  lc_place_succs(0) <= clear_lc_place;

  lt_place : place generic map (
    capacity => 1,
    marking  => 0,
    name => "loop_terminator:lt_place")
    port map (
      preds => lt_place_preds,
      succs => lt_place_succs,
      token => lt_place_token,
      clk   => clk,
      reset => reset);
  lt_place_preds(0) <= loop_terminate;
  lt_place_succs(0) <= clear_lt_place;


  lbe_place : place generic map (
    capacity => 1,
    marking  => 0,
    name => "loop_terminator:lbe_place")
    port map (
      preds => lbe_place_preds,
      succs => lbe_place_succs,
      token => lbe_place_token,
      clk   => clk,
      reset => reset);
  lbe_place_preds(0) <= loop_body_exit;
  lbe_place_succs(0) <= clear_lbe_place;
  
  -- state machine:
  --   inputs
  --   lc_place_token, lt_place_token, lbe_place_token, available_iterations.
  --   outputs
  --   clear_lc_place, clear_lt_place, clear_lbe_place, loop_back,
  --   loop_exit, available_iterations.
  --   
  process(clk, reset,lc_place_token,lt_place_token,lbe_place_token,available_iterations)
    variable next_available_iterations : 
		unsigned(available_iterations'high downto available_iterations'low);
    variable incr,decr,rst : boolean;
  begin
    -- all outputs are deasserted by default.
    loop_back <= false;
    loop_exit <= false;
    clear_lc_place <= false;
    clear_lt_place <= false;
    clear_lbe_place <= false;
    
    -- incr, decr, rst are used to manage count.
    incr := false;
    decr := false;
    if(reset = '1') then
      rst := true;
    else
      rst := false;
    end if;

    -- lbe always increments counter.
    if(lbe_place_token) then
      incr := true;
      clear_lbe_place <= true;
    end if;

    -- loop-continue? emit loop-back if count > 0..
    -- and decrement count, clear lc place.      
    if(lc_place_token and (available_iterations > 0)) then
      decr := true;
      loop_back <= true;
      clear_lc_place <= true;
    end if;

    -- loop-terminate? check if count will reach M, and emit loop_exit, reset counter.
    if(lt_place_token and 
		((available_iterations = max_iterations_in_flight) or 
			-- dont waste a cycle... loop-body-exit should be applied
			-- right away
			(incr and (not decr) and 
				(available_iterations = (max_iterations_in_flight-1))))) then
      rst := true;
      loop_exit <= true;
      clear_lt_place <= true;          
    end if;

    -- manage count.
    if(rst) then
       next_available_iterations := To_Unsigned(max_iterations_in_flight - 1, available_iterations'length);
    elsif (incr and (not decr)) then
       next_available_iterations := (available_iterations + 1);
    elsif (decr and (not incr)) then
       next_available_iterations := (available_iterations - 1);
    else
       next_available_iterations := available_iterations;
    end if;

    if(clk'event and clk = '1') then
	available_iterations <= next_available_iterations;
    end if;

  end process;

  assert (available_iterations > 0)  report "available_iterations = 0 in " & name  severity note;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.utilities.all;

entity marked_join is
  generic(number_of_predecessors: integer; number_of_marked_predecessors: integer;
		place_capacity : integer := 1; bypass : boolean := true; name : string; marked_predecessor_bypass: BooleanArray);
  port ( preds      : in   BooleanArray(number_of_predecessors-1 downto 0);
         marked_preds : in BooleanArray(number_of_marked_predecessors-1 downto 0);
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end marked_join;

architecture default_arch of marked_join is
  signal symbol_out_sig : BooleanArray(0 downto 0);
  signal place_sigs: BooleanArray(preds'range);
  signal mplace_sigs: BooleanArray(marked_preds'range);  
  constant H: integer := preds'high;
  constant L: integer := preds'low;

  constant MH: integer := marked_preds'high;
  constant ML: integer := marked_preds'low;  

  constant mbypass: BooleanArray(MH downto ML) := marked_predecessor_bypass;

begin  -- default_arch
  
  placegen: for I in H downto L generate
    placeBlock: block
	signal place_pred: BooleanArray(0 downto 0);
    begin
	place_pred(0) <= preds(I);
      bypassgen: if (bypass) generate
	pI: place_with_bypass
		generic map(capacity => place_capacity, 
				marking => 0,
				name => name & ":(bypass):" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
      end generate bypassgen;

      nobypassgen: if (not bypass) generate
	pI: place
		generic map(capacity => place_capacity, 
				marking => 0,
				name => name & ":(no-bypass):" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,place_sigs(I),clk,reset);
      end generate nobypassgen;
    end block;
  end generate placegen;

  -- the marked places
  mplacegen: for I in MH downto ML generate
    mplaceBlock: block
	signal place_pred: BooleanArray(0 downto 0);
    begin
	place_pred(0) <= marked_preds(I);
	bypassGen: if mbypass(I)  generate
	   mpI: place_with_bypass generic map(capacity => place_capacity, marking => 1, 
				 name => name & ":marked(bypass):" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,mplace_sigs(I),clk,reset);
	end generate bypassGen;
	NobypassGen: if (not mbypass(I))  generate
	  mpI: place generic map(capacity => place_capacity, marking => 1, 
				 name => name & ":marked(no-bypass):" & Convert_To_String(I) )
		port map(place_pred,symbol_out_sig,mplace_sigs(I),clk,reset);
	end generate NobypassGen;

    end block;
  end generate mplacegen;
  
  -- The transition is enabled only when all preds are true.
  symbol_out_sig(0) <= AndReduce(place_sigs) and AndReduce(mplace_sigs);
  symbol_out <= symbol_out_sig(0);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;

entity out_transition is
  
  port (preds      : in   BooleanArray;
        symbol_out : out  boolean);

end out_transition;

architecture default_arch of out_transition is
begin  -- default_arch

  -- The transition is enabled only when all preds are true.
  symbol_out <= AndReduce(preds);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- phi-sequencer.. improved version
--  src-expressions are triggered only when needed
--  (as opposed to the old phi which was clumsy).
-- written by Madhav P. Desai, December 2015.
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.Utilities.all;
use ahir.GlobalConstants.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity phi_sequencer_v2  is
  generic (place_capacity : integer; 
	   ntriggers : integer; 
	   name : string);
  port (
  	triggers : in BooleanArray(0 to ntriggers-1); 	    -- there are nreq triggers.
  	src_sample_starts : out BooleanArray(0 to ntriggers-1);   -- sample starts for sources.
	src_sample_completes: in BooleanArray(0 to ntriggers-1);  -- sample completes from sources.
  	src_update_starts : out BooleanArray(0 to ntriggers-1);   -- update starts for sources.
	src_update_completes: in BooleanArray(0 to ntriggers-1);  -- update completes from sources.
  	phi_sample_req  : in Boolean;			   	  -- incoming sample-req to phi.
	phi_sample_ack  : out Boolean;				  -- outgoing sample-ack from phi.
  	phi_update_req  : in Boolean;			   	  -- incoming update-req to phi.
	phi_update_ack  : out Boolean;				  -- outgoing update-ack from phi.
  	phi_mux_select_reqs    : out BooleanArray(0 to ntriggers-1);	  -- phi-select mux select reqs.
	phi_mux_ack: in Boolean;				  -- ack from mux signifying select complete.
  	clk, reset: in std_logic);
end phi_sequencer_v2;


--
-- on reset, wait for a transition on any of the in_places.
-- the corresponding req is asserted..  A token in the
-- enable places is needed to allow firing of the reqs.
--
architecture Behave of phi_sequencer_v2 is
  signal trigger_tokens, trigger_clears : BooleanArray(0 to ntriggers-1);
  signal sample_wait_tokens, sample_wait_clears : BooleanArray(0 to ntriggers-1);
  signal src_update_start_tokens, src_update_start_clears : BooleanArray(0 to ntriggers-1);
  signal src_update_wait_tokens, src_update_wait_clears : BooleanArray(0 to ntriggers-1);
  signal src_sample_start_sigs : BooleanArray(0 to ntriggers-1);   -- sample starts for sources.
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  src_sample_starts <= src_sample_start_sigs;

  -- fatal: multiple triggers should never be active.
  ErrorFlag: if global_debug_flag generate
    process(clk, reset)
        variable found_flag : Boolean := false;
    begin
       found_flag := false;
       if(clk'event and clk = '1') then
         if(reset = '0') then
	   for I in 0 to ntriggers-1 loop
             if(triggers(I)) then
		if(found_flag) then
		   assert false report "Multiple triggers to phi " & name & " are active. "
				severity error;
		else
		   found_flag := true;
                end if;
             end if;
          end loop;
         end if;
       end if;
    end process;
  end generate ErrorFlag;
 
  --
  -- the sample/update pairs are totally independent.
  -- If the phi-sequencer drives an operator which does
  -- not couple the sample-req/ack pair with the
  -- update req/ack pair (as can happen if the operation
  -- is guarded, for example), then we need to introduce an additional
  -- external dependency in the control-path...
  --
  trigForkSample: conditional_fork
		generic map (place_capacity => place_capacity,
				ntriggers => ntriggers,
					name => name & ":trigFork")
		port map (triggers => triggers,
				in_transition => phi_sample_req,
					out_transitions => src_sample_start_sigs, 
						clk => clk, reset => reset);
  trigForkUpdate: conditional_fork
		generic map (place_capacity => place_capacity,
				ntriggers => ntriggers,
					name => name & ":trigFork")
		port map (triggers => triggers,
				in_transition => phi_update_req,
					out_transitions => src_update_starts, 
						clk => clk, reset => reset);
					
					

  -- mux-selects triggered by src-update completes.
  phi_mux_select_reqs <= src_update_completes;

  -- phi-sample-ack is reduced or src-sample-completes.
  phi_sample_ack <= OrReduce(src_sample_completes);

  -- phi-mux-ack goes back as phi_update_ack.
  phi_update_ack <= phi_mux_ack; 

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- phi-sequencer..
-- written by Madhav P. Desai, December 2012.
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##


entity phi_sequencer  is
  generic (place_capacity : integer; nreqs : integer; nenables : integer; name : string);
  port (
  selects : in BooleanArray(0 to nreqs-1); -- there are nreq triggers.
  reqs : out BooleanArray(0 to nreqs-1);   -- generated reqs for the phis. one for each trigger.
  ack  : in Boolean;			   -- incoming sample-ack from phi.
  enables  : in BooleanArray(0 to nenables-1);  -- enables (all have to be asserted)
  done : out Boolean;
  clk, reset: in std_logic);
end phi_sequencer;


--
-- on reset, wait for a transition on any of the in_places.
-- the corresponding req is asserted..  A token in the
-- enable places is needed to allow firing of the reqs.
--
architecture Behave of phi_sequencer is
  signal select_token, select_clear : BooleanArray(0 to nreqs-1);
  signal enable_token, enable_clear : BooleanArray(0 to nenables-1);

  signal enabled, ack_token, ack_clear, req_being_fired: Boolean;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  -- instantiate unmarked places for the in_places.
  InPlaces: for I in 0 to nreqs-1 generate
    placeBlock: block
	signal place_pred, place_succ: BooleanArray(0 downto 0);
    begin
	place_pred(0) <= selects(I);
	place_succ(0) <= select_clear(I);

        -- a bypass place: in order to speed up loop turnaround times.
	pI: place_with_bypass generic map(capacity => place_capacity, marking => 0,
		   name => name & ":select:" & Convert_To_String(I))
		port map(place_pred,place_succ,select_token(I),clk,reset);
    end block;
  end generate InPlaces;

  -- place for enables: places are unmarked.. initial state
  -- should be consistently generated by the instantiator.
  EnablePlaces: for J in 0 to nenables-1 generate
    rnb_block: block
      signal place_pred, place_succ: BooleanArray(0 downto 0);    
    begin
      place_pred(0) <= enables(J);
      place_succ(0) <= enable_clear(J);
      pRnb: place_with_bypass generic map(capacity => place_capacity, marking => 0,
		  name => name & ":enable:" & Convert_To_String(J))
        port map(place_pred,place_succ,enable_token(J),clk,reset);    
    end block;
  end generate EnablePlaces;  
    
 
  -- sequencer is enabled by this sig.
  enabled <= AndReduce(enable_token) and ack_token;

  -- a marker to indicate that a req is being fired.
  req_being_fired <= OrReduce(select_token) and enabled;

  -- outgoing reqs can fire only when the sequencer is enabled.
  reqs <= select_token when enabled else (others => false);

  -- clear the selects and reenables when the req is being fired.
  select_clear <= select_token when req_being_fired else (others => false);
  enable_clear <= (others => true) when req_being_fired else (others => false);

  -- ack should be received to reenable the sequencer.
  -- this place is initially marked (it is internal
  -- to the sequencer).
  ack_block: block
      signal place_pred: BooleanArray(0 downto 0);    
      signal place_succ: BooleanArray(0 downto 0);    
  begin
      place_pred(0) <= ack;
      place_succ(0) <= ack_clear;
      pack: place generic map(capacity => place_capacity, marking => 1,
	  	 name => name & ":ack")
        port map(place_pred,place_succ,ack_token,clk,reset);    
  end block;

  -- clear the ack place when req is fired.
  ack_clear <= req_being_fired;

  -- outgoing exit.. is the incoming ack..
  done <= ack;

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.subprograms.all;
use ahir.BaseComponents.all;

entity pipeline_interlock is
  port (trigger: in boolean;
        enable : in boolean;
    	symbol_out : out  boolean;
	clk: in std_logic;
	reset: in std_logic);
end pipeline_interlock;

architecture default_arch of pipeline_interlock is
  signal symbol_out_sig : BooleanArray(0 downto 0);
  signal enable_place_pred : BooleanArray(0 downto 0);
  signal enable_place : Boolean;
  signal trigger_place_pred : BooleanArray(0 downto 0);
  signal trigger_place : Boolean;
  

begin  -- default_arch
  

  trigger_place_pred(0) <= trigger;
  pTrig: place generic map(name => "pipeline-interlock-trigger", capacity => 1, marking => 0)
    port map(trigger_place_pred, symbol_out_sig,trigger_place,clk,reset);

  enable_place_pred(0) <= enable;
  pEnable: place generic map(name => "pipeline-interlock-enable", capacity => 1, marking => 1)
    port map(enable_place_pred, symbol_out_sig,enable_place,clk,reset);
  
  symbol_out_sig(0) <= enable_place and trigger_place;
  symbol_out <= symbol_out_sig(0);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity place is

  generic (
    capacity: integer := 1;
    marking : integer := 0;
    name   : string
    );
  port (
    preds : in  BooleanArray;
    succs : in  BooleanArray;
    token : out boolean;
    clk   : in  std_logic;
    reset : in  std_logic);

end place;

architecture default_arch of place is

  signal incoming_token : boolean;      -- true if a pred fires
  signal backward_reset : boolean;      -- true if a succ fires
  signal token_sig      : boolean;  -- asynchronously computed value of the token
  signal token_latch    : unsigned (LogWidth(capacity)-1 downto 0);
  
  constant debug_flag : boolean := global_debug_flag;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch

  assert capacity > 0 report "in place " & name & ": place must have capacity > 0." severity error;
  assert marking <= capacity report "in place " & name & ": initial marking must be less than place capacity." severity error;


  -- At most one of the preds can send a pulse.
  -- We detect it with an OR over all inputs
  incoming_token <= OrReduce(preds);

  -- At most one of the succs can send a pulse.
  -- We detect it with an OR over all inputs
  backward_reset <= OrReduce(succs);

  latch_token : process (clk, reset, token_latch, backward_reset, incoming_token)
    variable next_token_latch_var: unsigned (token_latch'high downto token_latch'low);
  begin

    next_token_latch_var := token_latch;
    if (backward_reset and (not incoming_token)) then
	if(token_latch> 0) then
            next_token_latch_var := (token_latch - 1);
        end if;
    elsif (incoming_token and (not backward_reset)) then
	if(token_latch < capacity) then
            next_token_latch_var := (token_latch + 1);
        end if;
    end if;
    
    if clk'event and clk = '1' then  -- rising clock edge
      if reset = '1' then            -- synchronous reset (active high)
        token_latch <= To_Unsigned(marking,token_latch'length);
      else
        token_latch <= next_token_latch_var;
  
        if(debug_flag) then
           if (backward_reset and (not incoming_token)) then
              assert token_latch > 0 report "in place " & name &  ": number of tokens cannot become negative!" severity error;
              assert false report "in place " & name & ": token count decremented from " & Convert_To_String(To_Integer(token_latch)) 
	severity note;
  	   elsif (incoming_token and (not backward_reset)) then
          	assert token_latch < capacity report "in place " & name & " number of tokens "
			 	& Convert_To_String(To_Integer(token_latch)+1) & " cannot exceed capacity " 
			 	& Convert_To_String(capacity) severity error;
          	assert false report "in place " & name & " token count incremented from " & Convert_To_String(To_Integer(token_latch))
		 	severity note;
       	    end if;
        end if; -- if debug_flag
      end if; -- if reset
    end if; -- if clk'event
  end process latch_token;

  token <= true when (token_latch > 0) else false;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity place_with_bypass is

  generic (
    capacity: integer := 1;
    marking : integer := 0;
    name   : string
    );
  port (
    preds : in  BooleanArray;
    succs : in  BooleanArray;
    token : out boolean;
    clk   : in  std_logic;
    reset : in  std_logic);

end place_with_bypass;

architecture default_arch of place_with_bypass is

  signal incoming_token : boolean;      -- true if a pred fires
  signal backward_reset : boolean;      -- true if a succ fires
  signal token_latch    : unsigned (LogWidth(capacity)-1 downto 0);
  constant U0    : unsigned (LogWidth(capacity)-1 downto 0) := (others => '0');

  signal non_zero       : boolean;

  constant debug_flag : boolean := global_debug_flag;
  
-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- default_arch

  assert capacity > 0 report "in place " & name & ": place must have capacity > 0." severity error;
  assert marking <= capacity report "in place " & name & ": initial marking must be less than place capacity." severity error;

  -- At most one of the preds can send a pulse.
  -- We detect it with an OR over all inputs
  incoming_token <= OrReduce(preds);

  -- At most one of the succs can send a pulse.
  -- We detect it with an OR over all inputs
  backward_reset <= OrReduce(succs);


  CapGtOne: if (capacity > 1) generate
  
    non_zero <= (token_latch /= U0);

    latch_token_cap_gt_one : process (clk, reset,incoming_token, backward_reset, token_latch, non_zero)
	variable incr, decr          : boolean;
    	variable next_token_latch_var: unsigned (token_latch'high downto token_latch'low);
    begin

      incr := incoming_token and (not backward_reset);
      decr := backward_reset and (not incoming_token);
      next_token_latch_var := token_latch;
  
      if(incr) then
          next_token_latch_var := token_latch + 1;
      elsif (decr) then
          next_token_latch_var := token_latch - 1;
      end if;
      
      if clk'event and clk = '1' then  -- rising clock edge

        if reset = '1' then            -- synchronous reset (active high)
          token_latch <= To_Unsigned(marking, token_latch'length);
        else
          token_latch <= next_token_latch_var;
        end if;
  
        if((reset /= '1') and debug_flag and decr) then
             
        	  if (token_latch = 0) then
          		  assert false report "in place-with-bypass: " & name &  ": number of tokens cannot become negative!" severity error;
        	  end if;
           	  assert false report "in place " & name & ": token count decremented from " & Convert_To_String(to_integer(token_latch))
		 	  severity note;
        end if;
  
        if ((reset /= '1') and debug_flag and incr) then
  
       		  if(token_latch = capacity) then
         		  assert false report "in place-with-bypass: " & name & " number of tokens "
			 	  & Convert_To_String(to_integer(token_latch)+1) & " cannot exceed capacity " 
			 	  & Convert_To_String(capacity) severity error;
       		  end if;
           	  assert false report "in place " & name & " token count incremented from " & Convert_To_String(to_integer(token_latch))
		  	  severity note;
	  end if;

      end if;
    end process latch_token_cap_gt_one;
  end generate CapGtOne;


  -- When capacity = 1, we will write this process in a slightly optimized
  -- manner in order to save a flip-flop.
  CapEqOne: if (capacity = 1) generate

    latch_token_cap_eq_one : process (clk, reset,incoming_token, backward_reset, non_zero)
	variable incr, decr          : boolean;
	variable next_non_zero_var        : boolean; 
    begin

      incr := incoming_token and (not backward_reset);
      decr := backward_reset and (not incoming_token);

      next_non_zero_var := non_zero;
  
      if(incr) then
          next_non_zero_var := true;
      elsif (decr) then
          next_non_zero_var := false;
      end if;
      
  
      if clk'event and clk = '1' then  -- rising clock edge

        if reset = '1' then            -- synchronous reset (active high)
          non_zero <= (marking > 0);
        else
          non_zero    <= next_non_zero_var;
        end if;
  
        if((reset /= '1') and debug_flag and decr) then
             
        	  if (not non_zero) then
          		  assert false report "in place-with-bypass: " & name &  ": number of tokens cannot become negative!" severity error;
        	  end if;
           	  assert false report "in place " & name & ": token count decremented from 1 to 0 " severity note;
        end if;
  
        if ((reset /= '1') and debug_flag and incr) then
  
       		  if(non_zero) then
         		  assert false report "in place-with-bypass: " & name & " number of tokens "
			 	  & " cannot exceed capacity " 
			 	  & Convert_To_String(capacity) severity error;
       		  end if;
           	  assert false report "in place " & name & " token count incremented from 0 to 1" severity note;
	  end if;

      end if;
    end process latch_token_cap_eq_one;
  end generate CapEqOne;

  token <= incoming_token or non_zero;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;

-- a short-hand model to implement a merge
-- from transitions to transitions.entity
entity transition_merge is
  generic (name: string);
  port (
    preds      : in   BooleanArray;
    symbol_out : out  boolean);
end transition_merge;

architecture default_arch of transition_merge is
begin  -- default_arch

  -- The transition fires when any of its preds is true.
  symbol_out <= OrReduce(preds);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ahir;
use ahir.Types.all;
use ahir.subprograms.all;

entity transition is
  port (
    preds      : in   BooleanArray;
    symbol_in  : in   boolean;
    symbol_out : out  boolean);
end transition;

architecture default_arch of transition is
begin  -- default_arch

  -- The transition is enabled only when all preds are true.
  symbol_out <= symbol_in and AndReduce(preds);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity BinaryEncoder is
  generic (name:string; iwidth: integer := 3; owidth: integer := 3);
  port(din: in std_logic_vector(iwidth-1 downto 0);
       dout: out std_logic_vector(owidth-1 downto 0));
end BinaryEncoder;


architecture LowLevel of BinaryEncoder is
  signal ival : integer range 0 to iwidth-1;
  constant awidth : integer := Minimum(Maximum(Ceil_Log2(iwidth),1),owidth);
begin  -- LowLevel

  process(din)
    variable ivar : integer range 0 to iwidth-1;
  begin
    ivar := 0;
    for I in 0 to iwidth-1 loop
      if(din(I) = '1') then
        ivar := I;
        exit;
      end if;
    end loop;
    ival <= ivar;
  end process;

  process(ival)
    variable doutvar : std_logic_vector(owidth-1 downto 0);
  begin
    doutvar := (others => '0');
    doutvar(awidth-1 downto 0) := To_SLV(To_Unsigned(ival,awidth));
    dout <= doutvar;
  end process;
    

end LowLevel;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Utilities.all;
use ahir.SubPrograms.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity BranchBase is
  generic (name: string; condition_width: integer := 1; bypass_flag: boolean := false);
  port (condition: in std_logic_vector(condition_width-1 downto 0);
        clk,reset: in std_logic;
        req: in Boolean;
        ack0: out Boolean;
        ack1: out Boolean);
end entity;


architecture Behave of BranchBase is

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin

 noBypass: if not bypass_flag generate
  process(clk)
    variable c_reduce : std_logic;
  begin
    if(clk'event and clk = '1') then
      if(reset = '1') then
        ack0 <= false;
        ack1 <= false;
      elsif req then

	assert(not is_X(condition)) report 
		"branch condition is X" severity error;

        c_reduce := OrReduce(condition);
	
        if(c_reduce = '1') then
          ack1 <= true;
          ack0 <= false;
        else
          ack0 <= true;
          ack1 <= false;
        end if;
      else
        ack0 <= false;
        ack1 <= false;
      end if;
    end if;
  end process;
 end generate noBypass;

 yesBypass: if bypass_flag generate

    process(condition, req)
	variable c_reduce: std_logic;
    begin
        c_reduce := OrReduce(condition);
	if(req) then
		ack0 <= (c_reduce = '0');
		ack1 <= (c_reduce = '1');
	else
		ack0 <= false;
		ack1 <= false;
	end if;
    end process;
 end generate yesBypass;

end Behave;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity FullRateRepeater is
  generic(name : string;  data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity FullRateRepeater;

architecture behave of FullRateRepeater is

-- see comment above..
--##decl_synopsys_sync_set_reset##

       type RepeaterState is (Empty, Full);
       signal repeater_state: RepeaterState;

       signal data_reg: std_logic_vector(data_width-1 downto 0);
begin  -- SimModel

    process(clk, reset, repeater_state, push_req, pop_req, data_in)
	variable nstate: RepeaterState;
	variable push_ack_v, pop_ack_v : std_logic;
	variable load_reg : boolean;
    begin
	
	nstate := repeater_state;
	push_ack_v := '0';
	pop_ack_v  := '0';
	load_reg := false;

	case repeater_state is
		when Empty =>
			push_ack_v := '1';
			if(push_req = '1')  then
				load_reg := true;
				nstate   := Full;
			end if;
		when Full =>
			pop_ack_v := '1';
			if(pop_req = '1') then
				push_ack_v := '1';
				if(push_req = '0') then
					nstate := Empty;
				else
					load_reg := true;
				end if;
			end if;
	end case;

	push_ack <= push_ack_v;
	pop_ack  <= pop_ack_v;
		
	if(clk'event and clk = '1') then
		if(reset = '1') then
			repeater_state <= Empty;
		else
			repeater_state <= nstate;
			if(load_reg) then
				data_reg <= data_in;
			end if;
		end if;
	end if;
    end process;

    data_out <= data_reg;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.OperatorPackage.all;
use ahir.FloatOperatorPackage.all;


library ahir_ieee_proposed;
use ahir_ieee_proposed.float_pkg.all;

entity GenericCombinationalOperator is
  generic
    (
      name: string;
      operator_id   : string := "ApIntAdd";          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer := 4;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer := 0;    -- width of input2
      num_inputs    : integer := 1;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer := 4;          -- width of output.
      constant_operand : std_logic_vector := "0001"; -- constant operand.. (it is always the second operand)
      constant_width: integer := 4;
      use_constant  : boolean := true
      );
  port (
    data_in       : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
    result      : out std_logic_vector(owidth-1 downto 0)
    );
end GenericCombinationalOperator;


architecture Vanilla of GenericCombinationalOperator is
  constant iwidth : integer := iwidth_1 + iwidth_2;
begin  -- Behave

  assert((num_inputs = 1) or (num_inputs = 2)) report "either 1 or 2 inputs" severity failure;

  TwoOperand : if num_inputs = 2 generate
    -- int x int -> int
    TwoOpIntIntInt: if input1_is_int and input2_is_int and output_is_int generate
      process(data_in)
        variable   result_var : std_logic_vector(owidth-1 downto 0);
        variable op1: std_logic_vector(iwidth_1-1 downto 0);
        variable op2: std_logic_vector(iwidth_2-1 downto 0);
      begin
        op1 := data_in(iwidth-1 downto iwidth_2);
        op2 := data_in(iwidth_2-1 downto 0);
        result_var := (others => '0');
        TwoInputOperation(operator_id, op1, op2,result_var);
        result <= result_var;
      end process;
    end generate TwoOpIntIntInt;

    -- float x float -> float
    TwoOpFloatFloatFloat: if (not input1_is_int) and (not input2_is_int) and (not output_is_int) generate
      assert(iwidth_1 = iwidth_2) report "floatXfloat -> float operation: inputs must be of the same width." severity error;
      assert(input1_characteristic_width = input2_characteristic_width) report "floatXfloat -> float operation: input exponent sizes must be the same."
        severity error;
      
      process(data_in)
        variable op1: std_logic_vector(iwidth_1-1 downto 0);
        variable op2: std_logic_vector(iwidth_2-1 downto 0);
        variable   result_var: std_logic_vector(owidth-1 downto 0);
      begin
        op1 := data_in(iwidth-1 downto iwidth_2);
        op2 := data_in(iwidth_2-1 downto 0);
        result_var := (others => '0');
        TwoInputFloatArithOperation(operator_id, op1,op2,input1_characteristic_width, input1_mantissa_width, result_var);
        result <= result_var;
      end process;
    end generate TwoOpFloatFloatFloat;

    -- float x float -> int
    TwoOpFloatFloatInt: if ((not input1_is_int) and (not input2_is_int) and output_is_int) generate
      assert(iwidth_1 = iwidth_2) report "floatXfloat -> int operation: inputs must be of the same width." severity error;
      assert(input1_characteristic_width = input2_characteristic_width) report "floatXfloat -> int operation: input exponent sizes must be the same."
        severity error;
      
      process(data_in)
        variable op1: std_logic_vector(iwidth_1-1 downto 0);
        variable op2: std_logic_vector(iwidth_2-1 downto 0);
        variable   result_var: std_logic_vector(owidth-1 downto 0);        
      begin
        result_var := (others => '0');

	op1 := data_in(iwidth-1 downto iwidth_2);
	op2 := data_in(iwidth_2-1 downto 0);

        TwoInputFloatCompareOperation(operator_id, op1,op2, input1_characteristic_width, input1_mantissa_width, result_var);
        result <= result_var;
      end process;
    end generate TwoOpFloatFloatInt;

    -- float x int -> * and int x float -> * are not permitted.
    assert(input1_is_int = input2_is_int) report "both operands of two input operators should be either ints or floats"
      severity failure;

    -- int x int -> float is not permitted.
    assert((not input1_is_int) or output_is_int) report "if the inputs to a two-input operation are ints, the output cannot be a float!" severity failure;

  end generate TwoOperand;


  SingleOperandNoConstant : if num_inputs = 1 and not use_constant generate

    SingleOperandNoConstantIntInt: if input1_is_int and output_is_int generate
      process(data_in)
        variable   result_var    : std_logic_vector(owidth-1 downto 0);
      begin
        result_var := (others => '0');
        SingleInputOperation(operator_id, data_in, result_var);
        result <= result_var;
      end process;
    end generate SingleOperandNoConstantIntInt;
    
    SingleOperandNoConstantFloatFloat: if (not input1_is_int) and (not output_is_int) generate

      -- the resize operation is to be treated specially, since
      -- there are two different conversions..
      ResizeFloat: if (operator_id = "ApFloatResize") generate

        Trivial: if ((output_mantissa_width = input1_mantissa_width) and
			(output_characteristic_width = input1_characteristic_width)) generate
		result <= data_in;
	end generate Trivial;

        NonTrivial: if ((output_mantissa_width /= input1_mantissa_width) or
			(output_characteristic_width /= input1_characteristic_width)) generate
          process(data_in)
            variable op1: std_logic_vector(iwidth_1-1 downto 0);
            variable   result_var: std_logic_vector(owidth-1 downto 0);                
          begin
            op1 := data_in;
            result_var := (others => '0');
            ApFloatResize_proc(To_Float(op1, input1_characteristic_width, input1_mantissa_width),
                               output_characteristic_width,
                               output_mantissa_width,
                               result_var);
            result <= result_var;
          end process;        
	end generate NonTrivial;
      end generate ResizeFloat;

      NotResizeFloat: if (operator_id /= "ApFloatResize") generate
        
        process(data_in)
          variable op1: std_logic_vector(iwidth_1-1 downto 0);
          variable   result_var: std_logic_vector(owidth-1 downto 0);                
        begin
          op1 := data_in;
          result_var := (others => '0');
          SingleInputFloatOperation(operator_id, op1, input1_characteristic_width, input1_mantissa_width, result_var);
          result <= result_var;
        end process;
      end generate NotResizeFloat;
      
    end generate SingleOperandNoConstantFloatFloat;

    SingleOperandNoConstantFloatInt: if (not input1_is_int) and output_is_int generate
      process(data_in)
        variable op1: std_logic_vector(iwidth_1-1 downto 0);
        variable   result_var: std_logic_vector(owidth-1 downto 0);                
      begin
        op1 := data_in;
        result_var := (others => '0');
        SingleInputFloatOperation(operator_id, op1, input1_characteristic_width, input1_mantissa_width, result_var);
        result <= result_var;
      end process;
    end generate SingleOperandNoConstantFloatInt;

    SingleOperandNoConstantIntFloat: if (input1_is_int) and (not output_is_int) generate
      process(data_in)
        variable   result_var: std_logic_vector(owidth-1 downto 0);                
      begin
        result_var := (others => '0');
        SingleInputFloatOperation(operator_id, data_in, output_characteristic_width, output_mantissa_width, result_var);
        result <= result_var;
      end process;
    end generate SingleOperandNoConstantIntFloat;
  end generate SingleOperandNoConstant;

  SingleOperandWithConstant : if num_inputs = 1 and use_constant generate

    SingleOperandWithConstantIntInt: if input1_is_int and output_is_int generate
      SigBlock: block
        signal op2_sig : std_logic_vector(constant_width-1 downto 0);
      begin  -- block SigBlock
        -- TODO: changes here.
        op2_sig <= constant_operand;

        process(data_in,op2_sig)
          variable   result_var    : std_logic_vector(owidth-1 downto 0);
        begin
          result_var := (others => '0');
          TwoInputOperation(operator_id,
                            data_in,
                            op2_sig,
                            result_var); 
          result <= result_var;
        end process;
      end block SigBlock;
    end generate SingleOperandWithConstantIntInt;

    SingleOperandWithConstantFloatInt: if (not input1_is_int) and output_is_int generate

      SigBlock: block
      	signal op2_sig: std_logic_vector(constant_width-1 downto 0);
      begin
      op2_sig <= constant_operand;
      process(data_in, op2_sig)
        variable   result_var: std_logic_vector(owidth-1 downto 0);                        
      begin
        result_var := (others => '0');
       	TwoInputFloatCompareOperation(operator_id, data_in, op2_sig,input1_characteristic_width, input1_mantissa_width, result_var);
        result <= result_var;
      end process;
      end block SigBlock;
    end generate SingleOperandWithConstantFloatInt;

    SingleOperandWithConstantFloatFloat: if (not input1_is_int) and (not output_is_int) generate
      SigBlock: block
      	signal op2_sig: std_logic_vector(constant_width-1 downto 0);
      begin
      op2_sig <= constant_operand;
      process(data_in, op2_sig)
        variable   result_var: std_logic_vector(owidth-1 downto 0);                        
      begin
        result_var := (others => '0');
       	TwoInputFloatArithOperation(operator_id, data_in, op2_sig, input1_characteristic_width, input1_mantissa_width, result_var);
        result <= result_var;
      end process;
    end block SigBlock;
    end generate SingleOperandWithConstantFloatFloat;
  end generate SingleOperandWithConstant;
  
end Vanilla;



------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- if guards(I) is true, let the handshake proceed, else
-- shunt it.  This interface is inserted in between the
-- req/ack signals from/to the CP and the operators in the
-- datapath.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity GuardInterface is
	generic (nreqs: integer; delay_flag:boolean);
	port (reqL: in BooleanArray(nreqs-1 downto 0);
	      ackL: out BooleanArray(nreqs-1 downto 0); 
	      reqR: out BooleanArray(nreqs-1 downto 0);
	      ackR: in BooleanArray(nreqs-1 downto 0); 
	      guards: in std_logic_vector(nreqs-1 downto 0);
	      clk: in std_logic;
	      reset: in std_logic);
end entity;


architecture Behave of GuardInterface is
	signal ackL_un_guarded: BooleanArray(nreqs-1 downto 0);
begin

	process(reqL,ackR,guards,ackL_un_guarded)
	begin
		for I in 0 to nreqs-1 loop
			if(guards(I) = '1') then
				reqR(I) <= reqL(I);
				ackL(I) <= ackR(I);
			else
				reqR(I) <= false;
				ackL(I) <= ackL_un_guarded(I);
			end if;
		end loop;
	end process;

	nodelay: if not delay_flag generate
		ackL_un_guarded <= reqL;
	end generate nodelay;

	yesdelay: if delay_flag generate
		process(clk)
		begin
			if(clk'event and clk = '1') then 
				if(reset = '1') then
					ackL_un_guarded <= (others => false);
				else
					ackL_un_guarded <= reqL;
				end if;
			end if;
		end process;
	end generate yesdelay;

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity InputMuxBaseNoData is
  generic (name: string;
	   twidth: integer;
	   nreqs: integer;
	   no_arbitration: Boolean := false);
  port (
    -- req/ack follow pulse protocol
    reqL                 : in  BooleanArray(nreqs-1 downto 0);
    ackL                 : out BooleanArray(nreqs-1 downto 0);
    -- output side req/ack level protocol
    reqR                 : out std_logic;
    ackR                 : in  std_logic;
    -- tag specifies the requester index 
    tagR                : out std_logic_vector(twidth-1 downto 0);
    clk, reset          : in std_logic);
end InputMuxBaseNoData;


architecture Behave of InputMuxBaseNoData is

  signal reqP,ackP,ssig : std_logic_vector(nreqs-1 downto 0);
  signal fEN: std_logic_vector(nreqs-1 downto 0);  

  constant tag0 : std_logic_vector(twidth-1 downto 0) := (others => '0');

  -- one-cycle delay between req and ack => in order to break long
  -- combinational (false) paths.
  constant suppress_immediate_ack : BooleanArray(reqL'length-1 downto 0) := (others => true);
begin  -- Behave


  -----------------------------------------------------------------------------
  -- pulse to level translate
  -----------------------------------------------------------------------------
  P2L: for I in nreqs-1 downto 0 generate
      P2LBlk: block
      begin  -- block P2L          
        p2Linst: Pulse_To_Level_Translate_Entity
	   generic map (name => name & "-p2Linst-" & Convert_To_String(I))
          port map (rL => reqL(I), rR => reqP(I), aL => ackL(I), aR => ackP(I),
                                 clk => clk, reset => reset);
      end block P2LBlk;

  end generate P2L;
  


  -----------------------------------------------------------------------------
  -- priority encoding or pass through
  -----------------------------------------------------------------------------
  NoArbitration: if no_arbitration generate
    fEN <= reqP;
    reqR <= OrReduce(fEN);
    ackP <= fEN when ackR = '1' else (others => '0');
  end generate NoArbitration;

  Arbitration: if not no_arbitration generate
    rpeInst: Request_Priority_Encode_Entity
      generic map (name => name & "-rpeInst", num_reqs => reqP'length)
      port map( clk => clk,
                reset => reset,
                reqR => reqP,
                ackR => ackP,
                forward_enable => fEN,
                req_s => reqR,
                ack_s => ackR);
    
  end generate Arbitration;

  -----------------------------------------------------------------------------
  -- tag generation
  -----------------------------------------------------------------------------
  taggen : BinaryEncoder generic map (
    name => name & "-taggen", 
    iwidth => nreqs,
    owidth => twidth)
    port map (
      din  => fEN,
      dout => tagR);

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity InputMuxBase is
  generic (name: string; iwidth: integer := 10;
	   owidth: integer := 10;
	   twidth: integer := 3;
	   nreqs: integer := 1;
	   no_arbitration: Boolean := false;
	   registered_output: Boolean := true);
  port (
    -- req/ack follow pulse protocol
    reqL                 : in  BooleanArray(nreqs-1 downto 0);
    ackL                 : out BooleanArray(nreqs-1 downto 0);
    dataL                : in  std_logic_vector(iwidth-1 downto 0);
    -- output side req/ack level protocol
    reqR                 : out std_logic;
    ackR                 : in  std_logic;
    dataR                : out std_logic_vector(owidth-1 downto 0);
    -- tag specifies the requester index 
    tagR                : out std_logic_vector(twidth-1 downto 0);
    clk, reset          : in std_logic);
end InputMuxBase;


architecture Behave of InputMuxBase is

  signal reqP,ackP,fEN : std_logic_vector(nreqs-1 downto 0);

  type WordArray is array (natural range <>) of std_logic_vector(owidth-1 downto 0);
  signal dataP : WordArray(nreqs-1 downto 0);

  constant tag0 : std_logic_vector(twidth-1 downto 0) := (others => '0');

  -- one-cycle delay between req and ack => in order to break long
  -- combinational (false) paths.
  constant suppress_immediate_ack : BooleanArray(reqL'length-1 downto 0) := (others => true);

  -- intermediate signals.
  signal reqR_sig                : std_logic;
  signal ackR_sig                : std_logic;
  signal dataR_sig               : std_logic_vector(owidth-1 downto 0);
  signal tagR_sig                : std_logic_vector(twidth-1 downto 0);
  signal fair_reqP, fair_ackP    : std_logic_vector(nreqs-1 downto 0);

begin  -- Behave


  assert(iwidth = owidth*nreqs) report "mismatched i/o widths in InputMuxBase" severity error;

  -----------------------------------------------------------------------------
  -- "fairify" the level-reqs.
  -----------------------------------------------------------------------------
  fairify: NobodyLeftBehind generic map (name=> name & "-fairify", num_reqs => nreqs)
		port map (clk => clk, reset => reset, reqIn => reqP, ackOut => ackP,
					reqOut => fair_reqP, ackIn => fair_ackP);


  -----------------------------------------------------------------------------
  -- output queue if registered_output is set.
  -----------------------------------------------------------------------------
  OutputRepeater: if registered_output generate

    -- purpose: output queue
    OqBlock: block
      signal oq_data_in : std_logic_vector((twidth + owidth)-1 downto 0);
      signal oq_data_out : std_logic_vector((twidth + owidth)-1 downto 0);
    begin  -- block OqBlock

      oq_data_in <= dataR_sig & tagR_sig;
      dataR <= oq_data_out((twidth+owidth)-1 downto twidth);
      tagR <= oq_data_out(twidth-1 downto 0);

        
      oqueue : QueueBase generic map (
        name => name & "-oqueue",
        queue_depth => 2,
        data_width  => twidth + owidth)
        port map (
          clk      => clk,
          reset    => reset,
          data_in  => oq_data_in,
          push_req => reqR_sig,
          push_ack => ackR_sig,
          data_out => oq_data_out,
          pop_ack  => reqR,
          pop_req  => ackR);
      
    end block OqBlock;
  end generate OutputRepeater;

  NoOutputRepeater: if not registered_output generate
    
    dataR <= dataR_sig;
    reqR <= reqR_sig;
    ackR_sig <= ackR;
    tagR <= tagR_sig;
    
  end generate NoOutputRepeater;
  
  -----------------------------------------------------------------------------
  -- pulse to level translate
  -----------------------------------------------------------------------------
  P2L: for I in nreqs-1 downto 0 generate
    p2Linstance: Pulse_To_Level_Translate_Entity
      generic map (name => name & "-p2Linstance-" & Convert_To_String(I))
      port map(rL => reqL(I), rR => reqP(I), aL => ackL(I), aR => ackP(I),
               clk => clk, reset => reset);     

    process(dataL)
      variable regv : std_logic_vector(owidth-1 downto 0);
    begin
      Extract(dataL,I,regv);
      dataP(I) <= regv;
    end process;
    
  end generate P2L;

  -----------------------------------------------------------------------------
  -- priority encoding or pass through
  -----------------------------------------------------------------------------
  NoArbitration: if no_arbitration generate
    fEN <= fair_reqP;
    reqR_sig <= OrReduce(fEN);
    fair_ackP <= fEN when ackR_sig = '1' else (others => '0');
  end generate NoArbitration;

  Arbitration: if not no_arbitration generate
    fEN <= PriorityEncode(fair_reqP);
    reqR_sig <= OrReduce(fEN);
    fair_ackP <= fEN when ackR_sig = '1' else (others => '0');
  end generate Arbitration;

  -----------------------------------------------------------------------------
  -- final multiplexor
  -----------------------------------------------------------------------------
  process(fEN,dataP)
  begin
    dataR_sig <= (others => '0');
    for J in 0 to nreqs-1 loop
      if(fEN(J) = '1') then
        dataR_sig <= dataP(J);
        exit;
      end if;
    end loop;
  end process;    

  -----------------------------------------------------------------------------
  -- tag generation
  -----------------------------------------------------------------------------
  taggen : BinaryEncoder generic map (
    name => name & "-taggen",
    iwidth => nreqs,
    owidth => twidth)
    port map (
      din  => fEN,
      dout => tagR_sig);

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity InputPortLevelNoData is
  
  generic (num_reqs: integer; 
	no_arbitration: boolean := false);
  port (
    -- ready/ready interface with the requesters
    req       : in  std_logic_vector(num_reqs-1 downto 0);
    ack       : out std_logic_vector(num_reqs-1 downto 0);
    -- ready/ready interface with outside world
    oreq       : out std_logic;
    oack       : in  std_logic;
    clk, reset : in  std_logic);
  
end InputPortLevelNoData;

architecture default_arch of InputPortLevelNoData is

  signal req_active, ack_sig  : std_logic_vector(num_reqs-1 downto 0); 
  
begin  -- default_arch

  oreq <= OrReduce(req_active);

  NoArb: if no_arbitration generate
    req_active <= req;
  end generate NoArb;

  Arb: if not no_arbitration generate
    req_active <= PriorityEncode(req);
  end generate Arb;

  gen: for I in num_reqs-1 downto 0 generate

    ack_sig(I) <= req_active(I) and oack; 
    
    ack(I) <= ack_sig(I);
    
  end generate gen;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity InputPortLevel is
  
  generic (name: string;
	num_reqs: integer := 5; 
	data_width: integer := 8;  
	no_arbitration: boolean := false);
  port (
    -- ready/ready interface with the requesters
    req       : in  std_logic_vector(num_reqs-1 downto 0);
    ack       : out std_logic_vector(num_reqs-1 downto 0);
    data      : out std_logic_vector((num_reqs*data_width)-1 downto 0);
    -- ready/ready interface with outside world
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : in  std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
  
end InputPortLevel;

architecture default_arch of InputPortLevel is

  
  type IPWArray is array(integer range <>) of std_logic_vector(data_width-1 downto 0);
  signal data_final, data_reg : IPWArray(num_reqs-1 downto 0);
  signal req_active, ack_sig  : std_logic_vector(num_reqs-1 downto 0); 
  
  
begin  -- default_arch

  oreq <= OrReduce(req_active);

  NoArb: if no_arbitration generate
    req_active <= req;
  end generate NoArb;

  Arb: if not no_arbitration generate
    req_active <= PriorityEncode(req);
  end generate Arb;

  process(data_final)
    variable ldata: std_logic_vector((num_reqs*data_width)-1 downto 0);
  begin

    for J in 0 to num_reqs-1 loop
       ldata(((J+1)*data_width)-1 downto (J*data_width)) := data_final(J);
    end loop;

    data <= ldata;
  end process;

  gen: for I in num_reqs-1 downto 0 generate

    SingleReq: if (num_reqs = 1) generate 
    	ack_sig(I) <=  oack; 
    end generate SingleReq;

    MultipleReqs: if (num_reqs > 1) generate
    	ack_sig(I) <= req_active(I) and oack; 
    end generate MultipleReqs;
    
    ack(I) <= ack_sig(I);
    
    data_final(I) <= odata;
    
  end generate gen;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- a level to pulse translator used at the
-- output end of a data-path operator in order
-- to interface to the control path.
-- Madhav Desai.
entity Level_To_Pulse_Translate_Entity is
  generic (name : string);
  port(
	rL : out std_logic;
        rR : in  boolean;
        aL : in std_logic;
        aR : out boolean;
        clk : in std_logic;
        reset : in std_logic);
end entity;

architecture Behave of Level_To_Pulse_Translate_Entity is
  type L2PState is (Idle,WaitForAckL);
  signal l2p_state : L2PState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  process(clk, reset, aL, rR, l2p_state)
    variable nstate : L2PState;
  begin
    nstate := l2p_state;
    rL <= '0';
    aR <= false;

    case l2p_state is
        when Idle =>
          if(rR) then
              nstate := WaitForAckL;
          end if;
        when WaitForAckL =>
          rL <= '1';
          if(aL = '1') then
            aR <= true;
	    if(rR)  then
               nstate := WaitForAckL;
            else
               nstate := Idle;
	    end if;
          end if; 
        when others => null;
      end case;

    if(clk'event and clk = '1') then
	if reset = '1' then
		l2p_state <= Idle;
	else
      		l2p_state <= nstate;
	end if;
    end if;
  end process;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity LoadCompleteShared is
    generic
    (
      name : string;
      data_width: integer := 8;
      tag_length:  integer := 1;
      num_reqs : integer := 1;
      no_arbitration: boolean := false;
      detailed_buffering_per_output: IntegerArray
    );
  port (
    -- req/ack follow level protocol
    reqR                     : in BooleanArray(num_reqs-1 downto 0);
    ackR                     : out BooleanArray(num_reqs-1 downto 0);
    dataR                    : out std_logic_vector((data_width*num_reqs)-1 downto 0);
    -- output data consists of concatenated pairs of ops.
    mdata                    : in std_logic_vector(data_width-1 downto 0);
    mreq                     : out  std_logic;
    mack                     : in std_logic;
    mtag                     : in std_logic_vector(tag_length-1 downto 0);
    -- with dataR
    clk, reset              : in std_logic);
end LoadCompleteShared;

architecture Vanilla of LoadCompleteShared is

begin  -- Behave


  odemux: OutputDeMuxBaseWithBuffering
    generic map (
      name => name & "-odemux ",
      iwidth => data_width,
      owidth =>  data_width*num_reqs,
      twidth =>  tag_length,
      nreqs  => num_reqs,
      detailed_buffering_per_output => detailed_buffering_per_output,
      full_rate => true )   -- always double buffered.
    port map (
      reqL   => mack,                   -- cross-over (mack from mem-subsystem)
      ackL   => mreq,                   -- cross-over 
      dataL =>  mdata,
      tagL  =>  mtag,
      reqR  => reqR,
      ackR  => ackR,
      dataR => dataR,
      clk   => clk,
      reset => reset);
  
  
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity LoadReqShared is
  generic
    (
	name: string;
	addr_width: integer := 8;
      	num_reqs : integer := 1; -- how many requesters?
	tag_length: integer := 1;
	no_arbitration: Boolean := false;
        min_clock_period: Boolean := true;
	time_stamp_width: integer := 0
    );
  port (
    -- req/ack follow pulse protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    -- concatenated address corresponding to access
    dataL                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
    -- address to memory
    maddr                   : out std_logic_vector((addr_width)-1 downto 0);
    mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);

    mreq                    : out std_logic;
    mack                    : in std_logic;
    -- clock, reset (active high)
    clk, reset              : in std_logic);
end LoadReqShared;

architecture Vanilla of LoadReqShared is

  constant iwidth: integer := addr_width*num_reqs;
  constant owidth: integer := addr_width;

  constant debug_flag : boolean := false;
-- constant registered_output : boolean := min_clock_period and (time_stamp_width = 0);

  -- must register..  ack implies that address has been sampled.
  constant registered_output : boolean := true; 

  signal imux_tag_out: std_logic_vector(tag_length-1 downto 0);
  
begin  -- Behave
  assert(tag_length >= Ceil_Log2(num_reqs)) report "insufficient tag width" severity error;

  TstampGen: if time_stamp_width > 0 generate

    Tstamp: block
	signal time_stamp: std_logic_vector(time_stamp_width-1 downto 0);
    begin 
    	mtag <= imux_tag_out & time_stamp; 


	-- ripple counter.
	process(clk)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				time_stamp <= (others => '0');
			else
				for I in 1 to time_stamp_width-1 loop
					time_stamp(I) <= time_stamp(I) xor AndReduce(time_stamp(I-1 downto 0));
				end loop;
				time_stamp(0) <= not time_stamp(0);
			end if;
		end if;
	end process;
    end block;
    
  end generate TstampGen;

  NoTstampGen: if time_stamp_width < 1 generate
	mtag <= imux_tag_out;
  end generate NoTstampGen;

  -- xilinx xst does not like this assertion...
  -- DbgAssert: if debug_flag generate
    -- assert( (not ((reset = '0') and (clk'event and clk = '1') and no_arbitration)) or Is_At_Most_One_Hot(reqL))
      -- report "in no-arbitration case, at most one request should be hot on clock edge (in SplitOperatorShared)" severity error;    
  -- end generate DbgAssert;

  
  imux: InputMuxBase
    generic map(name => name & "-imux",
		iwidth => iwidth,
                owidth => owidth, 
                twidth => tag_length,
                nreqs => num_reqs,
                no_arbitration => no_arbitration,
                registered_output => registered_output)
    port map(
      reqL       => reqL,
      ackL       => ackL,
      dataL      => dataL,
      reqR       => mreq,
      ackR       => mack,
      dataR      => maddr,
      tagR       => imux_tag_out,
      clk        => clk,
      reset      => reset);
  
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##


-- make sure that there is no starvation..
--
-- latch the incoming requests (reqIn) and present them
-- to the downstream user (reqOut).  As ackIn is received,
-- clear reqOut.  The latching of reqIn to reqOut is done
-- only if reqOut is cleared.  There is a bypass path
-- from reqIn to reqOut if reqIn_register is 0..  This
-- prevents a useless latency.
entity NobodyLeftBehind is
  generic ( name: string; num_reqs : integer := 1);
  port (
    clk,reset : in std_logic;
    reqIn : in std_logic_vector(num_reqs-1 downto 0);
    ackOut: out std_logic_vector(num_reqs-1 downto 0);
    reqOut : out std_logic_vector(num_reqs-1 downto 0);
    ackIn : in std_logic_vector(num_reqs-1 downto 0));
end entity;


architecture Fair of NobodyLeftBehind is
  signal reqIn_register: std_logic_vector(num_reqs-1 downto 0);
  signal reqIn_reg_is_non_zero: std_logic;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave


   -- if there is only one requester, there is really no point.
   Trivial: if num_reqs = 1 generate
     reqOut <= reqIn;
     ackOut <= ackIn;
   end generate Trivial;

   Nontrivial: if num_reqs > 1 generate

     reqIn_reg_is_non_zero <= OrReduce(reqIn_register);
     reqOut <= reqIn_register when reqIn_reg_is_non_zero = '1' else reqIn;
     
     process(clk, reset, reqIn_reg_is_non_zero, reqIn_register, reqIn, ackIn)
	  variable next_reqIn_register : std_logic_vector(num_reqs-1 downto 0);
     begin
	  next_reqIn_register := reqIn_register;
  
          if(reqIn_reg_is_non_zero = '0') then
              -- if reqIn_register is 0, then reqIn will be 
	      -- immediately forwarded to reqOut..  An ackIn
              -- may immediately appear.. in which case reqIn_register
              -- will stay 0.
	      next_reqIn_register := reqIn and (not ackIn); -- reqIn and (reqIn xor ackIn);
          else
              -- reqOut must come from reqIn_register.. the next
              -- state will be determined by reqIn_register and ackIn
	      next_reqIn_register := reqIn_register and (not ackIn); -- reqIn_register and (reqIn_register xor ackIn);
          end if;
  
          if(clk'event and clk = '1') then
		  if(reset = '1') then
			  reqIn_register <= (others => '0');
		  else
			  reqIn_register <= next_reqIn_register;
		  end if;
	  end if;
	  
     end process;

     ackOut <= ackIn;
   
   end generate NonTrivial;

end Fair;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##


-- does nothing really...
entity NullRepeater is
  generic(name : string;  data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity NullRepeater;

architecture behave of NullRepeater is

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- SimModel

   push_ack <= pop_req;
   pop_ack  <= push_req;
   data_out <= data_in;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity OutputDeMuxBaseNoData is
  generic(name : string;
          twidth: integer;
	  nreqs: integer;
	  detailed_buffering_per_output: IntegerArray);
  port (
    -- req/ack follow level protocol
    reqL                 : in  std_logic;
    ackL                 : out std_logic;
    -- tag identifies index to which demux
    -- should happen
    tagL                 : in std_logic_vector(twidth-1 downto 0);
    -- reqR/ackR follow pulse protocol
    -- and are of length n
    reqR                : in BooleanArray(nreqs-1 downto 0);
    ackR                : out  BooleanArray(nreqs-1 downto 0);
    clk, reset          : in std_logic);
end OutputDeMuxBaseNoData;

architecture Behave of OutputDeMuxBaseNoData is
  signal ackL_sig : std_logic_vector(nreqs-1 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  assert detailed_buffering_per_output'length = reqR'length report "Mismatch." severity failure;

  -----------------------------------------------------------------------------
  -- parallel generate across all requesters
  -----------------------------------------------------------------------------
  PGen: for I in reqR'range generate
    RegFSM: block
      signal valid: std_logic;
      signal lhs_clear : std_logic;
      signal rhs_state : std_logic;

      signal lhs_state : unsigned ((Ceil_Log2(detailed_buffering_per_output(I)+1))-1 downto 0); 
      signal lhs_valid: Boolean;

      signal aR, aR_reg: Boolean;

    begin  -- block Reg
      
      ---------------------------------------------------------------------------
      -- valid true if this I is mentioned in tag
      ---------------------------------------------------------------------------
      valid <= '1' when (reqL = '1') and (I = To_Integer(To_Unsigned(tagL))) else '0';

      ---------------------------------------------------------------------------
      -- lhs-state machine.. just a 3 bit counter which counts up everytime
      -- there is a valid input to this index, and down when the req appears 
      -- at the receiver end.
      ---------------------------------------------------------------------------
      process(clk,lhs_state, lhs_clear,reset,valid)
        variable nstate : unsigned ((Ceil_Log2(detailed_buffering_per_output(I)+1))-1 downto 0); 
        variable aL_var : std_logic;
	variable lhs_valid_var: Boolean;
      begin
        nstate := lhs_state;
        aL_var := '0';
        lhs_valid_var := false;
        
        if(lhs_state < detailed_buffering_per_output(I)) then
            aL_var := '1';
            if(valid = '1') then
              nstate := lhs_state + 1;
            end if;
        end if;

        if(nstate > 0) then
	    lhs_valid_var := true;
            if(lhs_clear = '1') then
              nstate := nstate-1;
            end if;
	end if;

        ackL_sig(I) <= aL_var;
        lhs_valid   <= lhs_valid_var;
        
        if(clk'event and clk = '1') then
           if(reset = '1') then
	      lhs_state <= (others => '0');
	   else
              lhs_state <= nstate;
           end if;        
        end if;

      end process;

      -------------------------------------------------------------------------
      -- rhs state machine
      -------------------------------------------------------------------------
     process(clk,rhs_state,reset,reqR(I),lhs_valid)
       variable nstate : std_logic;
       variable aR_var: boolean;
       variable lhs_clear_var : std_logic;
     begin
        nstate := rhs_state;
        aR_var     := false;
        lhs_clear_var := '0';
        
        case rhs_state is
          when '0' =>
            if(reqR(I)) then
	      nstate := '1';
            end if;
          when '1' =>
            if(lhs_valid) then
              aR_var := true;
              lhs_clear_var := '1';
	      if (not reqR(I)) then
                 nstate := '0';
	      end if;
            end if;
          when others => null;
        end case;

        lhs_clear <= lhs_clear_var;
        ackR(I) <= aR_var;
        
        if(clk'event and clk = '1') then
	  if(reset = '1') then 
          	rhs_state <= '0';
	  else
          	rhs_state <= nstate;
	  end if;
        end if;
     end process;
    end block RegFSM;
    
  end generate PGen;

  -----------------------------------------------------------------------------
  -- ackL
  -----------------------------------------------------------------------------
  ackL <= OrReduce(ackL_sig);

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-------------------------------------------------------------------------------
-- a single level requester on the left, and nreq requesters on the right.
--
-- reqR -> ackR has unit delay if pipeline_flag is true.
-- reqL -> ackL has at least a unit delay.
-------------------------------------------------------------------------------
entity OutputDeMuxBase is
  generic(name: string; iwidth: integer := 4;
	  owidth: integer := 12;
	  twidth: integer := 2;
	  nreqs: integer := 3;
	  no_arbitration: Boolean := false;
          pipeline_flag: Boolean := true);
  port (
    -- req/ack follow level protocol
    reqL                 : in  std_logic;
    ackL                 : out std_logic;
    dataL                : in  std_logic_vector(iwidth-1 downto 0);
    -- tag identifies index to which demux
    -- should happen
    tagL                 : in std_logic_vector(twidth-1 downto 0);
    -- reqR/ackR follow pulse protocol
    -- and are of length n
    reqR                : in BooleanArray(nreqs-1 downto 0);
    ackR                : out  BooleanArray(nreqs-1 downto 0);
    -- dataR is array(n,m) 
    dataR               : out std_logic_vector(owidth-1 downto 0);
    clk, reset          : in std_logic);
end OutputDeMuxBase;

architecture Behave of OutputDeMuxBase is

  type WordArray is array (natural range <>) of std_logic_vector(iwidth-1 downto 0);
  signal dfinal, dfinal_reg: WordArray(nreqs-1 downto 0);

  signal ackL_sig : std_logic_vector(nreqs-1 downto 0);
  signal ackR_sig : BooleanArray(nreqs-1 downto 0);
  
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  assert(owidth = iwidth*nreqs) report "word-length mismatch in output demux " & name severity failure;

  
  -----------------------------------------------------------------------------
  -- parallel generate across all requesters
  -----------------------------------------------------------------------------
  PGen: for I in reqR'range generate
    RegFSM: block
      signal valid: std_logic;
      signal lhs_clear : std_logic;
      signal rhs_state, lhs_state : std_logic;
    begin  -- block Reg
      
      ---------------------------------------------------------------------------
      -- valid true if this I is mentioned in tag
      ---------------------------------------------------------------------------
      valid <= '1' when (reqL = '1') and (I = To_Integer(To_Unsigned(tagL))) else '0';

      ---------------------------------------------------------------------------
      -- lhs-state machine.
      ---------------------------------------------------------------------------
      process(clk,lhs_state, lhs_clear,reset,valid)
        variable nstate : std_logic;
        variable latch_flag : boolean;
        variable aL_var : std_logic;
      begin
        nstate := lhs_state;
        latch_flag := false;
        aL_var := '0';
        
        case lhs_state is
          when '0' =>
            if(valid = '1') then
              nstate := '1';
              latch_flag := true;
              aL_var := '1';
            end if;
          when '1' =>
            if(lhs_clear = '1') then
              nstate := '0';
            end if;

	    -- to track down some mixup issues!
	    assert (valid = '0') report "In Outputdemux " & name & ": stalled request " & Convert_To_String(I)
			severity warning;

          when others => null;
        end case;

        ackL_sig(I) <= aL_var;
        
        if(clk'event and clk = '1') then
	  if(reset = '1') then
		lhs_state <= '0';
	  else
            	lhs_state <= nstate;
          end if;

          if(latch_flag) then
            dfinal(I) <= dataL;
          end if;          
        end if;
      end process;

      -------------------------------------------------------------------------
      -- rhs state machine
      -------------------------------------------------------------------------
     process(clk,rhs_state,reset,reqR(I),lhs_state)
       variable nstate : std_logic;
       variable aR_var : boolean;
       variable lhs_clear_var : std_logic;
     begin
        nstate := rhs_state;
        aR_var := false;
        lhs_clear_var := '0';
        
        case rhs_state is
          when '0' =>
            if(reqR(I)) then
              if(lhs_state = '1') then
                aR_var := true;
                lhs_clear_var := '1';
              else
                nstate := '1';
              end if;
            end if;
          when '1' =>
            if(lhs_state = '1') then
              lhs_clear_var := '1';
              aR_var := true;
              nstate := '0';
            end if;
          when others => null;
        end case;

        ackR_sig(I) <= aR_var;
        lhs_clear <= lhs_clear_var;
        
        if(clk'event and clk = '1') then
	  if(reset = '1') then
		rhs_state <= '0';
	  else
          	rhs_state <= nstate;
	  end if;
        end if;
     end process;
    end block RegFSM;
    
  end generate PGen;

  -----------------------------------------------------------------------------
  -- ackL
  -----------------------------------------------------------------------------
  ackL <= OrReduce(ackL_sig);

  -----------------------------------------------------------------------------
  -- non-pipelined case, ackR_sig goes straight to ackR, dfinal goes to dataR
  -----------------------------------------------------------------------------
  Nonpipelined: if (not pipeline_flag) generate

    ackR <= ackR_sig;

    process(dfinal)
      variable dataRv : std_logic_vector(owidth-1 downto 0);
    begin
      for I in dfinal'range loop
	dataRv(((I+1)*iwidth)-1 downto I*iwidth) := dfinal(I);
        --Insert(dataRv,I,dfinal(I));
      end loop;
      dataR <= dataRv;
    end process;
    
  end generate Nonpipelined;  

  -----------------------------------------------------------------------------
  -- pipelined case, ackR_sig delayed to ackR, dfinal delayed to dataR
  -----------------------------------------------------------------------------
  Pipelined: if pipeline_flag generate

    process(clk,reset)
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          ackR <= (others => false);
        else
          ackR <= ackR_sig;
        end if;
      end if;
    end process;

    Freggen: for I in 0 to nreqs-1 generate
      process(clk)
      begin
        if(clk'event and clk = '1') then
          if(ackR_sig(I)) then
            dfinal_reg(I) <= dfinal(I);
          end if;
        end if;
      end process;
    end generate Freggen;

    process(dfinal_reg)
      variable dataRv : std_logic_vector(owidth-1 downto 0);
    begin
      for I in dfinal_reg'range loop
	dataRv(((I+1)*iwidth)-1 downto I*iwidth) := dfinal_reg(I);
        -- Insert(dataRv,I,dfinal_reg(I));
      end loop;
      dataR <= dataRv;
    end process;
  end generate Pipelined;

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-------------------------------------------------------------------------------
-- a single level requester on the left, and nreq requesters on the right.
--
-- reqR -> ackR can be zero delay.
-- reqL -> ackL has at least a unit delay
--
-- This demux provides buffering for each output.
-- (potentially useful in loop-pipelining).
-------------------------------------------------------------------------------
entity OutputDeMuxBaseWithBuffering is
  generic(name: string;
          iwidth: integer := 4;
	  owidth: integer := 12;
	  twidth: integer := 2;
	  nreqs: integer := 3;
	  detailed_buffering_per_output: IntegerArray;
	  full_rate: boolean);
  port (
    -- req/ack follow level protocol
    reqL                 : in  std_logic;
    ackL                 : out std_logic;
    dataL                : in  std_logic_vector(iwidth-1 downto 0);
    -- tag identifies index to which demux
    -- should happen
    tagL                 : in std_logic_vector(twidth-1 downto 0);
    -- reqR/ackR follow pulse protocol
    -- and are of length n
    reqR                : in BooleanArray(nreqs-1 downto 0);
    ackR                : out  BooleanArray(nreqs-1 downto 0);
    -- dataR is array(n,m) 
    dataR               : out std_logic_vector(owidth-1 downto 0);
    clk, reset          : in std_logic);
end OutputDeMuxBaseWithBuffering;

architecture Behave of OutputDeMuxBaseWithBuffering is
  signal ackL_array : std_logic_vector(nreqs-1 downto 0);
  --alias buffer_sizes: IntegerArray(detailed_buffering_per_output'length-1 downto 0) is detailed_buffering_per_output;

begin  -- Behave
  assert(owidth = iwidth*nreqs) report "word-length mismatch in output demux " & name severity failure;

  bufGen: for I in 0 to nreqs-1 generate

    -- purpose: instantiate a buffer
    BufBlock: block
      signal write_req,write_ack : std_logic;
      signal unload_req,unload_ack : boolean;
      signal buf_data_in, buf_data_out : std_logic_vector(iwidth-1 downto 0);
      signal valid : std_logic;
      signal has_data: std_logic;

    begin  -- block BufBlock

       ub : UnloadBuffer generic map (
         name => name & " buffer " & Convert_To_String(I),
         buffer_size => detailed_buffering_per_output(I),
         data_width  => iwidth, 
	 bypass_flag => false,
	 use_unload_register => true)
         port map (
           write_req  => write_req,
           write_ack  => write_ack,
           write_data => buf_data_in,
           unload_req => unload_req,
           unload_ack => unload_ack,
           read_data  => buf_data_out,
           has_data   => has_data,
           clk        => clk,
           reset      => reset);

      
      ---------------------------------------------------------------------------
      -- valid true if this I is mentioned in tag
      ---------------------------------------------------------------------------
      valid <= '1' when (reqL = '1') and (I = To_Integer(To_Unsigned(tagL))) else '0';
      write_req <= valid;
      ackL_array(I) <= write_ack when (valid = '1') else '0';

      -------------------------------------------------------------------------
      -- dataL goes to each buffer.
      -------------------------------------------------------------------------
      buf_data_in <= dataL;


      -------------------------------------------------------------------------
      -- unload side is straightforward
      -------------------------------------------------------------------------
      unload_req <= reqR(I);
      ackR(I) <= unload_ack;
      dataR(((I+1)*iwidth)-1 downto I*iwidth) <= buf_data_out;
      
    end block BufBlock;
  end generate bufGen;

  -- ack is OrReduced from the Demux combinations.
  ackL <= OrReduce(ackL_array);
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity OutputPortLevelNoData is
  generic(name: string; num_reqs: integer;
	no_arbitration: boolean := false);
  port (
    req       : in  std_logic_vector(num_reqs-1 downto 0);
    ack       : out std_logic_vector(num_reqs-1 downto 0);
    oreq       : out std_logic;
    oack       : in  std_logic;
    clk, reset : in  std_logic);
end entity;

architecture Base of OutputPortLevelNoData is
  signal req_active, ack_sig , fair_reqs, fair_acks : std_logic_vector(num_reqs-1 downto 0);
begin
  
  fairify: NobodyLeftBehind generic map(name => name & "-fairify", num_reqs => num_reqs)
		port map(clk => clk, reset => reset,
				reqIn => req,
				ackOut => ack,
				reqOut => fair_reqs,
				ackIn => fair_acks);
  
  oreq <= OrReduce(req_active);

  NoArb: if no_arbitration generate
     req_active <= fair_reqs;
  end generate NoArb;

  Arb: if not no_arbitration generate
     req_active <= PriorityEncode(fair_reqs);
  end generate Arb;

  gen: for I in num_reqs-1 downto 0 generate
       ack_sig(I) <= req_active(I) and oack; 
       fair_acks(I) <= ack_sig(I);
  end generate gen;

end Base;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;

entity OutputPortLevel is
  generic(name: string; num_reqs: integer;
	data_width: integer;
	no_arbitration: boolean := true);
  port (
    req       : in  std_logic_vector(num_reqs-1 downto 0);
    ack       : out std_logic_vector(num_reqs-1 downto 0);
    data      : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : out std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
end entity;

architecture Base of OutputPortLevel is
  
  type OPWArray is array(integer range <>) of std_logic_vector(odata'range);
  signal data_array : OPWArray(num_reqs-1 downto 0);
  signal req_active, ack_sig , fair_reqs, fair_acks : std_logic_vector(num_reqs-1 downto 0);
  
begin

  fairify: NobodyLeftBehind generic map(name => name & "-fairify", num_reqs => num_reqs)
		port map(clk => clk, reset => reset,
				reqIn => req,
				ackOut => ack,
				reqOut => fair_reqs,
				ackIn => fair_acks);
  
  oreq <= OrReduce(req_active);

  NoArb: if no_arbitration generate
     req_active <= fair_reqs;
  end generate NoArb;

  Arb: if not no_arbitration generate
     req_active <= PriorityEncode(fair_reqs);
  end generate Arb;

  process (data_array)
    variable var_odata : std_logic_vector(data_width-1 downto 0) := (others => '0');
  begin  -- process
    var_odata := (others => '0');
    for I in 0 to num_reqs-1 loop
      var_odata := data_array(I) or var_odata;
    end loop;  -- I
    odata <= var_odata;
  end process;

  gen: for I in num_reqs-1 downto 0 generate

       debugGen: if global_pipe_report_flag generate
	process(clk)
	begin
		if(clk'event and clk = '1') then
			if (reset = '0') then
				if((req_active(I) = '1')  and (ack_sig(I) = '1')) then
					assert false report "RPIPE " & name & "requester=" &
						Convert_To_String(I) & " data=" &
							Convert_SLV_to_Hex_String(data_array(I)) severity note;
				end if;
			end if;
		end if;
	end process;
       end generate debugGen;

       SingleReq: if (num_reqs = 1) generate
          ack_sig(I) <=  oack; 
       	  data_array(I) <= data;
       end generate SingleReq;

       MultipleReq: if (num_reqs > 1) generate
          ack_sig(I) <= req_active(I) and oack; 
       	  process(data,req_active(I))
             variable target: std_logic_vector(data_width-1 downto 0);
          begin
            if(req_active(I) = '1') then
		target := data(((I+1)*data_width)-1 downto I*data_width);
		--Extract(data,I,target);
	    else
		target := (others => '0');
	    end if;	
       	    data_array(I) <= target;
          end process;
       end generate MultipleReq;

         
       fair_acks(I) <= ack_sig(I);
  end generate gen;

end Base;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity PhiBase is
  generic (
    name: string;
    num_reqs   : integer;
    data_width : integer;
    bypass_flag : boolean := false);
  port (
    req                 : in  BooleanArray(num_reqs-1 downto 0);
    ack                 : out Boolean;
    idata               : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
    odata               : out std_logic_vector(data_width-1 downto 0);
    clk, reset          : in std_logic);
end PhiBase;



architecture Behave of PhiBase is
   signal muxed_idata: std_logic_vector(data_width-1 downto 0);
   signal odata_reg: std_logic_vector(data_width-1 downto 0);
   signal there_is_a_req: boolean;
   signal ack_internal: boolean;
   signal req_registered, final_req : BooleanArray(num_reqs-1 downto 0);
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  assert(idata'length = (odata'length * req'length)) report "data size mismatch in PhiBase " & name severity failure;

  -- muxed data..
  odata <= MuxOneHot(idata,final_req);

  there_is_a_req <= OrReduce(req);
  ack_internal <= there_is_a_req;

  process(clk)
	variable mux_data : std_logic_vector(odata'length-1 downto 0);
  begin
     if(clk'event and clk = '1') then
	if(reset = '1') then
          req_registered <= (others => false);
	elsif (there_is_a_req) then
	  req_registered <= req;
	end if;
     end if;
  end process;

  -- bypass.
  Byp: if bypass_flag generate
  	final_req <= req when there_is_a_req else req_registered;
        ack <= ack_internal;
  end generate Byp;

  -- no-bypass.
  NoByp: if (not bypass_flag) generate
	final_req <= req_registered;
        process(clk)
        begin
 	   if(clk'event and clk = '1') then
		if(reset = '1') then
			ack <= false;
		else 
			ack <= ack_internal;
		end if;
	   end if;
        end process;
  end generate NoByp;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;

--
-- base Pipe.
--   Implementation guarantees registering of every in->out path
--   unless save_slot flag is true, in which case there will be
--   a combi path from write_req -> read_ack.
--

entity PipeBase is
  generic (name : string;
	   num_reads: integer;
           num_writes: integer;
           data_width: integer;
           lifo_mode: boolean := false;
           depth: integer := 1;
	   signal_mode: boolean := false;
           shift_register_mode: boolean := false;
	   save_slot: boolean := false;
	   bypass: boolean := false;
	   full_rate: boolean);
  port (
    read_req       : in  std_logic_vector(num_reads-1 downto 0);
    read_ack       : out std_logic_vector(num_reads-1 downto 0);
    read_data      : out std_logic_vector((num_reads*data_width)-1 downto 0);
    write_req       : in  std_logic_vector(num_writes-1 downto 0);
    write_ack       : out std_logic_vector(num_writes-1 downto 0);
    write_data      : in std_logic_vector((num_writes*data_width)-1 downto 0);
    clk, reset : in  std_logic);
  
end PipeBase;

architecture default_arch of PipeBase is

  signal pipe_data, pipe_data_repeated : std_logic_vector(data_width-1 downto 0);
  signal pipe_req, pipe_ack, pipe_req_repeated, pipe_ack_repeated: std_logic;
  signal signal_data : std_logic_vector(data_width-1 downto 0); 
  signal written_at_least_once: std_logic;

  --
  -- shallow => will be implemented using flip-flops.  Can be expensive!
  --
  constant shallow_flag : boolean :=    (depth < global_pipe_shallowness_threshold);
  -- constant shallow_flag : boolean :=   true;
  
  signal write_ack_sig: std_logic_vector(num_writes-1 downto 0);
  signal read_ack_sig: std_logic_vector(num_reads-1 downto 0);
  signal read_data_sig: std_logic_vector((num_reads*data_width)-1 downto 0);

begin  -- default_arch

 write_ack <= write_ack_sig;
 read_ack  <= read_ack_sig;
  
 read_data <= read_data_sig;
 debugGen: if global_pipe_report_flag generate
	-- super useful for tracing.

  process (clk)
	variable wvar : std_logic_vector(data_width-1 downto 0);
	variable rvar : std_logic_vector(data_width-1 downto 0);
  begin
	if(clk'event and clk = '1') then
		if(reset = '0') then
			for I in  0 to num_writes-1 loop
				wvar := write_data (((I+1)*data_width)-1 downto  I*data_width);
				if(write_req(I)= '1' and  write_ack_sig(I) = '1') then
					assert false report "WPIPE " & name & " requester=" & Convert_To_String(I) & " data= " & 
								Convert_SLV_to_Hex_String(wvar) severity note;
				end if;
			end loop;
			for J in  0 to num_reads-1 loop
				rvar := read_data_sig (((J+1)*data_width)-1 downto  J*data_width);
				if(read_req(J)= '1' and  read_ack_sig(J) = '1') then
					assert false report "RPIPE " & name & " requester=" & Convert_To_String(J) & " data= " & 
								Convert_SLV_to_Hex_String(rvar) severity note;
				end if;
			end loop;
		end if;
	end if;
  end process;
  end generate debugGen;

  manyWriters: if (num_writes > 1) generate
    wmux : OutputPortLevel generic map (
      name => name & "-wmux",
      num_reqs       => num_writes,
      data_width     => data_width,
      no_arbitration => false)
      port map (
        req   => write_req,
        ack   => write_ack_sig,
        data  => write_data,
        oreq  => pipe_req,                -- no cross-over, drives req
        oack  => pipe_ack,                -- no cross-over, receives ack
        odata => pipe_data,
        clk   => clk,
        reset => reset);
  end generate manyWriters;

  singleWriter: if (num_writes = 1) generate
    pipe_req <= write_req(0);
    write_ack_sig(0) <= pipe_ack;
    pipe_data <= write_data;
  end generate singleWriter;
 
  -- in signal mode, the pipe is just a flag
  SignalMode: if signal_mode generate

     -- write always succeeds.
     pipe_ack <= '1';
     process(clk,reset) 
     begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			signal_data <= (others => '0');	
  			written_at_least_once <= '0';
		else
			if(pipe_req = '1') then
				signal_data <= pipe_data;
  				written_at_least_once <= '1';
			end if;
		end if;
	end if;
     end process;

     ReaderGen: for R in 0 to num_reads-1 generate
	read_ack_sig(R) <= '1'; -- read-ack always succeeds..
	read_data_sig(((R+1)*data_width)-1 downto (R*data_width)) <= signal_data;
     end generate ReaderGen;

  end generate SignalMode;

  Shallow: if (not signal_mode) and shallow_flag and (not lifo_mode) generate

     saveSlot: if save_slot and (depth > 0) generate
      queue : QueueBaseSaveSlot generic map (	
        name => name & "-queue",	
        queue_depth => depth,
        data_width       => data_width)
        port map (
          push_req   => pipe_req,
          push_ack => pipe_ack,
          data_in  => pipe_data,
          pop_req  => pipe_req_repeated,
          pop_ack  => pipe_ack_repeated,
          data_out => pipe_data_repeated,
          clk      => clk,
          reset    => reset);
     end generate saveSlot;

     notSaveSlot: if ((not save_slot) and (not bypass)) or (depth = 0) generate

      queue : QueueBase generic map (	
        name => name & "-queue",	
        queue_depth => depth,
        data_width       => data_width)
        port map (
          push_req   => pipe_req,
          push_ack => pipe_ack,
          data_in  => pipe_data,
          pop_req  => pipe_req_repeated,
          pop_ack  => pipe_ack_repeated,
          data_out => pipe_data_repeated,
          clk      => clk,
          reset    => reset);
     end generate notSaveSlot;

     bypassCase: if (not save_slot) and bypass and (depth > 0) generate

      queue : QueueWithBypass generic map (	
        name => name & "-queue",	
        queue_depth => depth,
        data_width       => data_width)
        port map (
          push_req   => pipe_req,
          push_ack => pipe_ack,
          data_in  => pipe_data,
          pop_req  => pipe_req_repeated,
          pop_ack  => pipe_ack_repeated,
          data_out => pipe_data_repeated,
          clk      => clk,
          reset    => reset);
     end generate bypassCase;
  end generate Shallow;

  DeepFifo: if (not signal_mode) and (not shallow_flag) and (not lifo_mode) generate
    
   notShiftReg: if (not shift_register_mode) generate
    queue : SynchFifoWithDPRAM generic map (
      name => name & "-queue", 
      queue_depth => depth,
      data_width       => data_width)
      port map (
        push_req   => pipe_req,
        push_ack => pipe_ack,
        data_in  => pipe_data,
        pop_req  => pipe_req_repeated,
        pop_ack  => pipe_ack_repeated,
        data_out => pipe_data_repeated,
        nearly_full => open,
        clk      => clk,
        reset    => reset);
   end generate notShiftReg;
    
   shiftReg: if shift_register_mode generate
      srqueue : ShiftRegisterQueue generic map (	
        name => name & "-srqueue",	
        queue_depth => depth,
        data_width       => data_width)
        port map (
          push_req   => pipe_req,
          push_ack => pipe_ack,
          data_in  => pipe_data,
          pop_req  => pipe_req_repeated,
          pop_ack  => pipe_ack_repeated,
          data_out => pipe_data_repeated,
          clk      => clk,
          reset    => reset);
   end generate shiftReg;
 
  end generate DeepFifo;

  Lifo: if (not signal_mode) and  lifo_mode generate
    stack : SynchLifo generic map (
      name => name & "-stack",
      queue_depth => depth,
      data_width       => data_width)
      port map (
        push_req   => pipe_req,
        push_ack => pipe_ack,
        data_in  => pipe_data,
        pop_req  => pipe_req_repeated,
        pop_ack  => pipe_ack_repeated,
        data_out => pipe_data_repeated,
        nearly_full => open,
        clk      => clk,
        reset    => reset);
  end generate Lifo;
  

  manyReaders: if  (not signal_mode) and (num_reads > 1) generate
    rmux : InputPortLevel generic map (
	name => name & "-rmux",
      num_reqs       => num_reads,
      data_width     => data_width,
      no_arbitration => false)
      port map (
        req => read_req,
        ack => read_ack_sig,
        data => read_data_sig,
        oreq => pipe_req_repeated,       
        oack => pipe_ack_repeated,       
        odata => pipe_data_repeated,
        clk => clk,
        reset => reset);
  end generate manyReaders;

  singleReader: if  (not signal_mode) and (num_reads = 1) generate
    read_ack_sig(0) <= pipe_ack_repeated;
    pipe_req_repeated <= read_req(0);
    read_data_sig <= pipe_data_repeated;
  end generate singleReader;
  
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

--
-- in pull_mode, rL/aL accepts data which is sent by rR/aR.
-- rL -> rR is 0 delay, but aR -> aL MUST have a delay.
--
entity Pulse_To_Level_Translate_Entity is
  generic (name: string);
  port( rL : in boolean;
        rR : out std_logic;
        aL : out boolean;
        aR : in std_logic;
        clk : in std_logic;
        reset : in std_logic);
end entity;

architecture Behave of Pulse_To_Level_Translate_Entity is
  type PullModeState is (Idle,Ack,Waiting);
  signal pull_mode_state : PullModeState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  process(clk, rL, aR, pull_mode_state)
    variable nstate : PullModeState;
  begin
    nstate := pull_mode_state;
    rR <= '0';
    aL <= false;

      case pull_mode_state is
        when Idle =>
          if(rL) then
            rR <= '1';
            if(aR = '1') then
              nstate := Ack;
            else
              nstate := Waiting;
            end if;
          end if;
        when Ack =>
          aL <= true;
          if(rL) then
            rR <= '1' ;
	    if(aR = '0')  then
               	nstate := Waiting;
	    end if;
          else
            nstate := Idle;
          end if; 
        when Waiting =>
	  rR <= '1';
          if(aR = '1') then
            nstate := Ack;
          end if;
        when others => null;
      end case;

    if(clk'event and clk = '1') then
	if reset = '1' then
		pull_mode_state <= Idle;
	else
      		pull_mode_state <= nstate;
	end if;
    end if;
  end process;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity QueueBase is
  generic(name : string; queue_depth: integer := 1; data_width: integer := 32;
		save_one_slot: boolean := false);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity QueueBase;

architecture behave of QueueBase is

  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- SimModel

 --
 -- 0-depth queue is just a set of wires.
 --
 triv: if queue_depth = 0 generate
	push_ack <= pop_req;
	pop_ack  <= push_req;
	data_out <= data_in;
 end generate triv;

 qD1: if (queue_depth = 1) generate
   RB: block
      signal full_flag: boolean;
      signal data_reg: std_logic_vector(data_width-1 downto 0);

   begin

      push_ack <= '1' when (not full_flag) else '0';
      pop_ack  <= '1' when full_flag else '0';
      data_out <= data_reg;

      process(clk, reset, push_req, pop_req, full_flag, data_in, data_reg)
	variable next_full_flag_var: boolean;
        variable next_data_reg_var: std_logic_vector(data_width-1 downto 0);
      begin
	next_full_flag_var := full_flag;
        next_data_reg_var := data_reg;

        if (full_flag) then
           if (pop_req = '1') then
              next_full_flag_var := false;
           end if;
        else 
           if (push_req = '1') then
               next_full_flag_var := true;
               next_data_reg_var :=  data_in;
	   end if;
         end if;
  
       if (clk'event and clk='1') then
         if(reset  = '1') then
            full_flag <= false;
            data_reg <= (others => '0');
         else
             full_flag <= next_full_flag_var;
	     data_reg  <= next_data_reg_var;
         end if;
      end if;
     end process;
   end block;
 end generate qD1;


 qDGt1: if queue_depth > 1 generate 
  NTB: block 
   signal queue_array : QueueArray(queue_depth-1 downto 0);
   signal read_pointer, write_pointer: unsigned ((Ceil_Log2(queue_depth))-1 downto 0);
   signal next_read_pointer, next_write_pointer, write_pointer_plus_1: unsigned ((Ceil_Log2(queue_depth))-1 downto 0);

  constant URW0: unsigned ((Ceil_Log2(queue_depth))-1 downto 0):= (others => '0');

  signal full_flag, empty_flag: boolean;
  signal queue_size : unsigned ((Ceil_Log2(queue_depth+1))-1 downto 0);
  signal incr_read_pointer, incr_write_pointer: boolean;
  signal incr_queue_size, decr_queue_size: boolean;

  signal write_flag : boolean;
  signal eq_flag: boolean;

  begin
 
    assert (not full_flag) report "Queue " & name & " is full." severity note;

    write_pointer_plus_1 <= (others => '0') when (write_pointer = queue_depth-1) else (write_pointer+1);

    push_ack <= '1' when (not full_flag) else '0';
    pop_ack  <= '1' when (not empty_flag) else '0';

    -- next read pointer, write pointer.
    process(incr_read_pointer, read_pointer) 
    begin
	if(incr_read_pointer) then
		if(read_pointer = queue_depth-1) then
			next_read_pointer <= (others => '0');
		else
			next_read_pointer <= read_pointer + 1;
		end if;
	else
		next_read_pointer <= read_pointer;
	end if;
    end process;
    rdpReg: SynchResetRegisterUnsigned generic map (name => name & ":rpreg", data_width => read_pointer'length)
		port map (clk => clk, reset => reset, din => next_read_pointer, dout => read_pointer);

    process(incr_write_pointer, write_pointer, write_pointer_plus_1) 
    begin
	if(incr_write_pointer) then
		next_write_pointer <= write_pointer_plus_1;
	else
		next_write_pointer <= write_pointer;
	end if;
    end process;

    -- empty/full logic.
    eq_flag <= (next_read_pointer = next_write_pointer);
    fe_logic: QueueEmptyFullLogic 
	port map (clk => clk, reset => reset, 
			read => incr_read_pointer, write => incr_write_pointer,
				eq_flag => eq_flag,
				full => full_flag, empty => empty_flag);

    wrpReg: SynchResetRegisterUnsigned generic map (name => name & ":wrpreg", data_width => write_pointer'length)
		port map (clk => clk, reset => reset, din => next_write_pointer, dout => write_pointer);

    -- bottom pointer gives the data in FIFO mode..
    process (read_pointer, queue_array)
	variable data_out_var : std_logic_vector(data_width-1 downto 0);
    begin
	data_out_var := (others =>  '0');
        for I in 0 to queue_depth-1 loop
	    if(I = To_Integer(read_pointer)) then
    		data_out_var := queue_array(I);
	    end if;
	end loop;
	data_out <= data_out_var;
    end process;

    -- write to queue-array.
    Wgen: for W in 0 to queue_depth-1 generate
       process(clk, reset, write_flag, write_pointer, data_in) 
       begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
                             queue_array(W) <= (others => '0');
			elsif (write_flag and (W = write_pointer)) then
			     queue_array(W) <= data_in;
			end if;
		end if;
       end process;
    end generate Wgen;
  
    -- single process..  Synopsys mangles the logic... split it into two.
    process(read_pointer, write_pointer, empty_flag, full_flag, push_req, pop_req)
      variable push,pop : boolean;
    begin
      push  := false;
      pop   := false;
      
      if((not full_flag) and push_req = '1') then
          push := true;
      end if;
  
      if((not empty_flag) and pop_req = '1') then
          pop := true;
      end if;
  
      incr_read_pointer <= pop;
      incr_write_pointer <= push;
  
      write_flag <= push;
    end process;

   end block NTB;
  end generate qDGt1;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.GlobalConstants.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity QueueBaseWithEmptyFull is
  generic(name : string; 
		queue_depth: integer := 1; 
		reverse_bypass_flag: boolean := false;
		data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       empty, full: out std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity QueueBaseWithEmptyFull;

architecture behave of QueueBaseWithEmptyFull is

  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);

  signal base_push_req: std_logic;
  signal base_push_ack: std_logic;

  signal base_pop_req: std_logic;
  signal base_pop_ack: std_logic;

  signal base_empty: boolean;
  signal base_full: boolean;

  signal base_data_out: std_logic_vector(data_width-1 downto 0);
-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- SimModel

 pDZero:  if(queue_depth = 0) generate

	empty <= '1';
	full  <= '1';

	data_out <= data_in;

	push_ack <= pop_req;
	pop_ack  <= push_req;

 end generate pDZero;


 oSideQGt0: if (queue_depth > 0)  generate

     base_push_req <= push_req;
     push_ack <= base_push_ack;
     base_pop_req <= pop_req;
     pop_ack <= base_pop_ack;

     data_out <= base_data_out;

     empty <= '1' when base_empty else '0';
     full  <= '1' when base_full else '0';

 end generate oSideQGt0;

 qD1: if (queue_depth = 1) generate
   rbypGen: if reverse_bypass_flag generate
   RB: block
      signal full_flag: boolean;
      signal data_reg: std_logic_vector(data_width-1 downto 0);
   begin

      base_empty <= not full_flag;
      base_full  <= full_flag;

      base_push_ack <= '1' when (not full_flag) or (base_pop_req = '1')  else '0';
      base_pop_ack  <= '1' when full_flag else '0';
	
      base_data_out <= data_reg;

      process(clk, reset, base_push_req, base_pop_req, full_flag, data_in, data_reg)
	variable next_full_flag_var: boolean;
        variable next_data_reg_var: std_logic_vector(data_width-1 downto 0);
      begin
	next_full_flag_var := full_flag;
        next_data_reg_var := data_reg;

        if (full_flag) then
           if (base_pop_req = '1') then
		if(base_push_req = '1') then
               		next_data_reg_var :=  data_in;
		else
              		next_full_flag_var := false;
		end if;
           end if;
        else 
           if (base_push_req = '1') then
               next_full_flag_var := true;
               next_data_reg_var :=  data_in;
	   end if;
         end if;
  
       if (clk'event and clk='1') then
         if(reset  = '1') then
            full_flag <= false;
            data_reg <= (others => '0');
         else
             full_flag <= next_full_flag_var;
	     data_reg  <= next_data_reg_var;
         end if;
      end if;
     end process;
   end block;
   end generate rbypGen;

   not_rbypGen: if not reverse_bypass_flag generate
   RB: block
      signal full_flag: boolean;
      signal data_reg: std_logic_vector(data_width-1 downto 0);
   begin

      base_empty <= not full_flag;
      base_full  <= full_flag;

      base_push_ack <= '0' when full_flag else '1';
      base_pop_ack  <= '1' when full_flag else '0';
	
      base_data_out <= data_reg;

      process(clk, reset, base_push_req, base_pop_req, full_flag, data_in, data_reg)
	variable next_full_flag_var: boolean;
        variable next_data_reg_var: std_logic_vector(data_width-1 downto 0);
      begin
	next_full_flag_var := full_flag;
        next_data_reg_var := data_reg;

        if (full_flag) then
           if (base_pop_req = '1') then
              next_full_flag_var := false;
           end if;
        else 
           if (base_push_req = '1') then
               next_full_flag_var := true;
               next_data_reg_var :=  data_in;
	   end if;
         end if;
  
       if (clk'event and clk='1') then
         if(reset  = '1') then
            full_flag <= false;
            data_reg <= (others => '0');
         else
             full_flag <= next_full_flag_var;
	     data_reg  <= next_data_reg_var;
         end if;
      end if;
     end process;
   end block;
   end generate not_rbypGen;
 end generate qD1;


 qDGt1: if queue_depth > 1 generate 
  NTB: block 
   signal read_pointer, write_pointer, write_pointer_plus_1: unsigned ((Ceil_Log2(queue_depth))-1 downto 0);
   signal next_read_pointer, next_write_pointer: unsigned ((Ceil_Log2(queue_depth))-1 downto 0);

  constant URW0: unsigned ((Ceil_Log2(queue_depth))-1 downto 0):= (others => '0');

  signal incr_read_pointer, incr_write_pointer: boolean;
  signal write_flag : boolean;
  signal write_enable : std_logic;
  signal eq_flag : boolean;

  begin

    -- empty/full logic.
    eq_flag <= (next_read_pointer = next_write_pointer);
    fe_logic: QueueEmptyFullLogic 
	port map (clk => clk, reset => reset, 
			read => incr_read_pointer, write => incr_write_pointer,
				eq_flag => eq_flag,
				full => base_full, empty => base_empty);


    -- next read pointer, write pointer.
    process(incr_read_pointer, read_pointer) 
    begin
	if(incr_read_pointer) then
		if(read_pointer = queue_depth-1) then
			next_read_pointer <= (others => '0');
		else
			next_read_pointer <= read_pointer + 1;
		end if;
	else
		next_read_pointer <= read_pointer;
	end if;
    end process;
    rdpReg: SynchResetRegisterUnsigned generic map (name => name & ":rpreg", data_width => read_pointer'length)
		port map (clk => clk, reset => reset, din => next_read_pointer, dout => read_pointer);

    write_pointer_plus_1 <= (others => '0') when (write_pointer = queue_depth-1) else (write_pointer + 1);
    process(incr_write_pointer, write_pointer, write_pointer_plus_1) 
    begin
	if(incr_write_pointer) then
		next_write_pointer <= write_pointer_plus_1;
	else
		next_write_pointer <= write_pointer;
	end if;
    end process;
    wrpReg: SynchResetRegisterUnsigned generic map (name => name & ":wrpreg", data_width => write_pointer'length)
		port map (clk => clk, reset => reset, din => next_write_pointer, dout => write_pointer);

  -----------------------------------------  declared the array if not distrib ram case ------------------------
  notDistribRam: if not global_use_vivado_distributed_ram_queue generate
    QueueArrayBlock: block
   	signal queue_array : QueueArray(queue_depth-1 downto 0);
    begin 
        -- bottom pointer gives the data in FIFO mode..
        process (read_pointer, queue_array)
	    variable data_out_var : std_logic_vector(data_width-1 downto 0);
        begin
	    data_out_var := (others =>  '0');
            for I in 0 to queue_depth-1 loop
	        if(I = To_Integer(read_pointer)) then
    		    data_out_var := queue_array(I);
	        end if;
	    end loop;
	    base_data_out <= data_out_var;
        end process;

        -- write to queue-array.
        Wgen: for W in 0 to queue_depth-1 generate
           process(clk, reset, write_flag, write_pointer, data_in) 
           begin
		    if(clk'event and (clk = '1')) then
			    if(reset = '1') then
                                 queue_array(W) <= (others => '0');
			    elsif (write_flag and (W = write_pointer)) then
			         queue_array(W) <= data_in;
			    end if;
		    end if;
           end process;
        end generate Wgen;
    end block QueueArrayBlock;
  end generate notDistribRam;
  -----------------------------------------  end non distrib ram case -------------------------------------------

  -----------------------------------------  begin distrib ram case   -------------------------------------------
  write_enable <= '1' when write_flag else '0';
  DistribRam: if global_use_vivado_distributed_ram_queue generate
      distrib_ram_inst:
		fifo_mem_synch_write_asynch_read 
			generic map (name => name & ":distribRam", 
					address_width => read_pointer'length,
					data_width => data_width,
					mem_size => queue_depth)
			port map (
					write_enable => write_enable,
					write_data => data_in,
					write_address => std_logic_vector(write_pointer),
					read_data => base_data_out,
					read_address => std_logic_vector(read_pointer),
					clk => clk
				);
  end generate DistribRam;
  -----------------------------------------  end distrib ram case   -------------------------------------------
  
   not_rbypGen: if not reverse_bypass_flag generate

    base_push_ack <= '0' when base_full else '1';
    base_pop_ack  <= '0' when base_empty else '1';

    -- single process..  Synopsys mangles the logic... split it into two.
    process(base_empty, base_full, base_push_req, base_pop_req)
      variable push,pop : boolean;
    begin
      push  := false;
      pop   := false;
      
      if((not base_full) and base_push_req = '1') then
          push := true;
      end if;
  
      if((not base_empty) and base_pop_req = '1') then
          pop := true;
      end if;
  
      incr_read_pointer <= pop;
      incr_write_pointer <= push;
  
      write_flag <= push;
    end process;
   end generate not_rbypGen;

   rbypGen: if reverse_bypass_flag generate

    base_push_ack <= '1' when (not base_full) or (base_pop_req = '1')  else '0';
    base_pop_ack  <= '0' when base_empty else '1';

    -- single process..  Synopsys mangles the logic... split it into two.
    process(base_empty, base_full, base_push_req, base_pop_req)
      variable push,pop : boolean;
    begin
      push  := false;
      pop   := false;
      
      if(((base_pop_req = '1') or (not base_full)) and base_push_req = '1') then
          push := true;
      end if;
  
      if((not base_empty) and base_pop_req = '1') then
          pop := true;
      end if;
  
      incr_read_pointer <= pop;
      incr_write_pointer <= push;
  
      write_flag <= push;
    end process;
   end generate rbypGen;

   end block NTB;
  end generate qDGt1;

end behave;
library ieee;
use ieee.std_logic_1164.all;

entity QueueEmptyFullLogic is
	port (clk, reset: in std_logic;
		read,write,eq_flag: in boolean;
		full, empty: out boolean);
end entity;

architecture FSM of QueueEmptyFullLogic is

    type QFsmState is (EMPTYSTATE, INBETWEENSTATE, FULLSTATE);
    signal fsm_state: QFsmState;

begin
    
    process(clk, reset, fsm_state, read, write, eq_flag)
	variable ptrs_equal: boolean;
	variable next_fsm_state : QFsmState;
	variable full_var, empty_var: boolean;
    begin
	ptrs_equal := eq_flag;
	next_fsm_state := fsm_state;
	full_var := false;
	empty_var := false;
	case fsm_state is
		when EMPTYSTATE =>
			empty_var := true;
			if(write and (not read)) then
				next_fsm_state := INBETWEENSTATE;
			end if;
		when INBETWEENSTATE =>
			if(read and (not write) and
					ptrs_equal) then
				next_fsm_state := EMPTYSTATE;
			elsif ((not read) and write and
					ptrs_equal) then
				next_fsm_state := FULLSTATE;
			end if;
		when FULLSTATE => 
			full_var := true;
			if(read and (not write)) then
				next_fsm_state := INBETWEENSTATE;
			end if;
	end case;

	full <= full_var;
	empty <= empty_var;
			
			
 	if(clk'event and clk ='1') then
		if(reset = '1') then
			fsm_state <= EMPTYSTATE;
		else
			fsm_state <= next_fsm_state;
		end if;
	end if;

    end process;
end architecture FSM;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.Utilities.all;

entity QueueWithBypass is
  generic(name : string; queue_depth: integer := 1; data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity QueueWithBypass;

architecture behave of QueueWithBypass is

	signal number_of_elements_in_queue: unsigned( (Ceil_Log2(queue_depth+2))-1 downto 0); 

	signal qpush_req, qpush_ack, qpop_req, qpop_ack: std_logic;
	signal qdata_in, qdata_out: std_logic_vector(data_width-1 downto 0);

	signal qhas_data: Boolean;
	signal bypass_active : Boolean;

	signal empty, full: std_logic;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- SimModel

  assert (queue_depth > 0) report "QueueWithBypass "  &  name  & " must have depth > 0 "
				severity failure;

  qhas_data <= (empty = '0');

  -- queue will always accept if there is room.
  -- but it is possible that the accepted data goes 
  -- straight to the output.
  push_ack <= '1' when (full = '0') else '0';
 
  qinst: QueueBaseWithEmptyFull 
		generic map (name => name & "-qbase", queue_depth => queue_depth, data_width => data_width)
		port map (clk => clk, reset => reset, empty => empty, full => full,
				data_in => qdata_in, push_req => qpush_req, push_ack => qpush_ack,
				data_out => qdata_out, pop_req => qpop_req, pop_ack => qpop_ack);

  -- bypass is active?
  bypass_active <= (not qhas_data) and (pop_req = '1');

  -- push into the queue when queue-has-data = '1' or when the world does not care
  qpush_req <= push_req  when (not bypass_active) else  '0';
  qdata_in  <= data_in;

  -- pop from queue when queue-has-data = '1'.
  data_out <= qdata_out when qhas_data else data_in;
  qpop_req <= pop_req   when qhas_data else '0';
  
  -- Note: the forward path from push_req to pop_ack!
  pop_ack  <= qpop_ack  when qhas_data else push_req;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.Utilities.all;
use ahir.Subprograms.all;

-- a simple register
entity RegisterBase is
  generic(name: string; in_data_width: integer; out_data_width: integer);
  port(din: in std_logic_vector(in_data_width-1 downto 0);
       dout: out std_logic_vector(out_data_width-1 downto 0);
       req: in boolean;
       ack: out boolean;
       clk,reset: in std_logic);
end RegisterBase;


architecture arch of RegisterBase is
  constant min_data_width : integer := Minimum(in_data_width,out_data_width);
  signal out_reg : std_logic_vector(min_data_width-1 downto 0);
begin
  process(din,req,reset,clk)
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          ack <= false;
          out_reg <= (others => '0');
        elsif req then
          ack <= true;
          out_reg <= din(min_data_width-1 downto 0);
        else
          ack <= false;
        end if;
      end if;
  end process;

  process(out_reg)
  begin
	dout <= (others => '0');
	dout(min_data_width-1 downto 0) <= out_reg;
  end process;

end arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity Request_Priority_Encode_Entity is
  generic (
    name: string;
    num_reqs : integer := 1;
    pull_mode : boolean := false);
  port (
    clk,reset : in std_logic;
    reqR : in std_logic_vector(num_reqs-1 downto 0);
    forward_enable: out std_logic_vector(num_reqs-1 downto 0);
    ackR: out std_logic_vector(num_reqs-1 downto 0);
    req_s : out std_logic;
    ack_s : in std_logic);
end entity;

architecture Behave of Request_Priority_Encode_Entity is

  signal req_fsm_state : std_logic;
  signal reqR_priority_encoded : std_logic_vector(num_reqs-1 downto 0);
  signal reqR_fresh: std_logic_vector(num_reqs-1 downto 0);
  signal there_is_a_fresh_request  : std_logic;
  
  type RPEState is (idle,busy);
  signal rpe_state : RPEState;
begin  -- Behave

  reqR_fresh <= reqR and (not reqR_priority_encoded);
  there_is_a_fresh_request <= OrReduce(reqR_fresh);
  forward_enable <= reqR_priority_encoded;

  process(clk, rpe_state, there_is_a_fresh_request,ack_s)
	variable nstate: RPEState;
	variable latch_var : std_logic;
  begin
	nstate :=  rpe_state;
	latch_var := '0';
	req_s <= '0';
	if(rpe_state = idle) then
		if(there_is_a_fresh_request = '1') then
			latch_var := '1';
			nstate := busy;
		end if;
	elsif(rpe_state = busy) then
		req_s <= '1';
		if(ack_s = '1') then
			latch_var := '1';
			if(there_is_a_fresh_request = '1') then
				nstate := busy;
			else
				nstate := idle;
			end if;
		end if;
	end if;	

	if(clk'event and clk = '1') then
		if(reset = '1') then
			rpe_state <= idle;
			reqR_priority_encoded <= (others => '0');
		else
			if(latch_var = '1') then
				reqR_priority_encoded <= 
					PriorityEncode(reqR_fresh);
			end if;
			rpe_state <= nstate;
		end if;
	end if;

  end process;
  
  process(ack_s,reqR_priority_encoded)
  begin
    for I in reqR'range loop
      ackR(I) <= reqR_priority_encoded(I) and ack_s;
    end loop;  -- I
  end process;

  
end Behave;

architecture Fair of Request_Priority_Encode_Entity is
  signal reqR_register, reqR_priority_encoded : std_logic_vector(num_reqs-1 downto 0);
  signal reqR_reg_is_non_zero: std_logic;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

   SingleRequester: if num_reqs = 1 generate
	req_s <= reqR(0);
	ackR(0) <= ack_s;
	forward_enable <= reqR;
   end generate SingleRequester;

 
   MultipleRequesters: if num_reqs > 1 generate
   reqR_reg_is_non_zero <= OrReduce(reqR_register);
   req_s <= reqR_reg_is_non_zero;
   forward_enable <= reqR_priority_encoded;

   -- logic: in each cycle, reqR_register is updated
   --    1. if reqR_register is 0, then it is updated by reqR.
   --    2. if reqR_register is not-zero, then a forward request
   --         is enabled by a priority encode.  When this request
   --         is acked, the correspond reqR_register bit is set to 0.
   --

   process(clk, reset, reqR_reg_is_non_zero, reqR, reqR_register, ack_s, reqR_priority_encoded)
	variable next_reqR_register : std_logic_vector(num_reqs-1 downto 0);
   begin
	next_reqR_register := reqR_register;

        if(reqR_reg_is_non_zero = '0') then
	    next_reqR_register := reqR;
        elsif(ack_s = '1') then
	    next_reqR_register := reqR_register xor reqR_priority_encoded;

	    -- if next_reqR_register turns out to be 0, and if
	    -- there are waiting requests (other than the one that
	    -- was just acknowledge), then in principle, we could
	    -- fast track (reqR xor reqR_priority_encoded) into
            -- reqR_register...
	     if(OrReduce(next_reqR_register) = '0') then
            	 next_reqR_register := (reqR xor reqR_priority_encoded);
	     end if;
        end if;

        if(clk'event and clk = '1') then
		if(reset = '1') then
  			reqR_priority_encoded <= (others => '0');
			reqR_register <= (others => '0');
		else
			reqR_register <= next_reqR_register;
			reqR_priority_encoded <= PriorityEncode(next_reqR_register);
		end if;
	end if;
	
   end process;

  process(ack_s,reqR_priority_encoded)
  begin
    for I in reqR'range loop
      ackR(I) <= reqR_priority_encoded(I) and ack_s;
    end loop;  -- I
  end process;

  end generate MultipleRequesters;
end Fair;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- rL -> aL delay can be 0
entity Sample_Pulse_To_Level_Translate_Entity is
  generic (name: string);
  port( rL : in boolean;
        rR : out std_logic;
        aL : out boolean;
        aR : in std_logic;
        clk : in std_logic;
        reset : in std_logic);
end entity;

architecture Behave of Sample_Pulse_To_Level_Translate_Entity is
  type PullModeState is (Idle,Waiting);
  signal pull_mode_state : PullModeState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  process(clk, rL, aR, pull_mode_state)
    variable nstate : PullModeState;
  begin
    nstate := pull_mode_state;
    rR <= '0';
    aL <= false;

      case pull_mode_state is
        when Idle =>
          if(rL) then
            rR <= '1';
            if(aR = '1') then
              aL <= true;
            else
              nstate := Waiting;
            end if;
          end if;
        when Waiting =>
	  rR <= '1';
          if(aR = '1') then
            nstate := Idle;
	    aL <= true;
          end if;
        when others => null;
      end case;

    if(clk'event and clk = '1') then
	if reset = '1' then
		pull_mode_state <= Idle;
	else
      		pull_mode_state <= nstate;
	end if;
    end if;
  end process;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;

entity SelectBase is
  generic(name: string; data_width: integer; flow_through: boolean := false);
  port(x,y: in std_logic_vector(data_width-1 downto 0);
       sel: in std_logic_vector(0 downto 0);
       req: in boolean;
       z: out std_logic_vector(data_width-1 downto 0);
       ack: out boolean;
       clk,reset: in std_logic);
end SelectBase;


architecture arch of SelectBase is 
begin

  noFlowThrough: if (not flow_through) generate

    process(x,y,sel,req,reset,clk)
    begin
      
      if(clk'event and clk = '1') then
        if(reset = '1') then
          ack <= false;
          z <= (others => '0');
        elsif(sel(sel'right) = '1' and req = true) then
          ack <= req;
          z <= x;
        elsif(sel(sel'right) = '0' and req = true) then
          ack <= req;
          z <= y; 
        else 
          ack <= false;
        end if;
      end if;
    end process;
  end generate noFlowThrough;

  flowThrough: if flow_through generate
	ack <= req;
	z <= x when sel(sel'right) = '1' else y;
  end generate flowThrough;

end arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.Utilities.all;
use ahir.Subprograms.all;

-- a simple slicing element.
entity Slicebase is
  generic(name: string; in_data_width : integer; high_index: integer; low_index : integer; flow_through : boolean := false);
  port(din: in std_logic_vector(in_data_width-1 downto 0);
       dout: out std_logic_vector(high_index-low_index downto 0);
       req: in boolean;
       ack: out boolean;
       clk,reset: in std_logic);
end Slicebase;


architecture arch of Slicebase is

begin

  assert ((high_index < in_data_width) and (low_index >= 0) and (high_index >= low_index))
    report "inconsistent slice parameters" severity failure;
  
  flowThrough: if flow_through generate
    ack <= req;
    dout <= din(high_index downto low_index);
  end generate flowThrough;

  noFlowThrough: if not flow_through generate
    process(clk)
      variable ack_var  : boolean;
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          ack <= false;
        else
          ack <= req;
        end if;
      end if;
    end process;

    process(clk)
    begin
      if(clk'event and clk = '1') then
        if(req) then
          dout <= din(high_index downto low_index);
        end if;
      end if;
    end process;
  end generate noFlowThrough;
  
end arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity SplitCallArbiterNoInArgsNoOutArgs is
  generic(name: string;
	   num_reqs: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
end SplitCallArbiterNoInArgsNoOutArgs;


architecture Struct of SplitCallArbiterNoInArgsNoOutArgs is
   signal call_data   : std_logic_vector(num_reqs-1 downto 0); -- tie to 0
   signal call_mdata  : std_logic_vector(0 downto 0); -- ignore.

   signal return_data : std_logic_vector(num_reqs-1 downto 0); --ignore
   signal return_mdata : std_logic_vector(0 downto 0); -- tie to 0
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin
	call_data <= (others => '0');
	return_mdata <= (others => '0');

	baseArbiter:
		SplitCallArbiter
			generic map (name => name & "-base",
					num_reqs => num_reqs,
					call_data_width => 1, -- fake
					return_data_width => 1, --fake
					caller_tag_length => caller_tag_length,
					callee_tag_length => callee_tag_length
				    )
			port map (
					call_reqs => call_reqs,
					call_acks => call_acks,
					call_data => call_data,
					call_tag => call_tag,
					call_mreq => call_mreq,
					call_mack => call_mack,
					call_mdata => call_mdata,
					call_mtag => call_mtag,
					return_reqs => return_reqs,
					return_acks => return_acks,
					return_data => return_data,
					return_tag => return_tag,
					return_mreq => return_mreq,
					return_mack => return_mack,
					return_mdata => return_mdata,
					return_mtag => return_mtag,
					clk => clk, reset => reset			
				 );

end Struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity SplitCallArbiterNoInargs is
  generic(name: string;
	  num_reqs: integer;
	  return_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
end SplitCallArbiterNoInargs;


architecture Struct of SplitCallArbiterNoInargs is
   signal call_data   : std_logic_vector(num_reqs-1 downto 0); -- tie to 0
   signal call_mdata  : std_logic_vector(0 downto 0); -- ignore.
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin
	call_data <= (others => '0');
	
	baseArbiter:
		SplitCallArbiter
			generic map (name => name & "-base",
					num_reqs => num_reqs,
					call_data_width => 1, -- fake
					return_data_width => return_data_width,
					caller_tag_length => caller_tag_length,
					callee_tag_length => callee_tag_length
				    )
			port map (
					call_reqs => call_reqs,
					call_acks => call_acks,
					call_data => call_data,
					call_tag => call_tag,
					call_mreq => call_mreq,
					call_mack => call_mack,
					call_mdata => call_mdata,
					call_mtag => call_mtag,
					return_reqs => return_reqs,
					return_acks => return_acks,
					return_data => return_data,
					return_tag => return_tag,
					return_mreq => return_mreq,
					return_mack => return_mack,
					return_mdata => return_mdata,
					return_mtag => return_mtag,
					clk => clk, reset => reset			
				 );
end Struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity SplitCallArbiterNoOutArgs is
  generic(name: string;
	  num_reqs: integer;
	  call_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
end SplitCallArbiterNoOutArgs;


architecture Struct of SplitCallArbiterNoOutArgs is
    signal return_data : std_logic_vector(num_reqs-1 downto 0);
    signal return_mdata : std_logic_vector(0 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin
	return_mdata <= (others => '0');

	baseArbiter:
		SplitCallArbiter
			generic map (name => name & "-base",
					num_reqs => num_reqs,
					call_data_width => call_data_width,
					return_data_width => 1, -- fake
					caller_tag_length => caller_tag_length,
					callee_tag_length => callee_tag_length
				    )
			port map (
					call_reqs => call_reqs,
					call_acks => call_acks,
					call_data => call_data,
					call_tag => call_tag,
					call_mreq => call_mreq,
					call_mack => call_mack,
					call_mdata => call_mdata,
					call_mtag => call_mtag,
					return_reqs => return_reqs,
					return_acks => return_acks,
					return_data => return_data,
					return_tag => return_tag,
					return_mreq => return_mreq,
					return_mack => return_mack,
					return_mdata => return_mdata,
					return_mtag => return_mtag,
					clk => clk, reset => reset			
				 );
	
end Struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity SplitCallArbiter is
  generic(name: string;
	  num_reqs: integer;
	  call_data_width: integer;
	  return_data_width: integer;
	  caller_tag_length: integer;
          callee_tag_length: integer);
  port ( -- ready/ready handshake on all ports
    -- ports for the caller
    call_reqs   : in  std_logic_vector(num_reqs-1 downto 0);
    call_acks   : out std_logic_vector(num_reqs-1 downto 0);
    call_data   : in  std_logic_vector((num_reqs*call_data_width)-1 downto 0);
    call_tag    : in  std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- call port connected to the called module
    call_mreq   : out std_logic;
    call_mack   : in  std_logic;
    call_mdata  : out std_logic_vector(call_data_width-1 downto 0);
    call_mtag   : out std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    -- similarly for return, initiated by the caller
    return_reqs : in  std_logic_vector(num_reqs-1 downto 0);
    return_acks : out std_logic_vector(num_reqs-1 downto 0);
    return_data : out std_logic_vector((num_reqs*return_data_width)-1 downto 0);
    return_tag  : out std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
    -- return from function
    return_mreq : out std_logic;
    return_mack : in std_logic;
    return_mdata : in  std_logic_vector(return_data_width-1 downto 0);
    return_mtag : in  std_logic_vector(callee_tag_length+caller_tag_length-1 downto 0);
    clk: in std_logic;
    reset: in std_logic);
end SplitCallArbiter;


architecture Struct of SplitCallArbiter is
   signal pe_call_reqs, pe_call_reqs_reg: std_logic_vector(num_reqs-1 downto 0);
   signal return_acks_sig: std_logic_vector(num_reqs-1 downto 0);

   type TwordArray is array (natural range <>) of std_logic_vector(return_mdata'length-1 downto 0);
   signal return_data_sig : TwordArray(num_reqs-1 downto 0);

   type TagwordArray is array (natural range <>) of std_logic_vector(caller_tag_length-1 downto 0);
   signal return_tag_sig : TagwordArray(num_reqs-1 downto 0);

   type CallStateType is (idle, busy);
   signal call_state: CallStateType;


   signal latch_call_data : std_logic;
   signal call_mdata_prereg  : std_logic_vector(call_data_width-1 downto 0);
   signal callee_mtag_prereg, callee_mtag_reg  : std_logic_vector(callee_tag_length-1 downto 0);
   signal caller_mtag_reg  : std_logic_vector(caller_tag_length-1 downto 0);

   signal fair_call_reqs, fair_call_acks: std_logic_vector(num_reqs-1 downto 0);
   signal return_mreq_sig : std_logic_vector(num_reqs-1 downto 0); 

   constant ztag: std_logic_vector(callee_tag_length-1 downto 0) := (others => '0');

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

  --
  -- cut through when there is no contention.
  --
  singleRequester: if num_reqs = 1 generate

	call_mreq <= call_reqs(0);
	call_acks(0) <= call_mack;
	call_mdata <= call_data;
	call_mtag <= ztag & call_tag;

	return_mreq <= return_reqs(0);
	return_acks(0) <= return_mack;
	return_data <= return_mdata;
        return_tag <= return_mtag (caller_tag_length - 1 downto 0);

  end generate singleRequester;


 multipleRequesters: if num_reqs > 1 generate

  -----------------------------------------------------------------------------
  -- "fairify" the call-reqs.
  -----------------------------------------------------------------------------
  fairify: NobodyLeftBehind generic map (name => name & "-fairify", num_reqs => num_reqs)
		port map (clk => clk, reset => reset, reqIn => call_reqs, ackOut => call_acks,
					reqOut => fair_call_reqs, ackIn => fair_call_acks);

  -----------------------------------------------------------------------------
  -- priority encode incoming
  -----------------------------------------------------------------------------
   pe_call_reqs <= PriorityEncode(fair_call_reqs);

   ----------------------------------------------------------------------------
   -- process to handle call_reqs  --> call_mreq muxing
   ----------------------------------------------------------------------------
   process(clk,pe_call_reqs,call_state,call_mack,reset)
        variable nstate: CallStateType;
        variable there_is_a_call : std_logic;
   begin
	nstate := call_state;
        there_is_a_call := OrReduce(pe_call_reqs);
	latch_call_data <= '0';
	call_mreq <= '0';

	if(call_state = idle) then
		if(there_is_a_call = '1') then
			latch_call_data <=  '1';
			nstate := busy;
		end if;
	elsif (call_state = busy) then
		call_mreq <= '1';
		if(call_mack = '1') then
			if(there_is_a_call = '1') then
				latch_call_data <=  '1';
                        else
				nstate := idle;
			end if;
		end if;
	end if;
	
	if(clk'event and clk = '1') then
		if(reset = '1') then
			call_state <= idle;
			pe_call_reqs_reg <= (others => '0');
		else
			call_state <= nstate;
		end if;
	end if;
   end process;



   -- combinational process.. generate fair_call_acks, and also
   -- mux to input of call data register.
   process(pe_call_reqs,latch_call_data,call_data)
	variable out_data : std_logic_vector(call_data_width-1 downto 0);
   begin
	fair_call_acks <= (others => '0');
	out_data := (others => '0');
       	for I in num_reqs-1 downto 0 loop
       		if(pe_call_reqs(I) = '1') then
			out_data := call_data(((I+1)*call_data_width)-1 downto
							I*call_data_width);
       			-- Extract(call_data,I,out_data);
			if(latch_call_data = '1') then
				fair_call_acks(I) <= '1';
			end if;
       		end if;
	end loop;
	call_mdata_prereg <= out_data;
   end process;

   -- call data register.
   process(clk)
   begin
     if(clk'event and clk = '1') then
     	if(latch_call_data = '1') then
		call_mdata <= call_mdata_prereg;
		callee_mtag_reg <= callee_mtag_prereg;
        end if;  -- I
     end if;
   end process;
 

   -- tag generation.
   tagGen : BinaryEncoder generic map (name => name & "-tagGen", iwidth => num_reqs,
                                       owidth => callee_tag_length)
     port map (din => pe_call_reqs, dout => callee_mtag_prereg);

   -- on a successful call, register the tag from the caller
   -- side..
   process(clk, pe_call_reqs, call_tag, latch_call_data)
	variable tvar : std_logic_vector(caller_tag_length-1 downto 0);
   begin
	tvar := (others => '0');

	for T in 0 to num_reqs-1 loop
         if(pe_call_reqs(T) = '1') then
           tvar := call_tag(((T+1)*caller_tag_length)-1 downto T*caller_tag_length);
         end if;
        end loop;

       if(clk'event and clk = '1') then
	if(latch_call_data = '1') then
		caller_mtag_reg <= tvar;
	end if;
       end if;
   end process;     

   -- call tag.
   call_mtag <= callee_mtag_reg & caller_mtag_reg;


   ----------------------------------------------------------------------------
   -- reverse path
   ----------------------------------------------------------------------------
   -- pack registers into return data array
   process(return_data_sig)
     variable lreturn_data : std_logic_vector((num_reqs*return_data_width)-1 downto 0);
   begin
     for J in return_data_sig'high(1) downto return_data_sig'low(1) loop
       lreturn_data(((J+1)*return_data_width)-1 downto J*return_data_width)
		:= return_data_sig(J);
       -- Insert(lreturn_data,J,return_data_sig(J));
     end loop;  -- J
     return_data <= lreturn_data;
   end process;
 
   -- 2D to 1D packing.
   process(return_tag_sig)
     variable lreturn_tag : std_logic_vector((num_reqs*caller_tag_length)-1 downto 0);
   begin
     for J in return_tag_sig'high(1) downto return_tag_sig'low(1) loop
       lreturn_tag(((J+1)*caller_tag_length)-1 downto J*caller_tag_length)
		:= return_tag_sig(J);
       -- Insert(lreturn_tag,J,return_tag_sig(J));
     end loop;  -- J
     return_tag <= lreturn_tag;
   end process;

   -- always ready to accept return data!
   -- Sorry, this is broken..  What if successive returns
   -- arrive from a pipelined module aimed at the same destination?
   -- Back-pressure is needed!
   return_mreq <= OrReduce(return_mreq_sig);

   -- return to caller.
   return_acks <= return_acks_sig;
   
   -- incoming data written into appropriate register.
   RetGen: for I in num_reqs-1 downto 0 generate

     fsm: block
       signal ack_reg, valid_flag : std_logic;
       signal data_reg : std_logic_vector(return_mdata'length-1 downto 0);
       signal tag_reg  : std_logic_vector(caller_tag_length-1 downto 0);
       signal return_state : CallStateType;
     begin  -- block fsm

       -- valid = '1' implies this index is incoming
       valid_flag <= '1' when return_mack = '1' and (I = To_Integer(To_Unsigned(return_mtag(caller_tag_length+callee_tag_length-1 downto caller_tag_length)))) else '0';

       --------------------------------------------------------------------------
       -- ack FSM
       --------------------------------------------------------------------------
       process(clk,return_state,return_reqs(I),valid_flag,reset)
	variable nstate: CallStateType;
	variable latch_var: std_logic;
       begin

	 nstate := return_state;
	 latch_var := '0';
	 return_acks_sig(I) <= '0';

	 if(return_state = Idle) then
		if(valid_flag = '1') then
			latch_var := '1';
			nstate := Busy;
		end if;		
	 else 
		return_acks_sig(I) <= '1';
		if((valid_flag = '1') and (return_reqs(I) = '1')) then
			latch_var := '1';
		elsif (return_reqs(I) = '1') then
			nstate := Idle;
		end if;
	 end if;

	 return_mreq_sig(I) <= latch_var;

         if clk'event and clk= '1' then
           if(reset = '1') then
             return_state <= Idle;
	   else
	     return_state <= nstate;
	     if(latch_var = '1') then
             	data_reg <= return_mdata;
             	tag_reg  <= return_mtag(caller_tag_length-1 downto 0);
	     end if;
           end if;
         end if;
       end process;

       -- pass info out of the generate
       return_data_sig(I) <= data_reg;
       return_tag_sig(I)  <= tag_reg;

     end block fsm;
     
   end generate RetGen;

  end generate multipleRequesters;
end Struct;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.OperatorPackage.all;
use ahir.FloatOperatorPackage.all;
use ahir.BaseComponents.all;

entity SplitOperatorBase is
  generic
    (
      name: string;
      operator_id   : string := "ApIntAdd";          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer := 4;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer := 0;    -- width of input2
      num_inputs    : integer := 1;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer := 4;          -- width of output.
      constant_operand : std_logic_vector := "0001"; -- constant operand.. (it is always the second operand)
      constant_width: integer := 4;
      twidth        : integer := 1;          -- tag width
      use_constant  : boolean := true
      );
  port (
    -- req/ack follow level protocol
    reqR: out std_logic;
    ackR: in std_logic;
    reqL: in std_logic;
    ackL : out  std_logic;
    -- tagL is passed out to tagR
    tagL       : in  std_logic_vector(twidth-1 downto 0);
    -- input array consists of m sets of 1 or 2 possibly concatenated
    -- operands.
    dataL      : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
    dataR      : out std_logic_vector(owidth-1 downto 0);
    -- tagR is received from tagL, concurrent
    -- with dataR
    tagR       : out std_logic_vector(twidth-1 downto 0);
    clk, reset : in  std_logic);
end SplitOperatorBase;


architecture Vanilla of SplitOperatorBase is
  signal   result    : std_logic_vector(owidth-1 downto 0);
  signal   state_sig : std_logic;
  constant tag0      : std_logic_vector(tagR'length-1 downto 0) := (others => '0');
  constant iwidth : integer := iwidth_1  + iwidth_2;

begin  -- Behave

  assert((num_inputs = 1) or (num_inputs = 2)) report "either 1 or 2 inputs" severity failure;

  f2f: if (operator_id = "ApFloatResize") generate
	f2f_inst: GenericFloatToFloat
			generic map (
					name => name & "-f2f_inst",
					tag_width => twidth,
					in_exponent_width => input1_characteristic_width,
					in_fraction_width => input1_mantissa_width,
					out_exponent_width => output_characteristic_width,
					out_fraction_width => output_mantissa_width)
			port map (
					INF => dataL, 
					OUTF => dataR,
					clk => clk, reset => reset,
					env_rdy => reqL, accept_rdy => ackR,
					tag_in => tagL, tag_out => tagR,
					f2fi_rdy => ackL, f2fo_rdy => reqR		
				);
  end generate f2f;


  Not_f2f:  if(operator_id /= "ApFloatResize") generate
    reqR <= reqL;
    ackL <= ackR;
    tagR <= tagL;
    
    comb_block: GenericCombinationalOperator
      generic map (
	name => name & "-comb_block",
        operator_id                 => operator_id,
        input1_is_int               => input1_is_int,
        input1_characteristic_width => input1_characteristic_width,
        input1_mantissa_width       => input1_mantissa_width,
        iwidth_1                    => iwidth_1,
        input2_is_int               => input2_is_int,
        input2_characteristic_width => input2_characteristic_width,
        input2_mantissa_width       => input2_mantissa_width,
        iwidth_2                    => iwidth_2,
        num_inputs                  => num_inputs,
        output_is_int               => output_is_int,
        output_characteristic_width => output_characteristic_width,
        output_mantissa_width       => output_mantissa_width,
        owidth                      => owidth,
        constant_operand            => constant_operand,
        constant_width		  => constant_width,
        use_constant                => use_constant)
      port map (
        data_in => dataL,
        result  => dataR);
  end generate Not_f2f;
  
  
end Vanilla;
  
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity SplitOperatorShared is
    generic
    (
      name : string;
      operator_id   : string := "ApIntAdd";          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer := 4;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer := 0;    -- width of input2
      num_inputs    : integer := 1;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer := 4;          -- width of output.
      constant_operand : std_logic_vector := "0001"; -- constant operand.. (it is always the second operand)
      constant_width: integer := 4;
      use_constant  : boolean := true;
      no_arbitration: boolean := false;
      min_clock_period: boolean := true;
      num_reqs : integer := 3; -- how many requesters?
      detailed_buffering_per_output : IntegerArray := (0 => 0);
      detailed_buffering_per_input : IntegerArray  := (0 => 0);
      use_input_buffering: boolean := false;
      full_rate : boolean 
    );
  port (
    -- req/ack follow level protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackR                     : out BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    reqR                     : in  BooleanArray(num_reqs-1 downto 0);
    -- input data consists of concatenated pairs of ips
    dataL                    : in std_logic_vector(((iwidth_1 + iwidth_2)*num_reqs)-1 downto 0);
    -- output data consists of concatenated pairs of ops.
    dataR                    : out std_logic_vector((owidth*num_reqs)-1 downto 0);
    -- with dataR
    clk, reset              : in std_logic);
end SplitOperatorShared;

architecture Vanilla of SplitOperatorShared is

  constant num_operands : integer := num_inputs;
  constant iwidth : integer := iwidth_1 + iwidth_2;
  
  constant ignore_tag  : boolean := no_arbitration or (reqL'length = 1);

  signal idata : std_logic_vector(iwidth-1 downto 0);
  signal odata: std_logic_vector(owidth-1 downto 0);

  constant tag_length: integer := Maximum(1,Ceil_Log2(reqL'length));
  signal itag,otag : std_logic_vector(tag_length-1 downto 0);
  signal ireq,iack, oreq, oack: std_logic;

  constant debug_flag : boolean := global_debug_flag;
  
begin  -- Behave
  assert ackL'length = reqL'length report "mismatched req/ack vectors" severity error;
  

  -- DebugGen: if debug_flag generate 
    -- assert( (not ((reset = '0') and (clk'event and clk = '1') and no_arbitration)) or Is_At_Most_One_Hot(reqL))
    -- report "in no-arbitration case, at most one request should be hot on clock edge (in SplitOperatorShared)" severity error;
  -- end generate DebugGen;
  
   imuxWithInputBuf: InputMuxWithBuffering
      generic map(name => name & "-imux " , 
		iwidth => iwidth*num_reqs,
                owidth => iwidth, 
                twidth => tag_length,
                nreqs => num_reqs,
		buffering => detailed_buffering_per_input,
		full_rate => full_rate, 
                no_arbitration => no_arbitration,
                registered_output => false)
      port map(
        reqL       => reqL,
        ackL       => ackL,
        reqR       => ireq,
        ackR       => iack,
        dataL      => dataL,
        dataR      => idata,
        tagR       => itag,
        clk        => clk,
        reset      => reset);

  op: SplitOperatorBase
    generic map (
      name => name & "-op",
      operator_id   => operator_id,
      input1_is_int => input1_is_int,
      input1_characteristic_width => input1_characteristic_width,
      input1_mantissa_width => input1_mantissa_width,
      iwidth_1  => iwidth_1,
      input2_is_int => input2_is_int,
      input2_characteristic_width => input2_characteristic_width,
      input2_mantissa_width  => input2_mantissa_width,
      iwidth_2  => iwidth_2,
      num_inputs  => num_inputs,
      output_is_int => output_is_int,
      output_characteristic_width => output_characteristic_width,
      output_mantissa_width  => output_mantissa_width,
      owidth    => owidth,
      constant_operand => constant_operand,
      constant_width => constant_width,
      twidth     => tag_length,
      use_constant => use_constant
      )
    port map (
      reqL => ireq,
      ackL => iack,
      reqR => oreq,
      ackR => oack,
      dataL => idata,
      dataR => odata,
      tagR => otag,
      tagL => itag,
      clk => clk,
      reset => reset);


  odemux: OutputDeMuxBaseWithBuffering
    generic map (
        name => name & "-odemux ",
  	iwidth => owidth,
  	owidth =>  owidth*num_reqs,
	twidth =>  tag_length,
	nreqs  => num_reqs,
        detailed_buffering_per_output => detailed_buffering_per_output,
	full_rate => full_rate )  
    port map (
      reqL   => oreq,
      ackL   => oack,
      dataL => odata,
      tagL  => otag,
      reqR  => reqR,
      ackR  => ackR,
      dataR => dataR,
      clk   => clk,
      reset => reset);
  
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity StoreCompleteShared is
  generic (name : string; num_reqs: integer := 3;
	   tag_length: integer :=  3;
	    detailed_buffering_per_output: IntegerArray);
  port (
    -- in requester array, pulse protocol
    -- more than one requester can be active
    -- at any time
    reqR : in BooleanArray(num_reqs-1 downto 0);
    -- out ack array, pulse protocol
    -- more than one ack can be sent back
    -- at any time.
    --
    -- Note: req -> ack delay can be 0
    ackR : out BooleanArray(num_reqs-1 downto 0);
    -- mreq goes out to memory as 
    -- a response to mack.
    mreq : out std_logic;
    mack : in  std_logic;
    -- mtag to distinguish the 
    -- requesters.
    mtag : in std_logic_vector(tag_length-1 downto 0);
    -- rising edge of clock is used
    clk : in std_logic;
    -- synchronous reset, active high
    reset : in std_logic);
end StoreCompleteShared;

architecture Behave of StoreCompleteShared is
begin  -- Behave


  odemux: OutputDemuxBaseNoData
    generic map (
      name => name & "-odemux",
      twidth =>  tag_length,
      nreqs  => num_reqs,
      detailed_buffering_per_output => detailed_buffering_per_output)
    port map (
      reqL   => mack,                   -- cross-over (mack from mem-subsystem)
      ackL   => mreq,                   -- cross-over 
      tagL  =>  mtag,
      reqR  => reqR,
      ackR  => ackR,
      clk   => clk,
      reset => reset);

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity StoreReqShared is
    generic
    (
	name: string;
	addr_width: integer;
	data_width : integer;
	time_stamp_width : integer;
      	num_reqs : integer; -- how many requesters?
	tag_length: integer;
	no_arbitration: Boolean := false;
        min_clock_period: Boolean := true        
    );
  port (
    -- req/ack follow pulse protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    -- address corresponding to access
    addr                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
    data                    : in std_logic_vector((data_width*num_reqs)-1 downto 0);
    -- address to memory
    maddr                   : out std_logic_vector(addr_width-1 downto 0);
    mdata                   : out std_logic_vector(data_width-1 downto 0);
    mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);
    mreq                    : out std_logic;
    mack                    : in std_logic;
    -- clock, reset (active high)
    clk, reset              : in std_logic);
end StoreReqShared;

architecture Vanilla of StoreReqShared is

  constant iwidth: integer := addr_width*num_reqs;
  constant owidth: integer := addr_width;

  signal idata: std_logic_vector(((addr_width+data_width)*num_reqs)-1 downto 0);
  signal odata: std_logic_vector((addr_width+data_width)-1 downto 0);

  constant debug_flag : boolean := global_debug_flag;
--  constant registered_output: boolean := min_clock_period and (time_stamp_width = 0);

  -- must register..  ack implies that address has been sampled.
  constant registered_output: boolean := true;

  
  signal imux_tag_out: std_logic_vector(tag_length-1 downto 0);
begin  -- Behave

  TstampGen: if time_stamp_width > 0 generate

    Tstamp: block
	signal time_stamp: std_logic_vector(time_stamp_width-1 downto 0);
    begin 
  	mtag <= imux_tag_out & time_stamp;

	-- ripple counter.
	process(clk)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				time_stamp <= (others => '0');
			else
				for I in 1 to time_stamp_width-1 loop
					time_stamp(I) <= time_stamp(I) xor AndReduce(time_stamp(I-1 downto 0));
				end loop;
				time_stamp(0) <= not time_stamp(0);
			end if;
		end if;
	end process;
    end block;
    
  end generate TstampGen;

  NoTstampGen: if time_stamp_width < 1 generate
	mtag <= imux_tag_out;
  end generate NoTstampGen;

  process(addr,data)
  begin
     for I in num_reqs-1 downto 0 loop
	idata(((I+1)*(addr_width+data_width))-1 downto (I*(addr_width+data_width))) <= 
		addr(((I+1)*addr_width)-1 downto I*addr_width) & 
		data(((I+1)*data_width)-1 downto I*data_width);
     end loop;
  end process;

  maddr <= odata(addr_width+data_width-1 downto data_width);
  mdata <= odata(data_width-1 downto 0);

  assert(tag_length >= Ceil_Log2(num_reqs)) report "insufficient tag width" severity error;

  -- debugCase: if debug_flag generate
    -- assert( (not ((reset = '0') and (clk'event and clk = '1') and no_arbitration)) or Is_At_Most_One_Hot(reqL))
      -- report "in no-arbitration case, at most one request should be hot on clock edge (in SplitOperatorShared)" severity error;
  -- end generate debugCase;
  
  imux: InputMuxBase
  	generic map(name => name & "-imux",
		    iwidth => (addr_width+data_width)*num_reqs ,
                    owidth => addr_width+data_width, 
                    twidth => tag_length,
                    nreqs => num_reqs,
                    registered_output => registered_output,
                    no_arbitration => no_arbitration)
    port map(
      reqL       => reqL,
      ackL       => ackL,
      reqR       => mreq,
      ackR       => mack,
      dataL      => idata,
      dataR      => odata,
      tagR       => imux_tag_out,
      clk        => clk,
      reset      => reset);
  
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity SynchFifoWithDPRAM is
  generic(name: string; queue_depth: integer := 3; data_width: integer := 72);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack : out std_logic;
       nearly_full: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity SynchFifoWithDPRAM;

architecture behave of SynchFifoWithDPRAM is

  constant addr_width_of_dpram: integer := Ceil_Log2(queue_depth);
  signal read_pointer, write_pointer : unsigned(addr_width_of_dpram-1 downto 0);
  signal queue_size : integer range 0 to queue_depth;

  function Incr(x: unsigned; M: integer) return unsigned is
     variable ret_var: unsigned(1 to x'length);
  begin
    if(x < M) then
      	ret_var := (x + 1);
    else
	ret_var := (others => '0');
    end if;
    return(ret_var);
  end Incr;

  signal incr_read_pointer, incr_write_pointer : unsigned(addr_width_of_dpram-1 downto 0);

  signal write_to_dpram, read_from_dpram, latch_read_data: std_logic;
  
  type ReadFsmState is (Idle, Valid, WaitPop);
  signal read_state: ReadFsmState;
  signal read_data : std_logic_vector(data_width-1 downto 0);
  signal read_data_reg: std_logic_vector(data_width-1 downto 0);

  signal ready_for_bypass: std_logic;
-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- SimModel


  assert(queue_depth > 1) report "Synch FIFO depth must be greater than 1" severity failure;
  assert (queue_size < queue_depth) report "Queue " & name & " is full." severity note;

  incr_read_pointer <= Incr(read_pointer, queue_depth-1);
  incr_write_pointer <= Incr(write_pointer, queue_depth-1);

  -- pointer management process.
  process(clk, reset)
  begin
     if(clk'event and (clk = '1') ) then
	if(reset ='1') then
		read_pointer <= (others => '0');
		write_pointer <= (others => '0');
                queue_size <= 0;
	else
             if(write_to_dpram = '1') then
		write_pointer <= incr_write_pointer;
	     end if;
	     if (read_from_dpram = '1') then
		read_pointer <= incr_read_pointer;
	     end if;

	     if ((write_to_dpram = '1') and (read_from_dpram = '0')) then
		queue_size <= queue_size + 1;
	     elsif ((read_from_dpram = '1') and (write_to_dpram = '0')) then
		queue_size <= queue_size - 1;
	     end if;
	end if;
     end if;
  end process;

  -- write is easy.
  write_to_dpram <= '1' when ((push_req = '1') and (queue_size < queue_depth) and (ready_for_bypass = '0')) 
						else '0';
  push_ack <= '1' when (queue_size < queue_depth) else '0';
  nearly_full <= '1' when (queue_size = (queue_depth-1)) else '0';


  
  -- read process.
  process(clk,reset,read_state, pop_req, queue_size, push_req) 
	variable next_read_state:  ReadFsmState;
	variable read_from_dpram_var: std_logic;
	variable latch_read_data_var: std_logic;
	variable ready_for_bypass_var: std_logic;
	variable pop_ack_var : std_logic;
  begin
	next_read_state := read_state;
	read_from_dpram_var := '0';
	latch_read_data_var := '0';
	ready_for_bypass_var := '0';

	pop_ack_var := '0';
	
	
	case read_state is 
		when Idle =>
			if (queue_size > 0) then
				read_from_dpram_var := '1';
				next_read_state := Valid;	
			elsif (push_req = '1') then
				ready_for_bypass_var := '1';
				latch_read_data_var := '1';
				next_read_state := WaitPop;
			end if;
		when Valid =>
			pop_ack_var := '1';
			if (pop_req = '1') then
				if(queue_size > 0) then 
					read_from_dpram_var := '1';
				elsif (push_req = '1') then
					ready_for_bypass_var := '1';
					latch_read_data_var := '1';
					next_read_state := WaitPop;
				else
					next_read_state := Idle;
				end if;
			else
				next_read_state := WaitPop;
				latch_read_data_var := '1';
			end if;
		when WaitPop =>
			pop_ack_var := '1';
			if(pop_req = '1') then
				if(queue_size > 0) then
					read_from_dpram_var := '1';
					next_read_state := Valid;
				elsif (push_req = '1') then
					ready_for_bypass_var := '1';
					latch_read_data_var := '1';
					next_read_state := WaitPop;
				else
					next_read_state := Idle;
				end if;
			end if;
	end case;

	read_from_dpram <= read_from_dpram_var;
	latch_read_data <= latch_read_data_var;
	ready_for_bypass <= ready_for_bypass_var;

	pop_ack <= pop_ack_var;

	if(clk'event and (clk = '1')) then
		if(reset = '1') then
			read_state <= Idle;
		else
			read_state <= next_read_state;
		end if;
	end if;
  end process;

  rf_1w_1r_inst: register_file_1w_1r_port
		generic map (name => name & "-register_file_1w_1r", 
				g_addr_width => addr_width_of_dpram,
				g_data_width => data_width)
		port map (
				-- port 0 for write
				datain_0 =>  data_in,
				addrin_0 =>  std_logic_vector(write_pointer),
				enable_0 => write_to_dpram,
				-- port 1 for read.
				dataout_1 => read_data,
				addrin_1 =>  std_logic_vector(read_pointer),
				enable_1 => read_from_dpram,
				-- clock pos edge..
				clk => clk, 
				-- reset active high.
				reset => reset
			 );
   -- registering
   process(clk, reset)
   begin
       if(clk'event and (clk = '1')) then
		if(reset = '1') then
			read_data_reg <= (others => '0');
		elsif (latch_read_data = '1') then
			if(ready_for_bypass = '1') then
				read_data_reg <= data_in;
			else
				read_data_reg <= read_data;
			end if;
		end if;
       end if;
   end process;

   -- output mux
   data_out <= read_data when (read_state = Valid) else read_data_reg;

end behave;


------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- written by Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;

entity SynchLifo is
  generic(name : string; queue_depth: integer := 3; data_width: integer := 72);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack : out std_logic;
       nearly_full: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity SynchLifo;

architecture behave of SynchLifo is

  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);

  signal queue_array : QueueArray(queue_depth-1 downto 0);
  signal tos_pointer, write_pointer : integer range 0 to queue_depth-1;
  signal queue_size : integer range 0 to queue_depth;

  signal bypass_reg, mem_out_reg : std_logic_vector(data_width-1 downto 0);

  function Incr(x: integer; M: integer) return integer is
  begin
    if(x < M) then
      return(x + 1);
    else
      return(0);
    end if;
  end Incr;

  signal nearly_empty_sig, empty_sig, full_sig : std_logic;
  signal select_bypass : std_logic;
  signal pop_req_int: std_logic;
begin  -- SimModel
  assert (queue_size < queue_depth) report "LIFO " & name & " is full." severity note;

  full_sig  <= '1' when (queue_size = queue_depth) else '0';
  empty_sig <= '1' when (queue_size = 0) else '0';
  nearly_empty_sig <= '1' when (queue_size = 1) else '0';
  nearly_full <= '1' when (queue_size = (queue_depth-1)) else '0';


  -- single process
  process(clk,reset,
          empty_sig,
          full_sig,
          queue_size,
          push_req,
          pop_req, pop_req_int,
          tos_pointer,
          write_pointer)
    variable qsize : integer range 0 to queue_depth;
    variable push,pop,bypass : boolean;
    variable next_tos_ptr, next_write_ptr : integer range 0 to queue_depth-1;
  begin
    qsize := queue_size;
    push  := false;
    pop   := false;
    next_tos_ptr := tos_pointer;
    next_write_ptr := write_pointer;
    
    if((queue_size < queue_depth) and push_req = '1') then
      push := true;
    end if;

    if((queue_size > 0) and pop_req_int = '1') then
      pop := true;
    end if;

    bypass := push and pop;
    
    if push and (not pop) then
      -- increment write pointer and tos-pointer.
      next_write_ptr := Incr(write_pointer,queue_depth-1);
      if(queue_size > 0) then
        next_tos_ptr := Incr(tos_pointer,queue_depth-1);
      else
        next_tos_ptr := 0;
      end if;
      qsize := queue_size + 1;      
    elsif pop and (not push) then
      if(write_pointer > 0) then
      	next_write_ptr := write_pointer-1;
      else
	-- if write-ptr is 0, it must have wrapped around
        -- in the increment function.
	next_write_ptr := queue_depth - 1;
      end if;

      if(tos_pointer > 0) then
        next_tos_ptr := tos_pointer - 1;
      else
        next_tos_ptr := 0;
      end if;
      qsize := queue_size - 1;            
    end if;
    
    if(clk'event and clk = '1') then
      
      if(reset = '1') then
	queue_size <= 0;
        tos_pointer <= 0;
        write_pointer <= 0;
        select_bypass <= '0';
      else
        queue_size <= qsize;
        tos_pointer <= next_tos_ptr;
        write_pointer <= next_write_ptr;
      end if;

      if(bypass) then
        select_bypass <= '1';
        bypass_reg <= data_in;
      elsif push then
        queue_array(write_pointer) <= data_in;
        select_bypass <= '1';
        bypass_reg <= data_in;
      elsif pop then
        select_bypass <= '0';        
	if(tos_pointer > 0) then
        	mem_out_reg <= queue_array(tos_pointer-1);        
	end if;
      end if;
    end if;  
  end process;

  push_ack <= not full_sig;
  pop_ack  <= not empty_sig;
  pop_req_int <= pop_req;
  data_out <= bypass_reg when select_bypass = '1' else mem_out_reg;
  
end behave;


------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- a simple register
entity SynchResetRegisterSlv is
  generic(name: string; data_width: integer);
  port(din: in std_logic_vector(data_width-1 downto 0);
       dout: out std_logic_vector(data_width-1 downto 0);
       clk,reset: in std_logic);
end SynchResetRegisterSlv;


architecture Simplest of SynchResetRegisterSlv is
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

  process(din,reset,clk)
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          dout <= (others => '0');
        else
          dout <= din;
 	end if;
      end if;
  end process;

end architecture Simplest;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- a simple register
entity SynchResetRegisterUnsigned is
  generic(name: string; data_width: integer);
  port(din: in unsigned(data_width-1 downto 0);
       dout: out unsigned(data_width-1 downto 0);
       clk,reset: in std_logic);
end SynchResetRegisterUnsigned;


architecture Simplest of SynchResetRegisterUnsigned is
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

  process(din,reset,clk)
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          dout <= (others => '0');
        else
          dout <= din;
 	end if;
      end if;
  end process;

end architecture Simplest;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity SynchToAsynchReadInterface is
  generic (
    name: string;
    data_width : integer);
  port (
    clk : in std_logic;
    reset  : in std_logic;
    synch_req : in std_logic;  -- indicates that synch side has data.
    synch_ack : out std_logic; -- indicates that synch-side should do a read 
				-- (there is a 1-cycle delay between the assertion of this signal
				--   and availability of synch data).
    asynch_req : out std_logic; --  indicates that asynch side wishes to forward data
    asynch_ack: in std_logic;  -- indicates that forwarded data is accepte.
    synch_data: in std_logic_vector(data_width-1 downto 0); -- synch data in
    asynch_data : out std_logic_vector(data_width-1 downto 0)); -- forwarded data out.
end SynchToAsynchReadInterface;


architecture Behave of SynchToAsynchReadInterface is

  type InMatchingFSMState is (Idle,LatchSynchData,WaitForAsynchAck);
  signal in_fsm_state : InMatchingFSMState;

  signal synch_data_reg: std_logic_vector(data_width-1 downto 0);
  
begin

  process(clk,reset, in_fsm_state, synch_req, asynch_ack)
    variable next_state: InMatchingFSMState;
    variable synch_ack_var, asynch_req_var: std_logic;
    variable latch_var: std_logic;
    
  begin
    next_state := in_fsm_state;

    synch_ack_var := '0';
    asynch_req_var := '0';
    latch_var := '0';
    
    case in_fsm_state is
      when idle =>
        if(synch_req = '1') then
            synch_ack_var := '1';
	    next_state := LatchSynchData;
	end if;
      when LatchSynchData =>
	-- latch the data from the synch side
        -- because that data is guarateed to be valid
        -- only in this cycle.
        latch_var := '1';
        asynch_req_var := '1';
        if(asynch_ack = '1') then
          synch_ack_var := '1';
	  -- if synch-req is '1', then stay
          -- here... 
          if(synch_req = '0') then
          	next_state :=  Idle;
	  end if;
        else
           next_state := WaitForAsynchAck;
        end if;
      when WaitForAsynchAck =>
	-- wait for ack from asynch-side
        asynch_req_var := '1';
        if(asynch_ack = '1')  then
            -- if synch-requests then latch
            -- synch data.
	    if(synch_req = '1') then
               synch_ack_var := '1';
               next_state := LatchSynchData;
            else
               next_state := Idle;
            end if;
        end if;
      when others => null;
    end case;
    
    synch_ack <= synch_ack_var;
    asynch_req <= asynch_req_var;

    if(clk'event and clk = '1') then
       if(reset = '1') then
         in_fsm_state <= Idle;
         synch_data_reg <= (others => '0');
       else 
         in_fsm_state <= next_state;
	 if(latch_var = '1') then
		synch_data_reg <= synch_data;
	 end if;
       end if;
    end if;
  end process;

  asynch_data <= synch_data when (in_fsm_state = LatchSynchData) else synch_data_reg; 
  
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

--
-- The deep version of the unload buffer.
--   When a synch-fifo is used, the in->out latency is two cycles.
--   To avoid this, we use a pass-around from in->out when the queue
--   is empty.
--
entity UnloadBufferDeep is
  generic (name: string; buffer_size: integer ; data_width : integer ; nonblocking_read_flag : boolean := false);
  port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data : out std_logic;
        clk : in std_logic;
        reset: in std_logic);
end UnloadBufferDeep;

architecture default_arch of UnloadBufferDeep is

  signal pop_req, pop_ack, push_req, push_ack: std_logic_vector(0 downto 0);
  signal pipe_data_out, data_to_unload_register:  std_logic_vector(data_width-1 downto 0);

  signal number_of_elements_in_pipe: unsigned ((Ceil_Log2(buffer_size+2))-1 downto 0); 
  signal pipe_has_data: boolean;

  signal unload_register_ready: boolean;

  signal pop_req_from_unload_register : std_logic;
  signal pop_ack_to_unload_register   : std_logic;

  signal write_to_pipe: boolean;
  signal unload_from_pipe : boolean;

begin  -- default_arch

  assert (buffer_size > 1) report "UnloadBufferDeep must have queue-size > 1" severity failure;


		-- count number of elements in pipe.
  process(clk, reset)
  begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			number_of_elements_in_pipe <= (others => '0');
		else
			if((pop_req(0) = '1') and (pop_ack(0) = '1')) then
				if(not ((push_req(0) = '1') and (push_ack(0) = '1'))) then
					number_of_elements_in_pipe <= (number_of_elements_in_pipe -1);
				end if;
			elsif((push_req(0) = '1') and (push_ack(0) = '1')) then
				number_of_elements_in_pipe <= (number_of_elements_in_pipe + 1);
			end if;
		end if;
	end if;
  end process;
	
  has_data <= '1' when pipe_has_data else '0';
  pipe_has_data <= (number_of_elements_in_pipe > 0);
  write_to_pipe <= (pipe_has_data or (not unload_register_ready));
  unload_from_pipe <= pipe_has_data;

  unload_register_ready <= (pop_req_from_unload_register = '1');
 
  -- if pipe does not have data, then we will be bypassing write-data straight
  -- to the unload-register, if it is ready to accept stuff.
  push_req(0) <= write_req when write_to_pipe else '0';
  write_ack   <= push_ack(0);

  pop_ack_to_unload_register <= pop_ack(0) when unload_from_pipe else write_req;
  pop_req(0)  <= pop_req_from_unload_register;
  data_to_unload_register <= pipe_data_out when unload_from_pipe else write_data;

  -- the input pipe.
  bufPipe : PipeBase generic map (
        	name =>  name & "-blocking_read-bufPipe",
        	num_reads  => 1,
        	num_writes => 1,
        	data_width => data_width,
        	lifo_mode  => false,
		shift_register_mode => false,
        	depth      => buffer_size,
		save_slot  => false,
		full_rate  => false)
      	port map (
        	read_req   => pop_req,
        	read_ack   => pop_ack,
        	read_data  => pipe_data_out,
        	write_req  => push_req,
        	write_ack  => push_ack,
        	write_data => write_data,
        	clk        => clk,
        	reset      => reset);

   ulReg: UnloadRegister 
			generic map (name => name & "-unload-register",
					data_width => data_width,
						bypass_flag => false,
						   nonblocking_read_flag => nonblocking_read_flag)
			port map (
					write_data => data_to_unload_register,
					write_req => pop_ack_to_unload_register,
					write_ack => pop_req_from_unload_register,
					unload_req => unload_req,
					unload_ack => unload_ack,
					read_data => read_data,
					clk => clk,  reset => reset
				);
							

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

--
-- An optimized version of the unload buffer, to be used when the buffer_size is > 1.
--     Uses a standard queue followed by a state machine..
--
entity UnloadBufferOptimized is
  generic (name: string; buffer_size: integer ; data_width : integer; 
		bypass_flag: boolean; nonblocking_read_flag : boolean := false);
  port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data : out std_logic;
        clk : in std_logic;
        reset: in std_logic);
end UnloadBufferOptimized;

architecture default_arch of UnloadBufferOptimized is

  signal pop_req, pop_ack : std_logic;
  signal unload_ack_sig: boolean; 
  signal empty, full: std_logic;

   type FsmState is (sA, sB, sC, sD);
   signal fsm_state: FsmState;

   signal queue_data_out: std_logic_vector(data_width-1 downto 0);

begin  -- default_arch

  assert (buffer_size /= 1) report "UnloadBufferOptimized must have queue-size != 1" severity failure;

  has_data <= not empty;

  qinst: QueueBaseWithEmptyFull
		generic map (name => name & ":qinst",
				queue_depth => buffer_size,
				data_width => data_width,
				reverse_bypass_flag => bypass_flag
			    )
		port map (
				empty => empty,
				full  => full,
				push_req => write_req,
				push_ack => write_ack,
				pop_req => pop_req,
				pop_ack => pop_ack,
				data_in => write_data,
				data_out => queue_data_out,
				clk => clk,
				reset => reset);	

	-- FSM
        process(clk, reset, pop_ack, fsm_state, unload_req, queue_data_out)
		variable next_fsm_state_var:  FsmState;
		variable unload_ack_var: boolean;
		variable pop_req_var: std_logic;
   		variable read_data_var: std_logic_vector(data_width-1 downto 0);
	begin
		next_fsm_state_var := fsm_state;
		unload_ack_var := false;
		pop_req_var := '0';
		read_data_var := queue_data_out;

		case fsm_state is
			when sA =>
				-- In the beginning, nothing has
				-- been read from the queue.
				if unload_req then
					next_fsm_state_var := sB;
				end if;
			when sB =>
				--
				-- Ack if queue has data 
				--
				-- Careful about the non-blocking
				-- behaviour.
				if (pop_ack = '1') then		     -- p
					unload_ack_var := true;
					if unload_req then
						-- pop from the queue
						-- since the next-req
						-- has arrived.
						pop_req_var := '1';
					else
						next_fsm_state_var := sC;
					end if;
				elsif nonblocking_read_flag then -- (~p).n
					-- non-blocking... as if pop_ack is
					-- asserted except that read data 
					-- will be zero-ed out.
					read_data_var := (others => '0');

					-- ack the zero data..
					unload_ack_var := true;

					if unload_req then
						-- do not pop here
						-- The queue data has not 
						-- been used yet.
						next_fsm_state_var := sB;
					else
						-- wait for update req
						-- but ensure that read_data
						-- is zero-ed out.
						next_fsm_state_var := sD;
					end if;
				end if;
			when sC =>
				--
				-- you will come to this state only
				-- if pop_ack = '1'... you are waiting
				-- for an update-req to start the
				-- next cycle.
				if unload_req then
					-- pop only when signaled by
					-- unload_req
					pop_req_var := '1';

					-- go to sB before reacting
					-- to the update-req.
					next_fsm_state_var := sB;
				end if;

			when SD =>
				--
				-- you got here because pop_ack was false
				-- and non-block was true.  zero out the
				-- read_data until the next unload_req.
				-- 
				-- you are waiting for an update-req to
				-- start the next cycle.
				--
				-- Keep read_data_var = 0 here.  you
				-- do not want the changed queue output
				-- to sneak to the user.
				--
				read_data_var := (others => '0');
				if unload_req then
					--
					-- do not pop!  
					-- 
					-- go to sB before reacting
					-- to the update-req.
					next_fsm_state_var := sB;
				end if;
		end case;

		pop_req <= pop_req_var;
		unload_ack <= unload_ack_var;
		read_data <= read_data_var;

		if(clk'event and (clk = '1')) then
			if (reset = '1') then
				fsm_state <= sA;
			else
				fsm_state <= next_fsm_state_var;
			end if;
		end if;
	end process;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;
-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

--
-- The unload buffer is used all over the place.  We will use
-- three forms
--     depth <= 1
--         fast cut through with buffering provided by a single register
--     depth >= 2
--         queue + wastes a buffer.  this needs to be sorted out.
--
--  Using shallow buffers (<= 1) will result in fast in->out 
--  performance but combinational through paths.  Using deeper
--  buffers will result in at least one unit of delay from in->out
--
-- Added Nov 2019.  Added use_unload_register generic.
--
--   This avoids wastage of an extra register in the unload-buffer.
--   but must be used with a cut-through that has a combinational
--   unload_ack to write_ack path.
-- 
entity UnloadBuffer is
  generic (name: string; buffer_size: integer ; data_width : integer ; 
			-- bypass = true means there are some combi paths.
			--   from write_req to unload_ack
			--   from unload_req to write_ack
			--   from write_data to read_data.
			bypass_flag : boolean := false; 
			-- self-explanatory.
			nonblocking_read_flag : boolean := false;
			-- if false use new revised version of the unload buffer (revised)
			-- which does not need an unload-register.
			use_unload_register: boolean := true);
  port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);
end UnloadBuffer;

architecture default_arch of UnloadBuffer is

  signal pop_req, pop_ack, push_req, push_ack: std_logic_vector(0 downto 0);
  signal pipe_data_out, data_to_unload_register:  std_logic_vector(data_width-1 downto 0);

  signal pipe_has_data: boolean;

  signal unload_register_ready: boolean;

  signal pop_req_from_unload_register : std_logic;
  signal pop_ack_to_unload_register   : std_logic;

  signal write_to_pipe: boolean;
  signal unload_from_pipe : boolean;

  signal empty, full: std_logic;
  --
  -- try to save a slot if buffer size is 1... this
  -- tries to prevent a 100% wastage of resources
  -- and allows us to use 2-depth buffers to cut long
  -- combinational paths.
  --
  function DecrDepth (buf_size: integer; bypass: boolean)
	return integer is
      variable ret_val: integer;
  begin
      ret_val := buf_size;
      if((not bypass) and (buffer_size = 1)) then
	ret_val := buf_size - 1;
      end if;
      return ret_val;
  end function DecrDepth;

  constant actual_buffer_size  : integer  := DecrDepth (buffer_size, bypass_flag);

  constant bypass_flag_to_ureg : boolean := (bypass_flag or (buffer_size = 0));

  constant shallow_flag : boolean :=    (buffer_size < global_pipe_shallowness_threshold);

  constant revised_case_blocking: boolean := 
		((buffer_size > 0) 
			and (bypass_flag or (buffer_size > 1))
                        and shallow_flag 
			and (not use_unload_register) 
			and (not nonblocking_read_flag));

  constant revised_case_non_blocking: boolean := 
		global_use_optimized_unload_buffer and
			((buffer_size > 1) and (not bypass_flag) and
				 shallow_flag and  nonblocking_read_flag);


  constant un_revised_case: boolean :=  (not revised_case_blocking) and 
						(not revised_case_non_blocking) and
							shallow_flag;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch

  RevisedCaseBlocking: if revised_case_blocking generate

         assert false report "ULB REVISED BLOCKING  " & name & ":" & Convert_To_String(data_width*buffer_size) 
			severity note;

	ulb_revised: UnloadBufferRevised
			generic map (name => name & "-revised",
					buffer_size => buffer_size, data_width => data_width,
						bypass_flag => bypass_flag)
			port map (
				write_req => write_req,
				write_ack => write_ack,
				unload_req => unload_req,
				unload_ack => unload_ack,
				write_data => write_data,
				read_data => read_data, 
				has_data => has_data,
				clk => clk, reset => reset);
  end generate RevisedCaseBlocking;

  RevisedCaseNonblocking: if revised_case_non_blocking generate

         assert false report "ULB REVISED NONBLOCKING  " & name & ":" & Convert_To_String(data_width*buffer_size) 
			severity note;

	ulb_revised: UnloadBufferRevisedNonblocking
			generic map (name => name & "-revised",
					buffer_size => buffer_size, data_width => data_width,
						bypass_flag => bypass_flag)
			port map (
				write_req => write_req,
				write_ack => write_ack,
				unload_req => unload_req,
				unload_ack => unload_ack,
				write_data => write_data,
				read_data => read_data, 
				has_data => has_data,
				clk => clk, reset => reset);
  end generate RevisedCaseNonblocking;

  DeepCase: if not shallow_flag generate
         assert false report "ULB DEEP " & name & ":" & Convert_To_String(data_width*buffer_size) 
			severity note;

	ulb_deep: UnloadBufferDeep
			generic map (name => name & "-deep",
					buffer_size => buffer_size, data_width => data_width,
						nonblocking_read_flag => nonblocking_read_flag)
			port map (
				write_req => write_req,
				write_ack => write_ack,
				unload_req => unload_req,
				unload_ack => unload_ack,
				write_data => write_data,
				read_data => read_data, 
				has_data => has_data,
				clk => clk, reset => reset);
  end generate DeepCase;

  NotRevisedCase: if un_revised_case generate

    ShallowCase: if shallow_flag  generate
      assert false report "ULB with ULREG " & name & ":" & Convert_To_String(data_width*buffer_size) 
			severity note;

      bufGt0: if actual_buffer_size > 0 generate

  	has_data <= '1' when pipe_has_data else '0';

  	pipe_has_data <= (empty = '0');
	write_to_pipe <= (pipe_has_data or (not unload_register_ready));
	unload_from_pipe <= pipe_has_data;

	unload_register_ready <= (pop_req_from_unload_register = '1');
 
	-- if pipe does not have data, then we will be bypassing write-data straight
	-- to the unload-register, if it is ready to accept stuff.
	push_req(0) <= write_req when write_to_pipe else '0';
	write_ack   <= push_ack(0);

	pop_ack_to_unload_register <= pop_ack(0) when unload_from_pipe else write_req;
	pop_req(0)  <= pop_req_from_unload_register;
	data_to_unload_register <= pipe_data_out when unload_from_pipe else write_data;

  	-- the input pipe.
  	bufPipe : QueueBaseWithEmptyFull generic map (
        	name =>  name & "-blocking_read-bufPipe",
        	data_width => data_width,
        	queue_depth      => actual_buffer_size)
      	port map (
        	pop_req   => pop_req(0),
        	pop_ack   => pop_ack(0),
        	data_out  => pipe_data_out,
        	push_req  => push_req(0),
        	push_ack  => push_ack(0),
        	data_in => write_data,
		empty => empty,
		full => full,
        	clk        => clk,
        	reset      => reset);

     end generate bufGt0;
	

     -- unload-register will provide bypassed buffering.
     bufEq0: if (actual_buffer_size = 0) generate

	empty <= '1';
	full  <= '0';

	has_data <= '0';

	data_to_unload_register <= write_data;
	pop_ack_to_unload_register <= write_req;
	write_ack  <= pop_req_from_unload_register;
     end generate bufEq0;

     ulReg: UnloadRegister 
			generic map (name => name & "-unload-register",
					data_width => data_width,
						bypass_flag => bypass_flag_to_ureg,
						   nonblocking_read_flag => nonblocking_read_flag)
			port map (
					write_data => data_to_unload_register,
					write_req => pop_ack_to_unload_register,
					write_ack => pop_req_from_unload_register,
					unload_req => unload_req,
					unload_ack => unload_ack,
					read_data => read_data,
					clk => clk,  reset => reset
				);
							
   end generate ShallowCase;
 end generate NotRevisedCase;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- The unshared operator uses a split protocol.
--    reqL/ackL  for sampling the inputs
--    reqR/ackR  for updating the outputs.
-- The two pairs should be used independently,
-- that is, there should be NO DEPENDENCY between
-- ackL and reqR!
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.OperatorPackage.all;
use ahir.BaseComponents.all;
use ahir.FloatOperatorPackage.all;

entity UnsharedOperatorBase is
  generic
    (
      name: string;
      operator_id   : string;          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer;    -- width of input2
      num_inputs    : integer := 2;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer;          -- width of output.
      constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
      constant_width : integer;
      use_constant  : boolean := false
      );
  port (
    -- req -> ack follow pulse protocol
    reqL:  in Boolean;
    ackL : out Boolean;
    reqR : in Boolean;
    ackR:  out Boolean;
    -- operands.
    dataL      : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
    dataR      : out std_logic_vector(owidth-1 downto 0);
    clk, reset : in  std_logic);
end UnsharedOperatorBase;


architecture Vanilla of UnsharedOperatorBase is
  signal   result: std_logic_vector(owidth-1 downto 0);
  constant iwidth : integer := iwidth_1  + iwidth_2;
  
  -- joined req, and joint ack.
  signal fReq,fAck: boolean;
 

begin  -- Behave


  assert((num_inputs = 1) or (num_inputs = 2)) report "either 1 or 2 inputs" severity failure;

  -----------------------------------------------------------------------------
  -- join the two reqs..
  -----------------------------------------------------------------------------
  rJ: join2 generic map (name => operator_id & "-join2", bypass => true)
		port map(pred0 => reqL, pred1 => reqR, symbol_out => fReq, clk => clk, reset => reset);

  
  dE: control_delay_element generic map(name => name & "-dE", delay_value  => 1)
		port map(req => fReq, ack => fAck, clk => clk, reset => reset);
  
  -- same ack to both.
  ackL <= fAck;
  ackR <= fAck;

  -----------------------------------------------------------------------------
  -- combinational block..
  -----------------------------------------------------------------------------
  comb_block: GenericCombinationalOperator
    generic map (
      name => name & "-comb_block", 
      operator_id                 => operator_id,
      input1_is_int               => input1_is_int,
      input1_characteristic_width => input1_characteristic_width,
      input1_mantissa_width       => input1_mantissa_width,
      iwidth_1                    => iwidth_1,
      input2_is_int               => input2_is_int,
      input2_characteristic_width => input2_characteristic_width,
      input2_mantissa_width       => input2_mantissa_width,
      iwidth_2                    => iwidth_2,
      num_inputs                  => num_inputs,
      output_is_int               => output_is_int,
      output_characteristic_width => output_characteristic_width,
      output_mantissa_width       => output_mantissa_width,
      owidth                      => owidth,
      constant_operand            => constant_operand,
      constant_width              => constant_width,
      use_constant                => use_constant)
    port map (data_in => dataL, result  => result);


  -----------------------------------------------------------------------------
  -- sample the output
  -----------------------------------------------------------------------------
  process(clk,reset)
  begin
    if(clk'event and clk = '1') then
      if(fReq) then
        dataR <= result;
      end if;
    end if;
  end process;
    
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Authors: Abhishek R. Kamath & Prashant Singhal
-- An IEEE-754 compliant Double-Precision pipelined multiplier
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity DoublePrecisionMultiplier is
  generic (name: string; tag_width : integer);
  port(
    INA, INB: in std_logic_vector(63 downto 0);   
    OUTM: out std_logic_vector(63 downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    NaN, oflow, uflow: out std_logic := '0';
    env_rdy, accept_rdy: in std_logic;
    muli_rdy, mulo_rdy: out std_logic);
end entity;

architecture rtl of DoublePrecisionMultiplier is

  type parpro is array (0 to 52) of std_logic_vector(52 downto 0);

  signal rdy1,rdy2,rdy3,rdy4,rdy5,rdy6,rdy7,rdy8,rdy9,rdy10,rdy11,rdy12: std_logic := '0';
  signal flag3,flag4,flag5,flag6,flag7,flag8,flag9,flag10,flag11: std_logic_vector(1 downto 0);
  signal fman11: std_logic_vector(51 downto 0);
  signal tag1,tag2,tag3,tag4,tag5,tag6,tag7,tag8,tag9,tag10,tag11: std_logic_vector(tag_width-1 downto 0);
  signal pipeline_stall: std_logic := '0';

  signal aman_1,aman_2,bman_1,bman_2: std_logic_vector(52 downto 0);
  signal anan1,bnan1,azero1,bzero1,ainf1,binf1,osgn1: std_logic := '0'; 
  signal aexp_s1,bexp_s1: std_logic_vector(10 downto 0);

  signal nocalc2,nocalc3,nocalc4,nocalc5,nocalc6,nocalc7,nocalc8,nocalc9,nocalc10,nocalc11: std_logic;-- := '0';
  signal output_s2,output_s23,output_s24,output_s25,output_s26,output_s27,output_s28,output_s29,output_s210,output_s211: std_logic_vector(2 downto 0);
  signal int_exp: std_logic_vector(11 downto 0);

  signal fexp3,fexp4,fexp5,fexp6,fexp7,fexp8,fexp9,fexp10,fexp11: std_logic_vector(10 downto 0);-- := X"00";

  signal pp: parpro;
  signal tr_400,tr_401,tr_402,tr_403,tr_404,tr_405,tr_406,tr_407,tr_408,tr_409,tr_410,tr_411,tr_412: std_logic_vector(105 downto 0);
  signal tr_413,tr_414,tr_415,tr_416,tr_417,tr_418,tr_419,tr_420,tr_421,tr_422,tr_423,tr_424,tr_425,tr_426: std_logic_vector(105 downto 0);

  signal tr501,tr502,tr503,tr504,tr505,tr506,tr507,tr508,tr509,tr510,tr511,tr512,tr513,tr514: std_logic_vector(105 downto 0);
  signal tr61,tr62,tr63,tr64,tr65,tr66,tr67: std_logic_vector(105 downto 0);
  signal tr71,tr72,tr73,tr74,tr71_int1,tr72_int1,tr71_int2: std_logic_vector(105 downto 0);


  signal tr401,tr402,tr403,tr404,tr405,tr406,tr407,tr408,tr409,tr410,tr411,tr412: std_logic_vector(105 downto 0);-- := X"000000000000";
  signal tr413,tr414,tr415,tr416,tr417,tr418,tr419,tr420,tr421,tr422,tr423,tr424: std_logic_vector(105 downto 0);-- := X"000000000000";
  signal tr425,tr426,tr427,tr428,tr429,tr430,tr431,tr432,tr433,tr434,tr435,tr436: std_logic_vector(105 downto 0);-- := X"000000000000";
  signal tr437,tr438,tr439,tr440,tr441,tr442,tr443,tr444,tr445,tr446,tr447,tr448: std_logic_vector(105 downto 0);-- := X"000000000000";
  signal tr449,tr450,tr451,tr452,tr453: std_logic_vector(105 downto 0);-- := X"000000000000";

begin

  stage_1: process(clk,reset)

    variable asgn,bsgn,osgn: std_logic := '0';
    variable aexp,bexp: std_logic_vector(10 downto 0);-- := "000" & X"00";
    variable aman,bman: std_logic_vector(52 downto 0);-- := "000000000000000000000000";
    variable anan,bnan,azero,bzero,ainf,binf: std_logic;-- := '0';

  begin
    if reset = '1' then
      rdy1 <= '0';
    else
      if clk'event and clk='1'then
        if env_rdy = '1' and pipeline_stall = '0' then
          --asgn1 <= INA(63);
          --bsgn1 <= INB(63);
          --aexp1 <= INA(62 downto 52);
          --bexp1 <= INB(62 downto 52);
          --aman1 <= '1' & INA(51 downto 0);
          --bman1 <= '1' & INB(51 downto 0);
          --rdy1 <= '1';
          

          --asgn := INA(63);
          --bsgn := INB(63);
          --osgn := INA(63) xor INB(63);

          
          aexp := INA(62 downto 52);
          bexp := INB(62 downto 52);
          aman := '1' & INA(51 downto 0);
          bman := '1' & INB(51 downto 0);
          
          
          
          if(aexp="111" & X"FF") then
            if(unsigned(aman)=0) then
              ainf := '1';
              anan := '0';
              azero := '0';
            else
              anan := '1';
              azero := '0';
              ainf := '0';
            end if;
          elsif(aexp="000"&X"00") then
            if unsigned(aman)=0 then
              azero := '1';
              ainf := '0';
              anan := '0';
            end if;
          else
            ainf := '0';
            anan := '0';
            azero := '0';
          end if;
          
          if(bexp="111"& X"FF") then
            if(unsigned(bman)=0) then
              binf := '1';
              bnan := '0';
              bzero := '0';
            else
              bnan := '1';
              bzero := '0';
              binf := '0';
            end if;
          elsif(bexp="000" & X"00") then
            if unsigned(bman)=0 then
              bzero := '1';
              binf := '0';
              bnan := '0';
            end if;
          else
            binf := '0';
            bnan := '0';
            bzero := '0';
          end if;

          osgn1 <= INA(63) xor INB(63);
          
          ainf1 <= ainf;
          binf1 <= binf;
          anan1 <= anan;
          bnan1 <= bnan;
          azero1 <= azero;
          bzero1 <= bzero;
          
          aexp_s1 <= aexp;
          bexp_s1 <= bexp;
          aman_1 <= aman;
          bman_1 <= bman;


          rdy1 <= '1';
          tag1 <= tag_in;
          
        elsif pipeline_stall = '1' then
        elsif env_rdy = '0' then
          rdy1 <= '0';
        end if;
      end if;
    end if;
  end process stage_1;





  stage_2: process(clk,reset)
  begin
    if reset = '1' then
      rdy2 <= '0';
    else
      if clk'event and clk='1'then
        if rdy1 = '1' and pipeline_stall = '0' then
          if (anan1 = '1' or bnan1 = '1') then
            output_s2 <= osgn1 & "10";
            nocalc2 <= '1';
          elsif (azero1 = '1' and binf1 = '1') or (ainf1 = '1' and bzero1 = '1') then
            output_s2 <= osgn1 & "10";
            nocalc2 <= '1';
          elsif azero1 = '1' or bzero1 = '1' then
            output_s2 <= osgn1 & "00";
            nocalc2 <= '1';
          elsif ainf1 = '1' or binf1 = '1' then
            output_s2 <= osgn1 & "11";
            nocalc2 <= '1';
          else
            int_exp <= std_logic_vector(unsigned('0' & aexp_s1) + unsigned('0' & bexp_s1));
            output_s2 <= osgn1 & "01";
            nocalc2 <= '0';
          end if;
          --aexp_s3 <= aexp_s2;
          --bexp_s3 <= bexp_s2;
          aman_2 <= aman_1;
          bman_2 <= bman_1;
          rdy2 <= '1';
          tag2 <= tag1;
          
          
        elsif pipeline_stall = '1' then
        elsif rdy1 = '0' then
          rdy2 <= '0';
        end if;
      end if;
    end if;
  end process stage_2;




  stage_3: process(clk,reset)

    variable exp3: unsigned(11 downto 0);

  begin
    if reset = '1' then
      rdy3 <= '0';
    else
      if clk'event and clk='1'then
        if rdy2 = '1' and pipeline_stall = '0' then
          if nocalc2 = '1' then
            nocalc3 <= '1';
            output_s23 <= output_s2;
            flag3 <= "00";
          elsif nocalc2 = '0' then
            exp3 := unsigned(int_exp);
            if(exp3 > 3069) then
              output_s23 <= output_s2(2) & "11";
              nocalc3 <= '1';
              flag3 <= "10";
            elsif(exp3 < 1023) then
              output_s23 <= output_s2(2) & "00";
              nocalc3 <= '1';
              flag3 <= "01";
            else
              exp3 := exp3 - 1023;
              output_s23 <= output_s2(2) & "01";
              nocalc3 <= '0';
              flag3 <= "00";
            end if;	
          end if;
          --aman_3 <= aman_2;
          --bman_3 <= bman_2;
          fexp3 <= std_logic_vector(exp3(10 downto 0));
          rdy3 <= '1';
          tag3 <= tag2;

          for i in 0 to 52 loop
            for j in 0 to 52 loop
              pp(i)(j) <= aman_2(j) and bman_2(i);
            end loop;
          end loop;

        elsif pipeline_stall = '1' then
        elsif rdy2 = '0' then
          rdy3 <= '0';
        end if;
      end if;
    end if;
  end process stage_3;





  stage_4: process(clk,reset)
  begin
    if reset = '1' then
      rdy4 <= '0';
    else
      if clk'event and clk='1'then
        if rdy3 = '1' and pipeline_stall = '0' then
          if nocalc3 = '1' then
            nocalc4 <= '1';
          elsif nocalc3 = '0' then
            
            tr401 <= X"0000000000000" & '0' & pp(0);
            tr402 <= X"0000000000000" & pp(1) & '0';
            tr403 <= X"000000000000" & "000" & pp(2) & "00";
            tr404 <= X"000000000000" & "00" & pp(3) & "000";	

            tr405 <= X"000000000000" & '0' & pp(4) & X"0";
            tr406 <= X"000000000000" & pp(5) & X"0" & '0';
            tr407 <= X"00000000000" & "000" & pp(6) & X"0" & "00";
            tr408 <= X"00000000000" & "00" & pp(7) & X"0" & "000";

            tr409 <= X"00000000000" & '0' & pp(8) & X"00";
            tr410 <= X"00000000000" & pp(9) & X"00" & '0';
            tr411 <= X"0000000000" & "000" & pp(10) & X"00" & "00";
            tr412 <= X"0000000000" & "00" & pp(11) & X"00" & "000";

            tr413 <= X"0000000000" & '0' & pp(12) & X"000";
            tr414 <= X"0000000000" & pp(13) & X"000" & '0';
            tr415 <= X"000000000" & "000" & pp(14) & X"000" & "00";
            tr416 <= X"000000000" & "00" & pp(15) & X"000" & "000";

            tr417 <= X"000000000" & '0' & pp(16) & X"0000";
            tr418 <= X"000000000" & pp(17) & X"0000" & '0';
            tr419 <= X"00000000" & "000" & pp(18) & X"0000" & "00";
            tr420 <= X"00000000" & "00" & pp(19) & X"0000" & "000";

            tr421 <= X"00000000" & '0' & pp(20) & X"00000";
            tr422 <= X"00000000" & pp(21) & X"00000" & '0';
            tr423 <= X"0000000" & "000" & pp(22) & X"00000" & "00";
            tr424 <= X"0000000" & "00" & pp(23) & X"00000" & "000";

            tr425 <= X"0000000" & '0' & pp(24) & X"000000";
            tr426 <= X"0000000" & pp(25) & X"000000" & '0';
            tr427 <= X"000000" & "000" & pp(26) & X"000000" & "00";
            tr428 <= X"000000" & "00" & pp(27) & X"000000" & "000";

            tr429 <= X"000000" & '0' & pp(28) & X"0000000";
            tr430 <= X"000000" & pp(29) & X"0000000" & '0';
            tr431 <= X"00000" & "000" & pp(30) & X"0000000" & "00";
            tr432 <= X"00000" & "00" & pp(31) & X"0000000" & "000";

            tr433 <= X"00000" & '0' & pp(32) & X"00000000";
            tr434 <= X"00000" & pp(33) & X"00000000" & '0';
            tr435 <= X"0000" & "000" & pp(34) & X"00000000" & "00";
            tr436 <= X"0000" & "00" & pp(35) & X"00000000" & "000";

            tr437 <= X"0000" & '0' & pp(36) & X"000000000";
            tr438 <= X"0000" & pp(37) & X"000000000" & '0';
            tr439 <= X"000" & "000" & pp(38) & X"000000000" & "00";
            tr440 <= X"000" & "00" & pp(39) & X"000000000" & "000";

            tr441 <= X"000" & '0' & pp(40) & X"0000000000";
            tr442 <= X"000" & pp(41) & X"0000000000" & '0';
            tr443 <= X"00" & "000" & pp(42) & X"0000000000" & "00";
            tr444 <= X"00" & "00" & pp(43) & X"0000000000" & "000";

            tr445 <= X"00" & '0' & pp(44) & X"00000000000";
            tr446 <= X"00" & pp(45) & X"00000000000" & '0';
            tr447 <= X"0" & "000" & pp(46) & X"00000000000" & "00";
            tr448 <= X"0" & "00" & pp(47) & X"00000000000" & "000";

            tr449 <= X"0" & '0' & pp(48) & X"000000000000";
            tr450 <= X"0" & pp(49) & X"000000000000" & '0';
            tr451 <= "000" & pp(50) & X"000000000000" & "00";
            tr452 <= "00" & pp(51) & X"000000000000" & "000";

            tr453 <= '0' & pp(52) & X"0000000000000";

            nocalc4 <= '0';
            
          end if;

          
          output_s24 <= output_s23;
          fexp4 <= fexp3;
          flag4 <= flag3;
          rdy4 <= '1';
          tag4 <= tag3;
          
        elsif pipeline_stall = '1' then
        elsif rdy3 = '0' then
          rdy4 <= '0';
        end if;
      end if;
    end if;
  end process stage_4;


  stage_5: process(clk,reset)
  begin
    if reset = '1' then
      rdy5 <= '0';
    else
      if clk'event and clk='1'then
        if rdy4 = '1' and pipeline_stall = '0' then
          if nocalc4 = '1' then
            nocalc5 <= '1';
          elsif nocalc4 = '0' then
            
            tr_400 <= std_logic_vector(unsigned(tr401) + unsigned(tr402));
            tr_401 <= std_logic_vector(unsigned(tr403) + unsigned(tr404));
            tr_402 <= std_logic_vector(unsigned(tr405) + unsigned(tr406));
            tr_403 <= std_logic_vector(unsigned(tr407) + unsigned(tr408));
            tr_404 <= std_logic_vector(unsigned(tr409) + unsigned(tr410));
            tr_405 <= std_logic_vector(unsigned(tr411) + unsigned(tr412));
            tr_406 <= std_logic_vector(unsigned(tr413) + unsigned(tr414));
            tr_407 <= std_logic_vector(unsigned(tr415) + unsigned(tr416));
            tr_408 <= std_logic_vector(unsigned(tr417) + unsigned(tr418));
            tr_409 <= std_logic_vector(unsigned(tr419) + unsigned(tr420));
            tr_410 <= std_logic_vector(unsigned(tr421) + unsigned(tr422));
            tr_411 <= std_logic_vector(unsigned(tr423) + unsigned(tr424));

            tr_412 <= std_logic_vector(unsigned(tr425) + unsigned(tr426));
            tr_413 <= std_logic_vector(unsigned(tr427) + unsigned(tr428));
            tr_414 <= std_logic_vector(unsigned(tr429) + unsigned(tr430));
            tr_415 <= std_logic_vector(unsigned(tr431) + unsigned(tr432));
            tr_416 <= std_logic_vector(unsigned(tr433) + unsigned(tr434));
            tr_417 <= std_logic_vector(unsigned(tr435) + unsigned(tr436));
            tr_418 <= std_logic_vector(unsigned(tr437) + unsigned(tr438));
            tr_419 <= std_logic_vector(unsigned(tr439) + unsigned(tr440));
            tr_420 <= std_logic_vector(unsigned(tr441) + unsigned(tr442));
            tr_421 <= std_logic_vector(unsigned(tr443) + unsigned(tr444));
            tr_422 <= std_logic_vector(unsigned(tr445) + unsigned(tr446));
            tr_423 <= std_logic_vector(unsigned(tr447) + unsigned(tr448));

            tr_424 <= std_logic_vector(unsigned(tr449) + unsigned(tr450));
            tr_425 <= std_logic_vector(unsigned(tr451) + unsigned(tr452));
            tr_426 <= tr453;

            nocalc5 <= '0';
            
          end if;

          
          output_s25 <= output_s24;
          fexp5 <= fexp4;
          flag5 <= flag4;
          rdy5 <= '1';
          tag5 <= tag4;
          
        elsif pipeline_stall = '1' then
        elsif rdy4 = '0' then
          rdy5 <= '0';
        end if;
      end if;
    end if;
  end process stage_5;



  stage_6: process(clk,reset)
  begin
    if reset = '1' then
      rdy6 <= '0';
    else
      if clk'event and clk='1'then
        if rdy5 = '1' and pipeline_stall = '0' then
          if nocalc5 = '1' then
            nocalc6 <= '1';
          else
            tr501 <= std_logic_vector(unsigned(tr_400) + unsigned(tr_401));
            tr502 <= std_logic_vector(unsigned(tr_402) + unsigned(tr_403));
            tr503 <= std_logic_vector(unsigned(tr_404) + unsigned(tr_405));
            tr504 <= std_logic_vector(unsigned(tr_406) + unsigned(tr_407));
            tr505 <= std_logic_vector(unsigned(tr_408) + unsigned(tr_409));
            tr506 <= std_logic_vector(unsigned(tr_410) + unsigned(tr_411));

            tr507 <= std_logic_vector(unsigned(tr_412) + unsigned(tr_413));
            tr508 <= std_logic_vector(unsigned(tr_414) + unsigned(tr_415));
            tr509 <= std_logic_vector(unsigned(tr_416) + unsigned(tr_417));
            tr510 <= std_logic_vector(unsigned(tr_418) + unsigned(tr_419));
            tr511 <= std_logic_vector(unsigned(tr_420) + unsigned(tr_421));
            tr512 <= std_logic_vector(unsigned(tr_422) + unsigned(tr_423));

            tr513 <= std_logic_vector(unsigned(tr_424) + unsigned(tr_425));
            tr514 <= tr_426;
            
            nocalc6 <= '0';
          end if;

          output_s26 <= output_s25;
          fexp6 <= fexp5;
          flag6 <= flag5;
          rdy6 <= '1';
          tag6 <= tag5;
          
        elsif pipeline_stall = '1' then
        elsif rdy5 = '0' then
          rdy6 <= '0';
        end if;
      end if;
    end if;
  end process stage_6;



  stage_7: process(clk,reset)
  begin
    if reset = '1' then
      rdy7 <= '0';
    else
      if clk'event and clk='1'then
        if rdy6 = '1' and pipeline_stall = '0' then
          if nocalc6 = '1' then
            nocalc7 <= '1';
          else
            tr61 <= std_logic_vector(unsigned(tr501) + unsigned(tr502));
            tr62 <= std_logic_vector(unsigned(tr503) + unsigned(tr504));
            tr63 <= std_logic_vector(unsigned(tr505) + unsigned(tr506));

            tr64 <= std_logic_vector(unsigned(tr507) + unsigned(tr508));
            tr65 <= std_logic_vector(unsigned(tr509) + unsigned(tr510));
            tr66 <= std_logic_vector(unsigned(tr511) + unsigned(tr512));

            tr67 <= std_logic_vector(unsigned(tr513) + unsigned(tr514));
            
            
            nocalc7 <= '0';
          end if;

          output_s27 <= output_s26;
          fexp7 <= fexp6;
          flag7 <= flag6;
          rdy7 <= '1';
          tag7 <= tag6;
          
        elsif pipeline_stall = '1' then
        elsif rdy6 = '0' then
          rdy7 <= '0';
        end if;
      end if;
    end if;
  end process stage_7;

  stage_8: process(clk,reset)
  begin
    if reset = '1' then
      rdy8 <= '0';
    else
      if clk'event and clk='1'then
        if rdy7 = '1' and pipeline_stall = '0' then
          if nocalc7 = '1' then
            nocalc8 <= '1';
          else
            tr71 <= std_logic_vector(unsigned(tr61) + unsigned(tr62));
            tr72 <= std_logic_vector(unsigned(tr63) + unsigned(tr64));
            tr73 <= std_logic_vector(unsigned(tr65) + unsigned(tr66));
            tr74 <= tr67;
            
            nocalc8 <= '0';
          end if;
          
          output_s28 <= output_s27;
          fexp8 <= fexp7;
          flag8 <= flag7;
          rdy8 <= '1';
          tag8 <= tag7;
          
        elsif pipeline_stall = '1' then
        elsif rdy7 = '0' then
          rdy8 <= '0';
        end if;
      end if;
    end if;
  end process stage_8;

  stage_9: process(clk,reset)
  begin
    if reset = '1' then
      rdy9 <= '0';
    else
      if clk'event and clk='1'then
        if rdy8 = '1' and pipeline_stall = '0' then
          if nocalc8 = '1' then
            nocalc9 <= '1';
          else
            tr71_int1 <= std_logic_vector(unsigned(tr71) + unsigned(tr72));
            tr72_int1 <= std_logic_vector(unsigned(tr73) + unsigned(tr74));
            nocalc9 <= '0';
          end if;
          
          output_s29 <= output_s28;
          fexp9 <= fexp8;
          flag9 <= flag8;
          rdy9 <= '1';
          tag9 <= tag8;
          
        elsif pipeline_stall = '1' then
        elsif rdy8 = '0' then
          rdy9 <= '0';
        end if;
      end if;
    end if;
  end process stage_9;


  stage_10: process(clk,reset)
  begin
    if reset = '1' then
      rdy10 <= '0';
    else
      if clk'event and clk='1'then
        if rdy9 = '1' and pipeline_stall = '0' then
          if nocalc9 = '1' then
            nocalc10 <= '1';
          else
            tr71_int2 <= std_logic_vector(unsigned(tr71_int1) + unsigned(tr72_int1));
            nocalc10 <= '0';
          end if;
          
          output_s210 <= output_s29;
          fexp10 <= fexp9;
          flag10 <= flag9;
          rdy10 <= '1';
          tag10 <= tag9;
          
        elsif pipeline_stall = '1' then
        elsif rdy9 = '0' then
          rdy10 <= '0';
        end if;
      end if;
    end if;
  end process stage_10;



  stage_11: process(clk,reset)
    variable man8: std_logic_vector(53 downto 0);
    variable exp8: unsigned(10 downto 0);
  begin
    if reset = '1' then
      rdy11 <= '0';
    else
      if clk'event and clk='1'then
        if rdy10 = '1' and pipeline_stall = '0' then
          if nocalc10 = '1' then
            nocalc11 <= '1';
            output_s211 <= output_s210;
            flag11 <= flag10;
          elsif nocalc10 = '0' then
            man8 := tr71_int2(105 downto 52);
            exp8 := unsigned(fexp10);
            if man8(53) = '1' then
              if	exp8 = 2046 then
                output_s211 <= output_s210(2) & "11";
                nocalc11 <= '1';
                flag11 <= "10";
              else
                exp8 := exp8 + 1;
                nocalc11 <= '0';
                fman11 <= man8(52 downto 1);
                output_s211 <= output_s210;
                flag11 <= flag10;
              end if;
            elsif exp8 = 0 then
              output_s211 <= output_s210(2) & "00";
              nocalc11 <= '1';
              flag11 <= "01";
            else
              fman11 <= man8(51 downto 0);
              output_s211 <= output_s210;
              nocalc11 <= '0';
              flag11 <= flag10;
            end if;
          end if;		
          rdy11 <= '1';
          tag11 <= tag10;
          fexp11 <= std_logic_vector(exp8);
        elsif pipeline_stall = '1' then
        elsif rdy10 = '0' then
          rdy11 <= '0';
        end if;
      end if;
    end if;
  end process stage_11;


  stage_12: process(clk,reset)
    variable temp: std_logic_vector(2 downto 0);
  begin
    if reset = '1' then
      rdy12 <= '0';
    else
      if clk'event and clk='1'then
        if rdy11 = '1' and pipeline_stall = '0' then
          rdy12 <= '1';
          temp := output_s211;
          if nocalc11 = '1' then
            case(temp(1 downto 0)) is
              when("00") => OUTM <= temp(2) & "000" & X"000000000000000"; NaN <= '0'; oflow <= '0'; uflow <= flag10(0);
            when("10") => OUTM <= temp(2) & "111" & X"FF" & "1000" & X"000000000000"; NaN <= '1'; oflow <= '0'; uflow <= '0';
            when("11") => OUTM <= temp(2) & "111" & X"FF" & X"0000000000000"; NaN <= '0'; oflow <= flag10(1); uflow <= '0';
            when others => null; 
          end case;
          else
            OUTM <= temp(2) & fexp11 & fman11; NaN <= '0'; oflow <='0'; uflow <= '0';
          end if;
          tag_out <= tag11;
        else
          rdy12 <= '0';
        end if;
      end if;
    end if;
  end process stage_12;

  pipeline_stall <= (rdy12 and (not accept_rdy));
  muli_rdy <= not (rdy12 and (not accept_rdy));  
  mulo_rdy <= rdy12;


end rtl;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- An IEEE-754 compliant arbitrary-precision pipelined adder/subtractor
-- which is basically, a 3-stage pipelined version of the add function
-- described in the ieee_proposed VHDL library float_pkg_c.vhd
-- originally written by David Bishop (dbishop@vhdl.org)
-- modified by Madhav Desai.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir_ieee_proposed;
use ahir_ieee_proposed.float_pkg.all;
use ahir_ieee_proposed.math_utility_pkg.all;

library ahir;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;


entity GenericFloatingPointAdderSubtractor is
  generic (name: string; tag_width : integer := 8;
           exponent_width: integer := 8;
           fraction_width : integer := 23;
           round_style : round_type := float_round_style;  -- rounding option
           addguard       : NATURAL := float_guard_bits;  -- number of guard bits
           check_error : BOOLEAN    := float_check_error;  -- check for errors
           denormalize : BOOLEAN    := float_denormalize;  -- Use IEEE extended FP           
	   use_as_subtractor: BOOLEAN := false
           );
  port(
    INA, INB: in std_logic_vector((exponent_width+fraction_width) downto 0);
    OUTADD: out std_logic_vector((exponent_width+fraction_width) downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    env_rdy, accept_rdy: in std_logic;
    addi_rdy, addo_rdy: out std_logic);
end entity;


-- architecture trivial of GenericFloatingPointAdderSubtractor is
	-- 
	-- signal stage_full, stall: std_logic;
  	-- signal lp, rp   : UNRESOLVED_float(exponent_width downto -fraction_width);  -- floating point input
-- begin
  -- -- construct l,r (user registers)
  -- lp <= to_float(INA, exponent_width, fraction_width);
 -- 
  -- AsAdder: if (not use_as_subtractor) generate
  	-- rp <= to_float(INB, exponent_width, fraction_width);
  -- end generate AsAdder;
-- 
  -- AsSubtractor: if (use_as_subtractor) generate
        -- process(INB)
           -- variable btmp: UNRESOLVED_float(exponent_width downto -fraction_width);
        -- begin
	   -- btmp := to_float(INB, exponent_width, fraction_width);
  	   -- rp <= - btmp;
	-- end process;
  -- end generate AsSubtractor;
-- 
  -- stall <= stage_full and (not accept_rdy);
  -- addi_rdy <= not stall;
  -- addo_rdy <= stage_full;
-- 
  -- process(clk)
  -- begin
	-- if(clk'event and clk = '1') then
		-- if(reset = '1') then
			-- stage_full <= '0';
		-- elsif stall = '0' then
			-- stage_full <= env_rdy;
		-- end if;
-- 
		-- if(stall = '0') then
			-- OUTADD <= to_slv(lp + rp);
		-- end if;
	-- end if;
  -- end process;
-- 
-- 
-- end trivial;


-- this is the pipelined version. works, and when synthesized
-- by xst 10.1 is ok.  synthesis produces incorrect circuit with
-- xst 9.2i.
architecture rtl of GenericFloatingPointAdderSubtractor is
  signal  l, r, l_1, r_1, lp, rp   : UNRESOLVED_float(exponent_width downto -fraction_width);  -- floating point input
  
  signal pipeline_stall : std_logic;
  signal stage_full : std_logic_vector(0 to 7);
  signal tag0, tag1, tag2, tag3, tag4, tag5, tag6, tag7: std_logic_vector(tag_width-1 downto 0);

  signal fpresult_1         : UNRESOLVED_float (exponent_width downto -fraction_width);
  signal fractl_1, fractr_1   : UNSIGNED (fraction_width+1+addguard downto 0);  -- fractions
  signal exponr_1, exponl_1 : SIGNED (exponent_width-1 downto 0);  -- result exponent
  signal sign_1             : STD_ULOGIC;   -- sign of the output
  signal exceptional_result_1 : std_ulogic; 
  signal shift_too_low_1, shift_too_high_1, shift_eq_zero_1, shift_lt_zero_1, shift_gt_zero_1: boolean;
  signal shiftx_1           : SIGNED (exponent_width downto 0);  -- shift fractions

  signal use_shifter_2  : std_ulogic;
  signal shifter_in_2, shifter_out   : UNSIGNED (fraction_width+1+addguard downto 0);  -- fractions
  signal shift_amount_2 : SIGNED (exponent_width downto 0);  -- shift fractions
  
  signal fpresult_2         : UNRESOLVED_float (exponent_width downto -fraction_width);
  signal rexpon_2           : SIGNED (exponent_width downto 0);  -- result exponent
  signal fractc_2, fracts_2 : UNSIGNED (fraction_width+1+addguard downto 0);  -- constant and shifted variables
  signal leftright_2 : boolean;
  signal sticky_2_vector: std_logic_vector(0 to 4);
  signal sticky_2: std_logic;
  signal exceptional_result_2 : std_ulogic; 
  signal sign_l_2, sign_r_2: std_ulogic;




  signal shifter_tag_in, shifter_tag_out: 
		std_logic_vector(tag_width + fpresult_2'length + fractc_2'length + fracts_2'length
				+ rexpon_2'length + 7 - 1 downto 0);
  signal shifter_full: std_logic;

  signal fpresult_4         : UNRESOLVED_float (exponent_width downto -fraction_width);
  signal addL_4             : UNSIGNED (fraction_width+1+addguard downto 0);
  signal addR_4             : UNSIGNED (fraction_width+1+addguard downto 0);
  signal subtract_4         : std_logic;
  signal rexpon_4           : SIGNED (exponent_width downto 0);  -- result exponent
  signal sign_4             : STD_ULOGIC;   -- sign of the output
  signal sticky_4           : STD_ULOGIC;   -- Holds precision for rounding
  signal exceptional_result_4 : std_ulogic; 

  signal ufract_5           : UNSIGNED (fraction_width+1+addguard downto 0);
  signal fpresult_5         : UNRESOLVED_float (exponent_width downto -fraction_width);
  signal adder_tag_in, adder_tag_out :
		std_logic_vector(tag_width + fpresult_4'length + rexpon_4'length + 3 - 1 downto 0);

  signal normalizer_tag_in, normalizer_tag_out: std_logic_vector(tag_width + fpresult_4'length downto 0);

  signal fpresult_6         : UNRESOLVED_float (exponent_width downto -fraction_width);

  signal fpresult_7         : std_logic_vector((exponent_width+fraction_width) downto 0);
  
  type FracMaskArray is array (natural range <> ) of unsigned(fractl_1'length-1 downto 0);
  function BuildFracMasks(width: natural) return FracMaskArray is
	variable ret_var: FracMaskArray(width-1 downto 0);
  begin
	for I in 0 to width-1 loop
		ret_var(I) := (others => '0');
		for J in 0 to I loop
			ret_var(I)(J) := '1';
		end loop;
	end loop;
	return(ret_var);
  end function BuildFracMasks;

  constant frac_masks: FracMaskArray(fractl_1'high downto fractl_1'low) := BuildFracMasks(fractl_1'length);
  constant SH: integer := frac_masks'high;
  constant SL: integer := frac_masks'low;
  function SelectFracMask(constant masks: FracMaskArray; shiftx: integer) 
	return unsigned is
	variable ret_mask: unsigned(SH downto SL);
  begin
	ret_mask := (others => '1');
	if(shiftx <= SH) then
		ret_mask := masks(shiftx);
	elsif (shiftx < 0) then
		ret_mask := (others => '0');
	end if;
	return(ret_mask);
  end function SelectFracMask;
begin

  pipeline_stall <= stage_full(7) and (not accept_rdy);
  addi_rdy <= not pipeline_stall;
  addo_rdy <= stage_full(7);
  tag_out <= tag7;

  -- construct l,r (user registers)
  lp <= to_float(INA, exponent_width, fraction_width);
 
  AsAdder: if (not use_as_subtractor) generate
  	rp <= to_float(INB, exponent_width, fraction_width);
  end generate AsAdder;

  AsSubtractor: if (use_as_subtractor) generate
        process(INB)
           variable btmp: UNRESOLVED_float(exponent_width downto -fraction_width);
        begin
	   btmp := to_float(INB, exponent_width, fraction_width);
  	   rp <= - btmp;
	end process;
  end generate AsSubtractor;

  -- return slv.
  OUTADD <= fpresult_7;

  -----------------------------------------------------------------------------
  -- Stage 0: register inputs.
  -----------------------------------------------------------------------------
  process(clk, env_rdy, pipeline_stall, reset)
    variable active_v : std_logic;
  begin
    active_v := env_rdy and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
      	stage_full(0) <= '0';
      elsif (pipeline_stall = '0') then
        stage_full(0) <= env_rdy;
      end if;

      if(active_v = '1') then
        tag0 <= tag_in;
        l <= lp;
        r <= rp;
      end if;
    end if;
  end process;
  
  -----------------------------------------------------------------------------
  -- Stage 1: detect NaN, deNorm, align exponents.
  -----------------------------------------------------------------------------
  process(clk, l, r, reset, pipeline_stall, stage_full)
    variable active_v : std_logic;
    variable lfptype, rfptype : valid_fpstate;
    variable fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable fractl, fractr   : UNSIGNED (fraction_width+1+addguard downto 0);  -- fractions
    variable fractc, fracts   : UNSIGNED (fraction_width+1+addguard downto 0);  -- constant and shifted variables
    variable urfract, ulfract : UNSIGNED (fraction_width downto 0);
    variable ufract           : UNSIGNED (fraction_width+1+addguard downto 0);
    variable exponl, exponr   : SIGNED (exponent_width-1 downto 0);  -- exponents
    variable rexpon           : SIGNED (exponent_width downto 0);  -- result exponent
    variable shiftx           : SIGNED (exponent_width downto 0);  -- shift fractions
    variable sign             : STD_ULOGIC;   -- sign of the output
    variable leftright        : BOOLEAN;      -- left or right used
    variable lresize, rresize : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable exceptional_result: std_ulogic;

    variable shift_too_low : boolean;
    variable shift_lt_zero : boolean;
    variable shift_eq_zero : boolean;
    variable shift_too_high : boolean;
    variable shift_gt_zero : boolean;

    variable sticky           : std_logic_vector(0 to 4);   -- Holds precision for rounding
  begin

    exceptional_result := '0';
    sticky := (others => '0');
    leftright := false;
    fracts := (others => '0');
    fractc := (others => '0');
    rexpon := (others => '0');
    fpresult := (others => '0');
   
    fractr := (others => '0');
    fractl := (others => '0');

    shift_too_low := false;
    shift_lt_zero := false;
    shift_eq_zero := false;
    shift_too_high := false;
    shift_gt_zero := false;
  
    exponl := (others => '0');
    exponr := (others => '0');

    shiftx := (others => '0');

    ---------------------------------------------------------------------------
    -- will need to set appropriate flags here!
    ---------------------------------------------------------------------------
    if (fraction_width = 0 or l'length < 7 or r'length < 7) then
      lfptype := isx;
    else
      lfptype := classfp (l, check_error);
      rfptype := classfp (r, check_error);
    end if;
    if (lfptype = isx or rfptype = isx) then
      fpresult := (others => 'X');
      exceptional_result := '1';
    elsif (lfptype = nan or lfptype = quiet_nan or
           rfptype = nan or rfptype = quiet_nan)
      -- Return quiet NAN, IEEE754-1985-7.1,1
      or (lfptype = pos_inf and rfptype = neg_inf)
      or (lfptype = neg_inf and rfptype = pos_inf) then
      -- Return quiet NAN, IEEE754-1985-7.1,2
      exceptional_result := '1';
      fpresult := qnanfp (fraction_width => fraction_width,
                          exponent_width => exponent_width);
    elsif (lfptype = pos_inf or rfptype = pos_inf) then   -- x + inf = inf
      exceptional_result := '1';
      fpresult := pos_inffp (fraction_width => fraction_width,
                             exponent_width => exponent_width);
    elsif (lfptype = neg_inf or rfptype = neg_inf) then   -- x - inf = -inf
      exceptional_result := '1';
      fpresult := neg_inffp (fraction_width => fraction_width,
                             exponent_width => exponent_width);
    elsif (lfptype = neg_zero and rfptype = neg_zero) then   -- -0 + -0 = -0
      exceptional_result := '1';
      fpresult := neg_zerofp (fraction_width => fraction_width,
                             exponent_width => exponent_width);
    else 
      lresize := resize (arg            => to_x01(l),
                           exponent_width => exponent_width,
                           fraction_width => fraction_width,
                           denormalize_in => denormalize,
                           denormalize    => denormalize);
      lfptype := classfp (lresize, false);    -- errors already checked
      rresize := resize (arg            => to_x01(r),
                           exponent_width => exponent_width,
                           fraction_width => fraction_width,
                           denormalize_in => denormalize,
                           denormalize    => denormalize);
      rfptype := classfp (rresize, false);    -- errors already checked
      break_number (
          arg         => lresize,
          fptyp       => lfptype,
          denormalize => denormalize,
          fract       => ulfract,
          expon       => exponl);
      fractl := (others => '0');
      fractl (fraction_width+addguard downto addguard) := ulfract;
      break_number (
        arg         => rresize,
        fptyp       => rfptype,
        denormalize => denormalize,
        fract       => urfract,
        expon       => exponr);
      fractr := (others => '0');
      fractr (fraction_width+addguard downto addguard) := urfract;
  
      shiftx := (exponl(exponent_width-1) & exponl) - exponr;
  
      shift_too_low := (shiftx < -fractl'high);
      shift_lt_zero := (shiftx < 0);
      shift_eq_zero := (shiftx = 0);
      shift_too_high := (shiftx > fractl'high);
      shift_gt_zero := (shiftx > 0);
    end if;

    active_v := stage_full(0) and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
	stage_full(1) <= '0';
      elsif (pipeline_stall = '0') then
	stage_full(1) <= stage_full(0);
      end if;

      if(active_v = '1') then
        tag1 <= tag0;
        fpresult_1 <= fpresult;
        fractr_1 <= fractr;
        fractl_1 <= fractl;
        exponr_1 <= exponr;
 	exponl_1 <= exponl;
        exceptional_result_1 <= exceptional_result;
        l_1 <= l;
        r_1 <= r;

	shift_too_low_1 <= shift_too_low;
	shift_lt_zero_1 <= shift_lt_zero;
	shift_eq_zero_1 <= shift_eq_zero;
	shift_too_high_1 <= shift_too_high;
	shift_gt_zero_1 <= shift_gt_zero;

        shiftx_1 <= shiftx;
      end if;        
    end if;
  end process;

  -----------------------------------------------------------------------------
  -- Stage 2: detect NaN, deNorm, align exponents.
  -----------------------------------------------------------------------------
  process(clk, reset, pipeline_stall, stage_full, fpresult_1, fractr_1, exceptional_result_1, shift_too_low_1, shift_lt_zero_1, shift_eq_zero_1,
				shift_too_high_1, shift_gt_zero_1, shiftx_1, exponr_1, exponl_1)
    variable active_v : std_logic;
    variable lfptype, rfptype : valid_fpstate;
    variable fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable fractl, fractr   : UNSIGNED (fraction_width+1+addguard downto 0);  -- fractions
    variable fractc, fracts   : UNSIGNED (fraction_width+1+addguard downto 0);  -- constant and shifted variables
    variable urfract, ulfract : UNSIGNED (fraction_width downto 0);
    variable ufract           : UNSIGNED (fraction_width+1+addguard downto 0);
    variable exponl, exponr   : SIGNED (exponent_width-1 downto 0);  -- exponents
    variable rexpon           : SIGNED (exponent_width downto 0);  -- result exponent
    variable shiftx           : SIGNED (exponent_width downto 0);  -- shift fractions
    variable leftright        : BOOLEAN;      -- left or right used
    variable lresize, rresize : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable exceptional_result: std_ulogic;

    -- to get stuff to the shifter.
    variable use_shifter  : std_ulogic;
    variable shifter_in   : UNSIGNED (fraction_width+1+addguard downto 0);  -- fractions
    variable shift_amount : SIGNED (exponent_width downto 0);  -- shift fractions

    variable shift_too_low : boolean;
    variable shift_lt_zero : boolean;
    variable shift_eq_zero : boolean;
    variable shift_too_high : boolean;
    variable shift_gt_zero : boolean;

    variable sticky           : std_logic_vector(0 to 4);   -- Holds precision for rounding
  begin
    fpresult := fpresult_1;

    fractr   := fractr_1;
    fractl   := fractl_1;

    rexpon   := (others => '0');


    exceptional_result := exceptional_result_1;

    shift_too_low := shift_too_low_1;
    shift_lt_zero := shift_lt_zero_1;
    shift_eq_zero := shift_eq_zero_1;
    shift_too_high := shift_too_high_1;
    shift_gt_zero := shift_gt_zero_1;
     
    shiftx := shiftx_1;

    exponr   := exponr_1;
    exponl   := exponl_1;
    fractc := (others => '0');
    fracts := (others => '0');
    leftright := false;
    sticky := (others => '0');
    use_shifter := '0';

    shifter_in := (others  => '0');
    shift_amount :=  (others => '0');

    if shift_too_low then
        rexpon    := exponr(exponent_width-1) & exponr;
        fractc    := fractr;
        fracts    := (others => '0');   -- add zero
        leftright := false;
        sticky(0)    := or_reduce (fractl);
    elsif shift_lt_zero then
        shiftx    := - shiftx;

        shift_amount := shiftx;
        use_shifter := '1';
        shifter_in := fractl;

        -- fracts    := shift_right (fractl, to_integer(shiftx));
        fractc    := fractr;
        rexpon    := exponr(exponent_width-1) & exponr;
        leftright := false;
        --sticky(1)    := smallfract (fractl, to_integer(shiftx));
        sticky(1)    := OrReduce(fractl and SelectFracMask(frac_masks,to_integer(shiftx)));
    elsif shift_eq_zero then
        rexpon := exponl(exponent_width-1) & exponl;
        sticky(2) := '0';
        if fractr > fractl then
          fractc    := fractr;
          fracts    := fractl;
          leftright := false;
        else
          fractc    := fractl;
          fracts    := fractr;
          leftright := true;
        end if;
    elsif shift_too_high then
        rexpon    := exponl(exponent_width-1) & exponl;
        fracts    := (others => '0');   -- add zero
        fractc    := fractl;
        leftright := true;
        sticky(3)    := or_reduce (fractr);
    elsif shift_gt_zero then

        shift_amount := shiftx;
        use_shifter := '1';
        shifter_in := fractr;

        -- fracts    := shift_right (fractr, to_integer(shiftx));
        fractc    := fractl;
        rexpon    := exponl(exponent_width-1) & exponl;
        leftright := true;
        -- sticky(4) := smallfract (fractr, to_integer(shiftx));
        sticky(1)    := OrReduce(fractr and SelectFracMask(frac_masks,to_integer(shiftx)));
    end if;
    
    active_v := stage_full(1) and not (pipeline_stall or reset);

    if(clk'event and clk = '1') then

      if(reset = '1') then
	stage_full(2) <= '0';
      elsif (pipeline_stall = '0') then
	stage_full(2) <= stage_full(1);
      end if;

      if(active_v = '1') then
        tag2 <= tag1;

        fpresult_2 <= fpresult;
        fractc_2 <= fractc;
        fracts_2 <= fracts;
        rexpon_2 <= rexpon;
        leftright_2 <= leftright;
        sticky_2_vector <= sticky;
        exceptional_result_2 <= exceptional_result;
	use_shifter_2 <= use_shifter;
        sign_l_2 <= l_1(l'high);
        sign_r_2 <= r_1(r'high);


	shift_amount_2 <= shift_amount;
	shifter_in_2 <= shifter_in;

        
      end if;        
    end if;
  end process;

  sticky_2 <= OrReduce(sticky_2_vector);

  -----------------------------------------------------------------------------
  -- stage 3: shifter.
  -----------------------------------------------------------------------------
  process(tag2, fpresult_2, fractc_2, fracts_2,rexpon_2, leftright_2,
		exceptional_result_2, use_shifter_2, sign_l_2, sign_r_2, sticky_2)
  begin
        -- concatenate the tag as well!
  	shifter_tag_in(shifter_tag_in'high downto 7) <= 
		tag2 & 
		Float_To_SLV(fpresult_2) & std_logic_vector(fractc_2) &
			std_logic_vector(fracts_2) & std_logic_vector(rexpon_2);
	shifter_tag_in(6) <= '0'; -- unused.
	if(leftright_2) then
		shifter_tag_in(5) <= '1';
	else
		shifter_tag_in(5) <= '0';
	end if;
	shifter_tag_in(4) <= sticky_2;
	shifter_tag_in(3) <= exceptional_result_2;
	shifter_tag_in(2) <= sign_l_2;
	shifter_tag_in(1) <= sign_r_2;
	shifter_tag_in(0) <= use_shifter_2;
 end process;

  shifter: UnsignedShifter generic map(name => name & "-shifter", 
					shift_right_flag => true,
					tag_width => shifter_tag_in'length,
					operand_width => shifter_in_2'length,
					shift_amount_width => shift_amount_2'length)
		port map( L => shifter_in_2, R => unsigned(shift_amount_2),
				RESULT => shifter_out,
				clk => clk, reset => reset,
				in_rdy => stage_full(2),
				out_rdy => stage_full(3),
				stall => pipeline_stall,
				tag_in => shifter_tag_in,
				tag_out => shifter_tag_out);


  -----------------------------------------------------------------------------
  -- Stage 4: prepare date for mantissa adder
  -----------------------------------------------------------------------------
  process(clk, reset, pipeline_stall, stage_full, shifter_out, shifter_tag_out)
    variable active_v : std_logic;
    variable lfptype, rfptype : valid_fpstate;
    variable fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable fractl, fractr   : UNSIGNED (fraction_width+1+addguard downto 0);  -- fractions
    variable fractc, fracts   : UNSIGNED (fraction_width+1+addguard downto 0);  -- constant and shifted variables
    variable urfract, ulfract : UNSIGNED (fraction_width downto 0);
    variable rexpon           : SIGNED (exponent_width downto 0);  -- result exponent
    variable shiftx           : SIGNED (exponent_width downto 0);  -- shift fractions
    variable sign,sign_l,sign_r          : STD_ULOGIC;   -- sign of the output
    variable leftright        : BOOLEAN;      -- left or right used
    variable sticky           : STD_ULOGIC;   -- Holds precision for rounding
    variable exceptional_result           : STD_ULOGIC;   -- set if exceptional.. Nan/-Zero/Inf
    variable tagv: std_logic_vector(tag_width-1 downto 0);
    variable use_shifter: std_logic;

    variable addL, addR : UNSIGNED (fraction_width+1+addguard downto 0); 
    variable subtract_v : std_logic;
    
  begin

    subtract_v := '0';
    addL := (others => '0');
    addR := (others => '0');

    tagv := shifter_tag_out(shifter_tag_out'high downto (shifter_tag_out'high - (tag_width-1)));
    fpresult := to_float(shifter_tag_out(shifter_tag_out'high - tag_width downto 
					(shifter_tag_out'high-(tag_width + fpresult'length - 1))),
					exponent_width, fraction_width);

    fractc := unsigned(shifter_tag_out((shifter_tag_out'high- (tag_width + fpresult'length)) downto 
					(shifter_tag_out'high-
						(tag_width + fpresult'length+fractc'length - 1))));
    fracts :=  unsigned(shifter_tag_out((shifter_tag_out'high-
					(tag_width + fpresult'length+fractc'length)) downto 
					(shifter_tag_out'high-
						(tag_width + fpresult'length+(2*fractc'length) - 1))));
    rexpon :=   signed(shifter_tag_out((shifter_tag_out'high-
					(tag_width + fpresult'length+(2*fractc'length))) downto 
					(shifter_tag_out'high-
					(tag_width + fpresult'length+(2*fractc'length)+rexpon'length-1))));

    sign := '0';

    if(shifter_tag_out(5)= '1') then
	leftright := true;
    else
	leftright := false;
    end if;
    sticky := shifter_tag_out(4);
    exceptional_result := shifter_tag_out(3);
    sign_l := shifter_tag_out(2);
    sign_r := shifter_tag_out(1);
    use_shifter := shifter_tag_out(0);

    if(use_shifter = '1') then
       fracts := shifter_out;
    end if;

      -- add
    fracts (0) := fracts (0) or sticky;     -- Or the sticky bit into the LSB

    -- inputs to the adder
    addL := fractc;
    addR := fracts;
    if sign_l = sign_r then
      -- ufract := fractc + fracts;
      sign   := sign_l;
    else                              -- signs are different
      subtract_v := '1';
      -- ufract := fractc - fracts;      -- always positive result
      if leftright then               -- Figure out which sign to use
        sign := sign_l;
      else
        sign := sign_r;
      end if;
    end if;
   

    active_v := stage_full(3) and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
	stage_full(4) <= '0';
      elsif (pipeline_stall = '0') then
	stage_full(4) <= stage_full(3);
      end if;

      if(active_v = '1') then
        tag4 <= tagv;
        fpresult_4 <= fpresult;
        rexpon_4 <= rexpon;
        sign_4 <= sign;
        sticky_4 <= sticky;
        exceptional_result_4 <= exceptional_result;
        addL_4 <= addL;
	addR_4 <= addR;
	subtract_4 <= subtract_v;
      end if;      
    end if;
  end process;

  -----------------------------------------------------------------------------
  -- Stage 5: mantissa adder.
  -----------------------------------------------------------------------------
  process(tag4, fpresult_4, rexpon_4, sign_4, sticky_4, exceptional_result_4)
  begin
	adder_tag_in(adder_tag_in'high downto 3)
		<= tag4 & Float_To_SLV(fpresult_4) & std_logic_vector(rexpon_4);
	adder_tag_in(2) <= sign_4;
	adder_tag_in(1) <= sticky_4;
	adder_tag_in(0) <= exceptional_result_4;
  end process;

  adder: UnsignedAdderSubtractor
		generic map(name => name & "-adder",
				tag_width => adder_tag_in'length,
				operand_width => addL_4'length,
				chunk_width => 32)
		port map( L => addL_4, R => addR_4, RESULT => ufract_5,
				subtract_op => subtract_4,
				clk => clk, reset => reset,
				in_rdy => stage_full(4),
				out_rdy => stage_full(5),
				stall => pipeline_stall,
				tag_in => adder_tag_in,
				tag_out => adder_tag_out);
				

  -----------------------------------------------------------------------------
  -- Stage 6: normalize.
  -----------------------------------------------------------------------------
  normalizer: block
    signal tagv: std_logic_vector(tag_width-1 downto 0);
    signal fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    signal rexpon           : SIGNED (exponent_width downto 0);  -- result exponent
    signal rexpon_padded    : SIGNED (exponent_width+1 downto 0);  -- result exponent
    signal sign             : STD_ULOGIC;   -- sign of the output
    signal sticky           : STD_ULOGIC;   -- Holds precision for rounding
    signal exceptional_result           : STD_ULOGIC;   -- set if exceptional.. Nan/-Zero/Inf
    signal ufract           : UNSIGNED (fraction_width+1+addguard downto 0);
  begin
    tagv <= adder_tag_out(adder_tag_out'high downto (adder_tag_out'high - (tagv'length-1)));
    fpresult <= to_float(adder_tag_out((adder_tag_out'high - tagv'length) downto 
				(adder_tag_out'high - (tagv'length+fpresult'length-1))),
			exponent_width, fraction_width);
    rexpon <= signed(adder_tag_out((adder_tag_out'high - (tagv'length+fpresult'length)) downto 
				(adder_tag_out'high - (tagv'length+fpresult'length+rexpon'length-1))));
    rexpon_padded <= resize(rexpon,exponent_width+2);
    ufract <= ufract_5;

    -- zero fraction => sign = '0'
    sign <= '0' when or_reduce(ufract) = '0' else adder_tag_out(2);

    sticky <= adder_tag_out(1);
    exceptional_result <= adder_tag_out(0);

    
    normalizer_tag_in(normalizer_tag_in'high downto 1) <= tagv & Float_To_SLV(fpresult);
    normalizer_tag_in(0) <= exceptional_result;

    normalizer: GenericFloatingPointNormalizer
		generic map (name => name & "-normalizer",
				tag_width => normalizer_tag_in'length,
				exponent_width => exponent_width,
				fraction_width => fraction_width,
				round_style => float_round_style,
				nguard => addguard,
				denormalize => denormalize)
		port map(fract => ufract,
			 expon => rexpon_padded,
			 sign => sign,
			 sticky => sticky,
			 in_rdy  => stage_full(5),
			 out_rdy => stage_full(6),
			 stall => pipeline_stall,
			 clk => clk,
			 reset => reset,
			 tag_in => normalizer_tag_in,
			 tag_out => normalizer_tag_out,
			 normalized_result => fpresult_6);
  end block;

  -----------------------------------------------------------------------------
  -- Stage 7: multiplexor.
  -----------------------------------------------------------------------------
  process(clk, reset, pipeline_stall, stage_full, normalizer_tag_out)
    variable active_v : std_logic;
    variable fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable fpresult_normalized         : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable exceptional_result           : STD_ULOGIC;   -- set if exceptional.. Nan/-Zero/Inf
    variable tagv: std_logic_vector(tag_width-1 downto 0);
  begin

    tagv := normalizer_tag_out(normalizer_tag_out'high downto (normalizer_tag_out'high - (tagv'length-1)));
    fpresult := to_float(normalizer_tag_out((normalizer_tag_out'high - tagv'length) downto 
				(normalizer_tag_out'high - (tagv'length+fpresult'length-1))),
			exponent_width, fraction_width);
    exceptional_result := normalizer_tag_out(0);

    active_v := stage_full(6) and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
	stage_full(7) <= '0';
      elsif (pipeline_stall = '0') then
	stage_full(7) <= stage_full(6);
      end if;

      if(active_v = '1') then
        tag7 <= tagv;
    	if(exceptional_result = '1') then 
        	fpresult_7 <= to_slv(fpresult);
	else
        	fpresult_7 <= to_slv(fpresult_6);
	end if;
      end if;
    end if;
  end process;
  
end rtl;


------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- An IEEE-754 compliant arbitrary-precision pipelined multiplier
-- which is basically, a pipelined version of the multiply function
-- described in the ahir_ieee_proposed VHDL library float_pkg_c.vhd
-- originally written by David Bishop (dbishop@vhdl.org)
-- modified by Madhav Desai.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir_ieee_proposed;
use ahir_ieee_proposed.float_pkg.all;
use ahir_ieee_proposed.math_utility_pkg.all;

library ahir;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;


entity GenericFloatingPointMultiplier is
  generic (name:string;
	  tag_width : integer := 8;
           exponent_width: integer := 11;
           fraction_width : integer := 52;
           round_style : round_type := float_round_style;  -- rounding option
           addguard       : NATURAL := float_guard_bits;  -- number of guard bits
           check_error : BOOLEAN    := float_check_error;  -- check for errors
           denormalize : BOOLEAN    := float_denormalize  -- Use IEEE extended FP           
           );
  port(
    INA, INB: in std_logic_vector((exponent_width+fraction_width) downto 0);
    OUTMUL: out std_logic_vector((exponent_width+fraction_width) downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    env_rdy, accept_rdy: in std_logic;
    muli_rdy, mulo_rdy: out std_logic);
end entity;

-- works, also when synthesized by xst 10.1.  xst 9.2is seems
-- to produce incorrect circuits.
architecture rtl of GenericFloatingPointMultiplier is

  constant operand_width : integer := exponent_width+fraction_width+1;

  signal lp, rp             : UNRESOLVED_float(exponent_width downto -fraction_width);  -- floating point input  
  signal pipeline_stall : std_logic;
  signal stage_full : std_logic_vector(0 to 4);


  constant multguard        : NATURAL := addguard;           -- guard bits


  -- stage 0 outputs.
  signal tag0: std_logic_vector(tag_width-1 downto 0);
  signal  l, r             : UNRESOLVED_float(exponent_width downto -fraction_width);  -- floating point input  

  -- stage 1 outputs
  signal lfptype_1, rfptype_1 : valid_fpstate;
  signal fpresult_1         : UNRESOLVED_float (exponent_width downto -fraction_width);
  signal fractl_1, fractr_1   : UNSIGNED (fraction_width downto 0);  -- fractions
  signal rfract_1           : UNSIGNED ((2*(fraction_width))+1 downto 0);  -- result fraction
  signal sfract_1           : UNSIGNED (fraction_width+1+multguard downto 0);  -- result fraction
  signal shifty_1           : INTEGER;      -- denormal shift
  signal exponl_1, exponr_1   : SIGNED (exponent_width-1 downto 0);  -- exponents
  signal rexpon_1           : SIGNED (exponent_width+1 downto 0);  -- result exponent
  signal fp_sign_1          : STD_ULOGIC;   -- sign of result
  signal lresize_1, rresize_1 : UNRESOLVED_float (exponent_width downto -fraction_width);
  signal sticky_1           : STD_ULOGIC;   -- Holds precision for rounding
  signal exceptional_result_1  : std_logic;
  
  signal tag1: std_logic_vector(tag_width-1 downto 0);
  signal tag1_extended : std_logic_vector(tag_width+operand_width+(exponent_width+2)+1+1-1 downto 0);  

  -- stage 2 outputs (note stage 2 itelf is a pipelined array multiplier)
  signal rfract_2           : UNSIGNED ((2*(fraction_width))+1 downto 0);  -- result fraction  
  signal tag2_extended : std_logic_vector(tag_width+operand_width+(exponent_width+2)+1+1-1 downto 0);

  -- normalizer
  signal normalizer_tag_in, normalizer_tag_out: std_logic_vector(tag_width+fpresult_1'length downto 0);
  signal fpresult_3         : UNRESOLVED_float (exponent_width downto -fraction_width);

  -- stage 4 outputs.
  signal tag4: std_logic_vector(tag_width-1 downto 0);  
  signal fpresult_4         : std_logic_vector((exponent_width+fraction_width) downto 0);
  
begin

  pipeline_stall <= stage_full(4) and (not accept_rdy);
  muli_rdy <= not pipeline_stall;
  mulo_rdy <= stage_full(4);
  tag_out <= tag4;

  -- construct l,r.
  lp <= to_float(INA, exponent_width, fraction_width);
  rp <= to_float(INB, exponent_width, fraction_width);

  -- return slv.
  OUTMUL <= fpresult_4;

  -----------------------------------------------------------------------------
  -- Stage 0: register inputs.
  -----------------------------------------------------------------------------
  process(clk, reset, pipeline_stall, stage_full, env_rdy)
    variable active_v : std_logic;
  begin
    active_v := env_rdy and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
      	stage_full(0) <= '0';
      elsif (pipeline_stall = '0') then
        stage_full(0) <= env_rdy;
      end if;

      if(active_v = '1') then
        tag0 <= tag_in;
        l <= lp;
        r <= rp;
      end if;
    end if;
  end process;

  
  -----------------------------------------------------------------------------
  -- Stage 1: detect NaN, deNorm, align exponents.
  -----------------------------------------------------------------------------
  process(clk, reset, pipeline_stall, stage_full, l, r)
    variable active_v : std_logic;
    variable exceptional_result: std_ulogic;
    variable lfptype, rfptype : valid_fpstate;
    variable fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable fractl, fractr   : UNSIGNED (fraction_width downto 0);  -- fractions
    variable rfract           : UNSIGNED ((2*(fraction_width))+1 downto 0);  -- result fraction
    variable sfract           : UNSIGNED (fraction_width+1+multguard downto 0);  -- result fraction
    variable shifty           : INTEGER;      -- denormal shift
    variable exponl, exponr   : SIGNED (exponent_width-1 downto 0);  -- exponents
    variable rexpon           : SIGNED (exponent_width+1 downto 0);  -- result exponent
    variable fp_sign          : STD_ULOGIC;   -- sign of result
    variable lresize, rresize : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable sticky           : STD_ULOGIC;   -- Holds precision for rounding
  begin
    exceptional_result := '0';    
    fp_sign := '0';
    rexpon := (others => '0');
    exponl := (others => '0');
    exponr := (others => '0');
    shifty := 0;
    fractl := (others => '0');
    fractr := (others => '0');
    lfptype := isx;
    rfptype := isx;
    fpresult := (others => '0');
     
    if (fraction_width = 0 or l'length < 7 or r'length < 7) then
      lfptype := isx;
      exceptional_result := '1';
    else
      lfptype := classfp (l, check_error);
      rfptype := classfp (r, check_error);
    end if;
    if (lfptype = isx or rfptype = isx) then
      fpresult := (others => 'X');
      exceptional_result := '1';      
    elsif ((lfptype = nan or lfptype = quiet_nan or
            rfptype = nan or rfptype = quiet_nan)) then
      -- Return quiet NAN, IEEE754-1985-7.1,1
      exceptional_result := '1';      
      fpresult := qnanfp (fraction_width => fraction_width,
                          exponent_width => exponent_width);
    elsif (((lfptype = pos_inf or lfptype = neg_inf) and
            (rfptype = pos_zero or rfptype = neg_zero)) or
           ((rfptype = pos_inf or rfptype = neg_inf) and
            (lfptype = pos_zero or lfptype = neg_zero))) then    -- 0 * inf
      -- Return quiet NAN, IEEE754-1985-7.1,3
      exceptional_result := '1';      
      fpresult := qnanfp (fraction_width => fraction_width,
                          exponent_width => exponent_width);
    elsif (lfptype = pos_inf or rfptype = pos_inf
           or lfptype = neg_inf or rfptype = neg_inf) then  -- x * inf = inf
      exceptional_result := '1';      
      fpresult := pos_inffp (fraction_width => fraction_width,
                             exponent_width => exponent_width);
      -- figure out the sign
      fp_sign := l(l'high) xor r(r'high);     -- figure out the sign
      fpresult (exponent_width) := fp_sign;
    else
      fp_sign := l(l'high) xor r(r'high);     -- figure out the sign
     
      -- mpd: this resize seems unnecessary..
      --lresize := resize (arg            => to_x01(l),
                         --exponent_width => exponent_width,
                         --fraction_width => fraction_width,
                         --denormalize_in => denormalize,
                         --denormalize    => denormalize);
      lresize := to_X01(l);

      lfptype := classfp (lresize, false);    -- errors already checked
      
      -- mpd: this resize is not necessary?
      -- rresize := resize (arg            => to_x01(r),
                         -- exponent_width => exponent_width,
                         -- fraction_width => fraction_width,
                         -- denormalize_in => denormalize,
                         -- denormalize    => denormalize);
      rresize := to_X01(r);
      rfptype := classfp (rresize, false);    -- errors already checked

      break_number (
        arg         => lresize,
        fptyp       => lfptype,
        denormalize => denormalize,
        fract       => fractl,
        expon       => exponl);
      break_number (
        arg         => rresize,
        fptyp       => rfptype,
        denormalize => denormalize,
        fract       => fractr,
        expon       => exponr);

      -- TODO: this shifter slows things down. perhaps its better to break
      --       and add a new stage at this point.
      if (rfptype = pos_denormal or rfptype = neg_denormal) then
        shifty := fraction_width - find_leftmost(fractr, '1');
        fractr := shift_left (fractr, shifty);
      elsif (lfptype = pos_denormal or lfptype = neg_denormal) then
        shifty := fraction_width - find_leftmost(fractl, '1');
        fractl := shift_left (fractl, shifty);
      else
        shifty := 0;
        -- Note that a denormal number * a denormal number is always zero.
      end if;
      -- multiply
      -- add the exponents
      rexpon := resize (exponl, rexpon'length) + exponr - shifty + 1;
    end if;

    active_v := stage_full(0) and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
	stage_full(1) <= '0';
      elsif (pipeline_stall = '0') then
	stage_full(1) <= stage_full(0);
      end if;

      if(active_v = '1') then
        tag1 <= tag0;
        
        fpresult_1 <= fpresult;
        fractl_1 <= fractl;
        fractr_1 <= fractr;
        rexpon_1 <= rexpon;
        fp_sign_1 <= fp_sign;
        exceptional_result_1 <= exceptional_result;
      end if;      
    end if;
  end process;

  -----------------------------------------------------------------------------
  -- Stage 2: instantiate array multiplier
  -----------------------------------------------------------------------------
  process(tag1, fpresult_1, rexpon_1, fp_sign_1, exceptional_result_1, fp_sign_1, exceptional_result_1)
    variable tex : std_logic_vector(tag_width+operand_width+(exponent_width+2)+1 downto 0);
    variable fp_slv : std_logic_vector(operand_width-1 downto 0);
    variable pad_bits : std_logic_vector(1 downto 0);
  begin

    fp_slv(operand_width-1) := fpresult_1(exponent_width);
    fp_slv(operand_width-2 downto fraction_width) := to_slv(fpresult_1(exponent_width-1 downto 0));
    fp_slv(fraction_width-1 downto 0) := to_slv(fpresult_1(-1 downto -fraction_width));

    pad_bits(1) := fp_sign_1;
    pad_bits(0) := exceptional_result_1;
    
    tex := tag1 & fp_slv & to_slv(rexpon_1) & pad_bits;
    
    tag1_extended <= tex;
  end process;
  
  amul : UnsignedMultiplier
    generic map (name => name & "-amul", tag_width => tag_width+operand_width+(exponent_width+2)+2,
                 operand_width => fraction_width+1,
		 chunk_width => 32)
    port map (
      L       => fractl_1,
      R       => fractR_1,
      RESULT  => rfract_2,
      clk     => clk,
      reset   => reset,
      in_rdy  => stage_full(1),
      out_rdy => stage_full(2),
      stall   => pipeline_stall,
      tag_in  => tag1_extended,
      tag_out => tag2_extended);
    


  -----------------------------------------------------------------------------
  -- Stage 3: normalize... 
  -----------------------------------------------------------------------------
  Normalizer: block
    signal rfract           : UNSIGNED ((2*(fraction_width))+1 downto 0);  -- result fraction
    signal sfract           : UNSIGNED (fraction_width+1+multguard downto 0);  -- result fraction
    signal rexpon           : SIGNED (exponent_width+1 downto 0);  -- result exponent
    signal fp_sign          : STD_ULOGIC;   -- sign of result
    signal sticky           : STD_ULOGIC;   -- Holds precision for rounding
    signal raw_tag          : std_logic_vector(tag_width-1 downto 0);
    signal fpresult         : UNRESOLVED_float (exponent_width downto -fraction_width);
    signal exceptional_result: std_logic;
  begin
    raw_tag <= tag2_extended((tag_width+operand_width+exponent_width+3) downto (operand_width+exponent_width+4));
    fpresult <= to_float(tag2_extended(operand_width+exponent_width+3 downto exponent_width+4), exponent_width, fraction_width);
    rexpon <= to_signed(tag2_extended(exponent_width+3 downto 2));
    fp_sign <= tag2_extended(1);
    exceptional_result <= tag2_extended(0);
    
    rfract <= rfract_2;
    sfract <= rfract (rfract'high downto
                      rfract'high - (fraction_width+1+multguard));
    sticky <= or_reduce (rfract (rfract'high-(fraction_width+1+multguard)
                                 downto 0));

    normalizer_tag_in(normalizer_tag_in'high downto 1) <= 
		raw_tag & Float_To_SLV(fpresult);
    normalizer_tag_in(0) <= exceptional_result;
   	
    normalizer: GenericFloatingPointNormalizer
		generic map (name => name & "-normalizer", tag_width => normalizer_tag_in'length,
				exponent_width => exponent_width,
				fraction_width => fraction_width,
				round_style => float_round_style,
				nguard => multguard,
				denormalize => denormalize)
		port map(fract => sfract,
			 expon => rexpon,
			 sign => fp_sign,
			 sticky => sticky,
			 in_rdy  => stage_full(2),
			 out_rdy => stage_full(3),
			 stall => pipeline_stall,
			 clk => clk,
			 reset => reset,
			 tag_in => normalizer_tag_in,
			 tag_out => normalizer_tag_out,
			 normalized_result => fpresult_3);
  end block;

  -----------------------------------------------------------------------------
  -- Stage 4: final multiplexor... 
  -----------------------------------------------------------------------------
  process(clk, reset, pipeline_stall, stage_full, normalizer_tag_out, fpresult_3)
    variable active_v : std_logic;
    variable exceptional_result: std_ulogic;
    variable fpresult, fpresult_normalized   : UNRESOLVED_float (exponent_width downto -fraction_width);
    variable raw_tag          : std_logic_vector(tag_width-1 downto 0);
    
  begin

    raw_tag := normalizer_tag_out(tag_width+operand_width downto operand_width+1);
    fpresult := to_float(normalizer_tag_out(operand_width downto 1), exponent_width, fraction_width);
    exceptional_result := normalizer_tag_out(0);
    
   fpresult_normalized := fpresult_3;

    active_v := stage_full(3) and not (pipeline_stall or reset);
    if(clk'event and clk = '1') then

      if(reset = '1') then
	stage_full(4) <= '0';
      elsif (pipeline_stall = '0') then
	stage_full(4) <= stage_full(3);
      end if;

      if(active_v = '1') then
        tag4 <= raw_tag;

        if(exceptional_result = '1') then
          fpresult_4 <= to_slv(fpresult);
	else
          fpresult_4 <= to_slv(fpresult_normalized);
        end if;
        
      end if;      
    end if;
  end process;
  
end rtl;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- An IEEE-754 compliant arbitrary-precision normalizer
-- originally written by David Bishop (dbishop@vhdl.org)
-- modified by Madhav Desai.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;

library ahir;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;


entity GenericFloatingPointNormalizer is
  generic (name:string; 
	   tag_width : integer := 8;
           exponent_width: integer := 11;
           fraction_width : integer := 52;
           round_style : round_type := float_round_style;  -- rounding option
           nguard       : NATURAL := float_guard_bits;  -- number of guard bits
           denormalize : BOOLEAN    := float_denormalize  -- Use IEEE extended FP           
           );
  port(
    fract  :in  unsigned(fraction_width+nguard+1 downto 0);
    expon  :in  signed(exponent_width+1 downto 0);
    sign   :in  std_ulogic;
    sticky :in  std_ulogic;
    tag_in :in  std_logic_vector(tag_width-1 downto 0);
    tag_out:out std_logic_vector(tag_width-1 downto 0);
    in_rdy :in  std_ulogic;
    out_rdy:out std_ulogic;
    stall  :in  std_ulogic;
    clk    :in  std_ulogic;
    reset  :in  std_ulogic;
    normalized_result :out UNRESOLVED_float (exponent_width downto -fraction_width)  -- result
   );
end entity;


architecture Simple of GenericFloatingPointNormalizer is

begin

	process(clk)
    	   variable result : UNRESOLVED_float (exponent_width downto -fraction_width);
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				out_rdy <= '0';
			elsif(stall = '0') then

				result := 
					normalize(fract,expon,sign,sticky,
					   	exponent_width, fraction_width,
						round_style, denormalize, 
						nguard);
				normalized_result <= result;

				tag_out <= tag_in;
				out_rdy <= in_rdy;
			end if;

			
		end if;
	end process;
end Simple;


-- this is the real stuff.
architecture rtl of GenericFloatingPointNormalizer is
    constant num_stages: integer := 6;
    constant operand_width: integer := fract'length;

    signal stage_full: std_logic_vector(0 to num_stages);

    type TagArray is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);
    signal stage_tags: TagArray(0 to num_stages);

    signal expon_1  : signed(exponent_width+1 downto 0);
    signal fract_1,fract_2,fract_3  :  unsigned(fraction_width+nguard+1 downto 0);
    signal round_1, zerores_1, infres_1 : BOOLEAN;
    signal round_2, zerores_2, infres_2 : BOOLEAN;

    signal shiftr_1,shiftr_2,shiftr_3     : INTEGER range -(2**(expon'length+1)) to (2**(expon'length+1));      -- shift amount

    signal exp_1,exp_2,exp_3        : SIGNED (exponent_width+1 downto 0);  -- exponent

    signal sticky_1,sticky_2, sticky_3    : STD_ULOGIC;   -- versions of sticky
    signal sign_1,sign_2, sign_3    : STD_ULOGIC;   -- versions of sign

    signal result_1,result_2,result_3, result_6: 
		UNRESOLVED_float (exponent_width downto -fraction_width);  -- result
    signal exceptional_result_flag_3: std_ulogic;

    signal shift_in, shift_out : unsigned(fraction_width+nguard+1 downto 0);
    signal shift_tag_in, shift_tag_out : 
		std_logic_vector(tag_width+expon'length+normalized_result'length+4-1 downto 0);
    signal shift_amount: unsigned(Ceil_Log2(fract'length)-1 downto 0);

begin

  stage_full(0) <= in_rdy;
  out_rdy <= stage_full(num_stages);

  stage_tags(0) <= tag_in;
  tag_out <= stage_tags(num_stages);

  normalized_result <= result_6;

  -------------------------------------------------------------------------------------------------------------
  -- stage 1: left-most 1
  -------------------------------------------------------------------------------------------------------------
  -- stage 1: find leftmost 1.
  process(clk)
    variable sfract     : UNSIGNED (fract'high downto 0);  -- shifted fraction
    variable rfract     : UNSIGNED (fraction_width-1 downto 0);   -- fraction
    variable exp        : SIGNED (exponent_width+1 downto 0);  -- exponent
    variable rexp       : SIGNED (exponent_width+1 downto 0);  -- result exponent
    variable rexpon     : UNSIGNED (exponent_width-1 downto 0);   -- exponent
    variable result     : UNRESOLVED_float (exponent_width downto -fraction_width);  -- result
    variable shiftr     : INTEGER range -(2**(expon'length+1)) to (2**(expon'length+1));      -- shift amount
    variable stickyx    : STD_ULOGIC;   -- version of sticky
    constant expon_base : SIGNED (exponent_width-1 downto 0) :=
      gen_expon_base(exponent_width);   -- exponent offset
    variable round, zerores, infres : BOOLEAN;
  begin  -- function normalize
    zerores := false;
    infres  := false;
    round   := false;
    shiftr  := find_leftmost (to_01(fract), '1')     -- Find the first "1"
               - fraction_width - nguard;  -- subtract the length we want
    exp := resize (expon, exp'length) + shiftr;
    if(clk'event and clk = '1') then
	if(reset = '1') then
		stage_full(1) <= '0';
	elsif(stall = '0') then
		zerores_1 <= zerores;
		infres_1  <= infres;
		round_1   <= round;
		shiftr_1  <= shiftr;
		exp_1 <= exp;
		fract_1 <= fract;
		sticky_1 <= sticky;
		sign_1 <= sign;
		expon_1 <= expon;
		stage_full(1) <= stage_full(0);
		stage_tags(1) <= stage_tags(0);
	end if;
    end if;
  end process;

  
  -------------------------------------------------------------------------------------------------------------
  -- stage 2,3,4: merged
  -------------------------------------------------------------------------------------------------------------
  process(fract_1, zerores_1, infres_1, round_1, shiftr_1, exp_1, expon_1, stage_full(1), stage_tags(1))
    variable sfract     : UNSIGNED (fract'high downto 0);  -- shifted fraction
    variable rfract     : UNSIGNED (fraction_width-1 downto 0);   -- fraction
    variable exp        : SIGNED (exponent_width+1 downto 0);  -- exponent
    variable rexp       : SIGNED (exponent_width+1 downto 0);  -- result exponent
    variable rexpon     : UNSIGNED (exponent_width-1 downto 0);   -- exponent
    variable result     : UNRESOLVED_float (exponent_width downto -fraction_width);  -- result
    variable shiftr     : INTEGER range -(2**(expon'length+1)) to (2**(expon'length+1));      -- shift amount
    variable stickyx    : STD_ULOGIC;   -- version of sticky
    constant expon_base : SIGNED (exponent_width-1 downto 0) :=
      gen_expon_base(exponent_width);   -- exponent offset
    variable round, zerores, infres : BOOLEAN;
  begin  -- function normalize
    zerores := zerores_1;
    infres  := infres_1;
    round   := round_1;
    shiftr  := shiftr_1;
    exp     := exp_1;

    if (or_reduce (fract_1) = '0') then   -- Zero
      zerores := true;
    elsif ((exp <= -resize(expon_base, exp'length)-1) and denormalize)
      or ((exp < -resize(expon_base, exp'length)-1) and not denormalize) then
      if (exp >= -resize(expon_base, exp'length)-fraction_width-1)
        and denormalize then
        exp    := -resize(expon_base, exp'length)-1;
        shiftr := -to_integer (expon_1 + expon_base);  -- new shift
      else                              -- return zero
        zerores := true;
      end if;
    elsif (exp > expon_base-1) then     -- infinity
      infres := true;
    end if;

    -- pass it to the next stage, combinationally..
    zerores_2 <= zerores;
    infres_2 <= infres;
    round_2 <= round;
    shiftr_2 <= shiftr;
    exp_2 <= exp;
    fract_2 <= fract_1;
    sticky_2 <= sticky_1;
    sign_2 <= sign_1;
    stage_full(2) <= stage_full(1);
    stage_tags(2) <= stage_tags(1);
  end process;

  -- stage 3: exceptional cases
  process(zerores_2, infres_2, round_2, shiftr_2, exp_2, fract_2, sticky_2, stage_full(2), stage_tags(2))
    variable sfract     : UNSIGNED (fract'high downto 0);  -- shifted fraction
    variable rfract     : UNSIGNED (fraction_width-1 downto 0);   -- fraction
    variable exp        : SIGNED (exponent_width+1 downto 0);  -- exponent
    variable rexp       : SIGNED (exponent_width+1 downto 0);  -- result exponent
    variable rexpon     : UNSIGNED (exponent_width-1 downto 0);   -- exponent
    variable result     : UNRESOLVED_float (exponent_width downto -fraction_width);  -- result
    variable shiftr     : INTEGER range -(2**(expon'length+1)) to (2**(expon'length+1));      -- shift amount
    variable stickyx    : STD_ULOGIC;   -- version of sticky
    constant expon_base : SIGNED (exponent_width-1 downto 0) :=
      gen_expon_base(exponent_width);   -- exponent offset
    variable round, zerores, infres : BOOLEAN;
    variable exceptional_result_flag: std_ulogic;
  begin  -- function normalize
    zerores := zerores_2;
    infres  := infres_2;
    round   := round_2;
    shiftr  := shiftr_2;
    exp     := exp_2;
    exceptional_result_flag := '0';
    result := (others => '0');

    if zerores then
      exceptional_result_flag := '1';
      result := zerofp (fraction_width => fraction_width,
                        exponent_width => exponent_width);
    elsif infres then
      exceptional_result_flag := '1';
      result := pos_inffp (fraction_width => fraction_width,
                           exponent_width => exponent_width);
    end if;
  
    fract_3 <= fract_2;	
    sticky_3 <= sticky_2;
    shiftr_3 <= shiftr;
    exp_3 <= exp;
    exceptional_result_flag_3 <= exceptional_result_flag;
    result_3 <= result;
    sign_3 <= sign_2;
    stage_full(3) <= stage_full(2);
    stage_tags(3) <= stage_tags(2);
  end process;

  
  -- stage 4:  prepare data for shifter.
  process(fract_3, sticky_3, shiftr_3, exp_3, exceptional_result_flag_3, result_3, sign_3, stage_full(3), stage_tags(3))
        variable reverse_flag, stickyx: std_ulogic;
        variable shiftu: unsigned(Ceil_Log2(fract'length)-1 downto 0);
        variable tmp: natural;
  begin 
   -- some variables depend on shift_3.
   if(shiftr_3 <= 0) then
	reverse_flag := '1';
        tmp := - shiftr_3;
	shiftu := to_unsigned(tmp,shiftu'length);
	stickyx := sticky_3;
   else 
        reverse_flag := '0';
	tmp := shiftr_3;
	shiftu := to_unsigned(tmp, shiftu'length);
	stickyx := sticky_3 or smallfract(fract_3, shiftr_3-1);
   end if;
    
    --- break 3 -----
   if(shiftr_3 <= 0) then
	shift_in <= reverse(fract_3);
   else
	shift_in <= fract_3;
   end if;
  
   shift_amount <= shiftu;

   shift_tag_in(shift_tag_in'high downto 4) <= std_logic_vector(stage_tags(3)) & 
			std_logic_vector(exp_3) & Float_To_SLV(result_3);
   shift_tag_in(3) <=  sign_3;
   shift_tag_in(2) <=  exceptional_result_flag_3;
   shift_tag_in(1) <=  reverse_flag;
   shift_tag_in(0) <=  stickyx;
   stage_full(4) <= stage_full(3);
   stage_tags(4) <= stage_tags(3);
  end process;
  
  ----------------------------------------------------------------------------------------------------------------
  -- stage 5: shifter:  sfract := fract srl shiftr;   
  ----------------------------------------------------------------------------------------------------------------
  us: UnsignedShifter generic map(name=> name & "-us", shift_right_flag => true,
					tag_width => shift_tag_in'length,
					operand_width => shift_in'length,
					shift_amount_width => shift_amount'length)
		port map(L => shift_in, R => shift_amount, RESULT => shift_out,
				clk => clk, reset => reset,
				in_rdy => stage_full(4),
				out_rdy => stage_full(5),
				stall => stall,
				tag_in => shift_tag_in,
				tag_out => shift_tag_out);


  ----------------------------------------------------------------------------------------------------------------
  -- stage 6: round.
  ----------------------------------------------------------------------------------------------------------------
  process(clk)
    variable sfract     : UNSIGNED (fract'high downto 0);  -- shifted fraction
    variable rfract     : UNSIGNED (fraction_width-1 downto 0);   -- fraction
    variable exp        : SIGNED (exponent_width+1 downto 0);  -- exponent
    variable rexp       : SIGNED (exponent_width+1 downto 0);  -- result exponent
    variable rexpon     : UNSIGNED (exponent_width-1 downto 0);   -- exponent
    variable result_exceptional   : UNRESOLVED_float (exponent_width downto -fraction_width);  -- result
    variable result     : UNRESOLVED_float (exponent_width downto -fraction_width);  -- result
    variable shiftr     : INTEGER range -(2**(expon'length+1)) to (2**(expon'length+1));      -- shift amount
    variable stickyx    : STD_ULOGIC;   -- version of sticky
    constant expon_base : SIGNED (exponent_width-1 downto 0) :=
      gen_expon_base(exponent_width);   -- exponent offset
    variable round, zerores, infres : BOOLEAN;
    variable exceptional_result_flag, reverse_flag: std_ulogic;
    variable shiftu : unsigned(Ceil_Log2(fract'length)-1 downto 0);
    variable signx: std_ulogic;
  begin  -- function normalize
    exp   := signed(shift_tag_out((shift_tag_out'high - tag_width) downto 
		(shift_tag_out'high - (tag_width+exp'length-1))));	
    result_exceptional := to_float(shift_tag_out((shift_tag_out'high - 
					(tag_width + exp'length)) downto 
				(shift_tag_out'high - (tag_width+exp'length+result'length-1))),
				exponent_width, fraction_width);	
    signx := shift_tag_out(3);
    exceptional_result_flag := shift_tag_out(2);
    reverse_flag := shift_tag_out(1);
    stickyx := shift_tag_out(0);
    result := (others => '0');
    rfract := (others => '0');

    if reverse_flag = '0' then
        sfract := shift_out;
    else
    	sfract := reverse(shift_out);
    end if;

    if nguard > 0 then
      round := check_round (
        fract_in    => sfract (nguard),
        sign        => signx,
        remainder   => sfract(nguard-1 downto 0),
        sticky      => stickyx,
        round_style => round_style);
    end if;
    if round then
      fp_round(fract_in  => sfract (fraction_width-1+nguard downto nguard),
               expon_in  => exp(rexp'range),
               fract_out => rfract,
               expon_out => rexp);
    else
      rfract := sfract (fraction_width-1+nguard downto nguard);
      rexp   := exp(rexp'range);
    end if;
      --- break 5 ----
      -- result
    rexpon := UNSIGNED (rexp(exponent_width-1 downto 0));
    rexpon (exponent_width-1)          := not rexpon(exponent_width-1);
    result (rexpon'range)              := UNRESOLVED_float(rexpon);
    result (-1 downto -fraction_width) := UNRESOLVED_float(rfract);

    result (exponent_width) := signx;    -- sign BIT

    if(clk'event and clk = '1') then
	if(reset = '1') then
		stage_full(6) <= '0';
	elsif (stall = '0') then
		if(exceptional_result_flag = '0') then
			result_6 <= result;
		else
			result_6 <= result_exceptional;
		end if;
		stage_full(6) <= stage_full(5);
		stage_tags(6) <= shift_tag_out(shift_tag_out'high downto 
					(shift_tag_out'high - (tag_width-1)));
	end if;
    end if;
  end process;

end rtl;


------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- An IEEE-754 compliant arbitrary-precision pipelined float-to-float
-- converter which is basically, a pipelined version of the resize function
-- described in the ahir_ieee_proposed VHDL library float_pkg_c.vhd
-- originally written by David Bishop (dbishop@vhdl.org)
-- modified by Madhav Desai.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir_ieee_proposed;
use ahir_ieee_proposed.float_pkg.all;
use ahir_ieee_proposed.math_utility_pkg.all;

library ahir;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;

entity GenericFloatToFloat is
  generic (name: string; 
	   tag_width : integer := 8;
           in_exponent_width: integer := 11;
           in_fraction_width : integer := 52;
           out_exponent_width: integer := 8;
           out_fraction_width : integer := 23;
           round_style : round_type := float_round_style;  -- rounding option
           addguard       : NATURAL := float_guard_bits;  -- number of guard bits
           check_error : BOOLEAN    := float_check_error;  -- check for errors
           denormalize_in : BOOLEAN := float_denormalize;  -- Use IEEE extended FP           
           denormalize : BOOLEAN    := float_denormalize  -- Use IEEE extended FP           
           );
  port(
    INF: in std_logic_vector((in_exponent_width+in_fraction_width) downto 0);
    OUTF: out std_logic_vector((out_exponent_width+out_fraction_width) downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    env_rdy, accept_rdy: in std_logic;
    f2fi_rdy, f2fo_rdy: out std_logic);
end entity;

-- works, also when synthesized by xst 10.1.  xst 9.2is seems
-- to produce incorrect circuits.
architecture rtl of GenericFloatToFloat is
        signal stage_full: std_logic_vector(1 to 2);
	signal pipeline_stall: std_logic;
	signal in_arg  : UNRESOLVED_float (in_exponent_width downto -in_fraction_width);

	signal sign_sig: std_logic;
    	signal expon_in_sig          : SIGNED (in_exponent_width-1 downto 0);
    	signal fract_in_sig          : UNSIGNED (in_fraction_width downto 0);
    	signal expon_out_sig         : SIGNED (out_exponent_width-1 downto 0);  -- output fract
    	signal fract_out_sig         : UNSIGNED (out_fraction_width downto 0);  -- output fract

	signal normalizer_result_out : std_logic_vector(OUTF'length-1 downto 0);
	signal normalizer_tag_in, normalizer_tag_out: std_logic_vector((tag_width + OUTF'length) downto 0);
begin

	in_arg <= to_float (INF, in_exponent_width, in_fraction_width);

	pipeline_stall <= stage_full(2) and (not accept_rdy);
	f2fo_rdy <= stage_full(2);
	f2fi_rdy <=  not pipeline_stall;

	-- stage 1 upto normalizer..
	process(clk, reset, pipeline_stall, stage_full, fract_in_sig)
    		variable result            : UNRESOLVED_float (out_exponent_width downto -out_fraction_width);
                                        -- result value
    		variable fptype            : valid_fpstate;
    		variable expon_in          : SIGNED (in_exponent_width-1 downto 0);
    		variable fract_in          : UNSIGNED (in_fraction_width downto 0);
    		variable round             : BOOLEAN;
    		variable expon_out         : SIGNED (out_exponent_width-1 downto 0);  -- output fract
    		variable fract_out         : UNSIGNED (out_fraction_width downto 0);  -- output fract
    		variable nguard            : NATURAL;
		variable use_normalizer : std_logic;
		variable fract_in_sign: std_logic;
    		constant check_error    : BOOLEAN    := float_check_error;
	begin
		result := (others => '0');
		expon_in := (others => '0');
		expon_out := (others => '0');
		fract_in := (others => '0');
		fract_out := (others => '0');
		nguard := 0;
		use_normalizer := '0';
		fract_in_sign := INF(in_exponent_width + in_fraction_width);

    		fptype := classfp(in_arg, check_error);
    		if ((fptype = pos_denormal or fptype = neg_denormal) and denormalize_in
        		and (in_exponent_width < out_exponent_width
             			or in_fraction_width < out_fraction_width))
      				or in_exponent_width > out_exponent_width
      				or in_fraction_width > out_fraction_width then
      			-- size reduction
      			classcase : case fptype is
        			when isx =>
          			  result := (others => 'X');
        			when nan | quiet_nan =>
          			  result := qnanfp (fraction_width => out_fraction_width,
                            				exponent_width => out_exponent_width);
        			when pos_inf =>
          			  result := pos_inffp (fraction_width => out_fraction_width,
                               				exponent_width => out_exponent_width);
        			when neg_inf =>
          			  result := neg_inffp (fraction_width => out_fraction_width,
                               				exponent_width => out_exponent_width);
        			when pos_zero | neg_zero =>
          			   result := zerofp (fraction_width => out_fraction_width,   -- hate -0
                            					exponent_width => out_exponent_width);
        			when others =>
          				break_number (
            					arg         => in_arg,
            					fptyp       => fptype,
            					denormalize => denormalize_in,
            					fract       => fract_in,
            					expon       => expon_in);
       					if out_fraction_width > in_fraction_width and denormalize_in then
						use_normalizer := '1';
           					-- You only get here if you have a denormal input
       						fract_out := (others => '0');              -- pad with zeros
       						fract_out (out_fraction_width downto
                       							out_fraction_width - in_fraction_width) := fract_in;
       						nguard := 0;
       					else
						use_normalizer := '1';
              					nguard := in_fraction_width - out_fraction_width;
          				end if;
      			end case classcase;
    		else                                -- size increase or the same size
      			if out_exponent_width > in_exponent_width then
        			expon_in := SIGNED(in_arg (in_exponent_width-1 downto 0));
        			if fptype = pos_zero or fptype = neg_zero then
          				result (out_exponent_width-1 downto 0) := (others => '0');
        			elsif expon_in = -1 then        -- inf or nan (shorts out check_error)
          				result (out_exponent_width-1 downto 0) := (others => '1');
        			else
          			-- invert top BIT
          				expon_in(expon_in'high)            := not expon_in(expon_in'high);
          				expon_out := resize (expon_in, expon_out'length);  -- signed expand
          			-- Flip it back.
          				expon_out(expon_out'high)          := not expon_out(expon_out'high);
          				result (out_exponent_width-1 downto 0) := UNRESOLVED_float(expon_out);
        			end if;
        			result (out_exponent_width) := in_arg (in_exponent_width);     -- sign
      			else                              -- exponent_width = in_exponent_width
        			result (out_exponent_width downto 0) := in_arg (in_exponent_width downto 0);
      			end if;
      			if out_fraction_width > in_fraction_width then
        			result (-1 downto -out_fraction_width) := (others => '0');  -- zeros
        			result (-1 downto -in_fraction_width) :=
          						in_arg (-1 downto -in_fraction_width);
      			else                              -- fraction_width = in_fraciton_width
        			result (-1 downto -out_fraction_width) :=
          						in_arg (-1 downto -in_fraction_width);
      			end if;
    		end if;
	
		if(clk'event and clk = '1') then
			if(reset = '1') then
				stage_full(1) <= '0';
				fract_in_sig <= (others => '0');
				fract_out_sig <= (others => '0');
				expon_in_sig <= (others => '0');
				expon_out_sig <= (others => '0');
				sign_sig <= '0';
				normalizer_tag_in <= (others =>  '0');
			elsif (pipeline_stall = '0') then
				fract_in_sig <= fract_in;
				fract_out_sig <= fract_out;
				expon_in_sig <= expon_in;
				expon_out_sig <= expon_out;
				normalizer_tag_in(0) <= use_normalizer;
				normalizer_tag_in((tag_width + result'length) downto 1) <= (tag_in & to_slv(result));
				sign_sig <= fract_in_sign;
				stage_full(1) <= env_rdy;
			end if;
		end if;
	end process;


	f2D: if (out_fraction_width >= in_fraction_width) generate
	    blk: block
			signal normalizer_fract: unsigned(out_fraction_width downto 0);
	    begin
		
		process(fract_in_sig)
		begin
			normalizer_fract  <=   (others => '0');
			normalizer_fract(in_fraction_width downto 0) <= fract_in_sig;
		end process;

		process(clk,reset,  pipeline_stall,  stage_full,  normalizer_fract)
    			variable result    : UNRESOLVED_float (out_exponent_width downto -out_fraction_width);
		begin
			result :=
				normalize (fract => normalizer_fract, 
						expon => expon_in_sig,
						sign => sign_sig,
						fraction_width => out_fraction_width,
						exponent_width => out_exponent_width,
						round_style => round_style,
						denormalize => denormalize,
						nguard => 0);

			if(clk'event and clk = '1') then
				if(reset = '1') then
					stage_full(2) <= '0';
					normalizer_tag_out <= (others => '0');
				elsif (pipeline_stall = '0') then
					stage_full(2) <= stage_full(1);
					normalizer_result_out <= to_slv(result);
					normalizer_tag_out <= normalizer_tag_in;	
				end if;
			end if;
		end process;
	    end block;
        end generate f2D;

	D2f: if (out_fraction_width < in_fraction_width) generate
		process(clk, reset, pipeline_stall, fract_in_sig, expon_in_sig, sign_sig)
    			variable result    : UNRESOLVED_float (out_exponent_width downto -out_fraction_width);
		begin
			result :=
				normalize (fract => fract_in_sig, 
						expon => expon_in_sig,
						sign => sign_sig,
						fraction_width => out_fraction_width,
						exponent_width => out_exponent_width,
						round_style => round_style,
						denormalize => denormalize,
						nguard => (in_fraction_width - out_fraction_width));

			if(clk'event and clk = '1') then
				if(reset = '1') then
					stage_full(2) <= '0';
					normalizer_tag_out <= (others => '0');
				elsif (pipeline_stall = '0') then
					stage_full(2) <= stage_full(1);
					normalizer_result_out <= to_slv(result);
					normalizer_tag_out <= normalizer_tag_in;	
				end if;
			end if;
		end process;
	end generate D2f;

	-- output multiplexor.
	OUTF <= normalizer_tag_out(OUTF'length downto 1) when
			(normalizer_tag_out(0) = '0')  else  normalizer_result_out;
	tag_out <= normalizer_tag_out((tag_width + OUTF'length) downto (OUTF'length + 1));
end rtl;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;

entity PipelinedFPOperator is
  generic (
      name : string;
      operator_id : string;
      exponent_width : integer := 8;
      fraction_width : integer := 23;
      no_arbitration: boolean := true;
      num_reqs : integer := 3; -- how many requesters?
      use_input_buffering: boolean := true;
      detailed_buffering_per_input: IntegerArray;
      detailed_buffering_per_output: IntegerArray;
      full_rate: boolean
    );
  port (
    -- req/ack follow level protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackR                     : out BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    reqR                     : in  BooleanArray(num_reqs-1 downto 0);
    -- input data consists of concatenated pairs of ips
    dataL                    : in std_logic_vector((2*(exponent_width+fraction_width+1)*num_reqs)-1 downto 0);
    -- output data consists of concatenated pairs of ops.
    dataR                    : out std_logic_vector(((exponent_width+fraction_width+1)*num_reqs)-1 downto 0);
    -- with dataR
    clk, reset              : in std_logic);
end PipelinedFPOperator;

architecture Vanilla of PipelinedFPOperator is

  constant num_operands : integer := 2;
  constant operand_width : integer := exponent_width+fraction_width+1;
  constant iwidth : integer := 2*operand_width;
  constant owidth : integer := operand_width;
  
  constant tag_length: integer := Maximum(1,Ceil_Log2(reqL'length));
  signal itag,otag : std_logic_vector(tag_length-1 downto 0);
  signal ireq,iack, oreq, oack: std_logic;

  constant debug_flag : boolean := global_debug_flag;

  signal idata: std_logic_vector(iwidth-1 downto 0);
  signal odata: std_logic_vector(owidth-1 downto 0);

  signal NaN, overflow, underflow : std_logic;
  constant use_as_subtractor : boolean := (operator_id = "ApFloatSub");


  -----------------------------------------------------------------------------
  -- for the moment..
  constant use_generic_multiplier : boolean := true;
  -----------------------------------------------------------------------------
  
begin  -- Behave
  assert ackL'length = reqL'length report "mismatched req/ack vectors" severity error;
  assert ((operand_width = 32) or (operand_width = 64)) report "32/64 bit operand-support only!" severity error;
  assert ((operator_id = "ApFloatMul") or (operator_id = "ApFloatAdd") or (operator_id = "ApFloatSub"))
    report "operator_id must be either add or mul or sub" severity error;  

  -- DebugGen: if debug_flag generate 
    -- assert( (not ((reset = '0') and (clk'event and clk = '1') and no_arbitration)) or Is_At_Most_One_Hot(reqL))
    -- report "in no-arbitration case, at most one request should be hot on clock edge (in SplitOperatorShared)" severity error;
  -- end generate DebugGen;
  NoInBuffers : if not use_input_buffering generate 
    imux: InputMuxBase
      generic map(name => name & "-imux",
		  iwidth => iwidth*num_reqs,
                  owidth => iwidth, 
                  twidth => tag_length,
                  nreqs => num_reqs,
                  no_arbitration => no_arbitration,
                  registered_output => false)
      port map(
          reqL       => reqL,
        ackL       => ackL,
        reqR       => ireq,
        ackR       => iack,
        dataL      => dataL,
        dataR      => idata,
        tagR       => itag,
        clk        => clk,
        reset      => reset);
   end generate NoInBuffers;

  InBuffers: if use_input_buffering generate
    imuxWithInputBuf: InputMuxWithBuffering
      generic map(name => name & "-imux" , 
		iwidth => iwidth*num_reqs,
                owidth => iwidth, 
                twidth => tag_length,
                nreqs => num_reqs,
		buffering => detailed_buffering_per_input,
                no_arbitration => no_arbitration,
		full_rate => full_rate,
                registered_output => false)
      port map(
        reqL       => reqL,
        ackL       => ackL,
        reqR       => ireq,
        ackR       => iack,
        dataL      => dataL,
        dataR      => idata,
        tagR       => itag,
        clk        => clk,
        reset      => reset);
  end generate InBuffers;

  IEEE754xMul:  if operator_id = "ApFloatMul" generate
    useGeneric: if use_generic_multiplier generate
    op: GenericFloatingPointMultiplier
      generic map(name => name & "-IEEE754-mul", tag_width     => tag_length,
                   exponent_width => exponent_width,
                   fraction_width => fraction_width,
                   round_style => round_nearest,
                   addguard => 3,
                   check_error => true,
                   denormalize => true)
      port map (
        env_rdy => ireq,
        muli_rdy => iack,
        accept_rdy => oack,
        mulo_rdy => oreq,
        INA => idata((2*operand_width)-1 downto operand_width),
        INB => idata(operand_width-1 downto 0),
        OUTMUL => odata,
        tag_in => itag,
        tag_out => otag,
        clk => clk,
        reset => reset);
    end generate useGeneric;
    
    SinglePrecision: if operand_width = 32 and (not use_generic_multiplier) generate 
    	op: SinglePrecisionMultiplier
          generic map(name => name & "-SinglePrecision-op",
					 tag_width     => tag_length)
          port map (
            env_rdy => ireq,
            muli_rdy => iack,
            accept_rdy => oack,
            mulo_rdy => oreq,
            INA => idata(63 downto 32),
            INB => idata(31 downto 0),
            OUTM => odata,
            tag_in => itag,
            tag_out => otag,
            NaN => NaN,
            oflow => overflow,
            uflow => underflow,
            clk => clk,
            reset => reset);
	end generate SinglePrecision;


    DoublePrecision: if operand_width = 64 and (not use_generic_multiplier) generate 
    	op: DoublePrecisionMultiplier
          generic map ( name => name & "-DoublePrecision-op",
					tag_width     => tag_length)
          port map (
            env_rdy => ireq,
            muli_rdy => iack,
            accept_rdy => oack,
            mulo_rdy => oreq,
            INA => idata(127 downto 64),
            INB => idata(63 downto 0),
            OUTM => odata,
            tag_in => itag,
            tag_out => otag,
            NaN => NaN,
            oflow => overflow,
            uflow => underflow,
            clk => clk,
            reset => reset);
    end generate DoublePrecision;
  end generate IEEE754xMul;

  IEEE754xAdd:  if ((operator_id = "ApFloatAdd") or (operator_id = "ApFloatSub")) generate
    op: GenericFloatingPointAdderSubtractor
      generic map(name => name & "-IEEE754-add", tag_width     => tag_length,
                   exponent_width => exponent_width,
                   fraction_width => fraction_width,
                   round_style => round_nearest,
                   addguard => 3,
                   check_error => true,
                   denormalize => true,
                   use_as_subtractor => use_as_subtractor)
      port map (
        env_rdy => ireq,
        addi_rdy => iack,
        accept_rdy => oack,
        addo_rdy => oreq,
        INA => idata((2*operand_width)-1 downto operand_width),
        INB => idata(operand_width-1 downto 0),
        OUTADD => odata,
        tag_in => itag,
        tag_out => otag,
        clk => clk,
        reset => reset);
  end generate IEEE754xAdd;


  odemux: OutputDeMuxBaseWithBuffering
    generic map (
        name => name & "-odemux",
  	iwidth => owidth,
  	owidth =>  owidth*num_reqs,
	twidth =>  tag_length,
	nreqs  => num_reqs,
	detailed_buffering_per_output => detailed_buffering_per_output,
	full_rate => full_rate)
    port map (
      reqL   => oreq,
      ackL   => oack,
      dataL => odata,
      tagL  => otag,
      reqR  => reqR,
      ackR  => ackR,
      dataR => dataR,
      clk   => clk,
      reset => reset);
  
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Authors: Abhishek R. Kamath & Prashant Singhal
-- An IEEE-754 compliant Single-Precision pipelined multiplier
--
--   rounding-scheme implemented is round-to-zero.
--   overflow/underflow exceptions are detected.
--
--   TODO: implement round-to-nearest since this
--         is preferred to reduce errors.
-- 
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity SinglePrecisionMultiplier is
  generic (name: string; tag_width : integer);
  port(
    INA, INB: in std_logic_vector(31 downto 0);
    OUTM: out std_logic_vector(31 downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    NaN, oflow, uflow: out std_logic := '0';
    env_rdy, accept_rdy: in std_logic;
    muli_rdy, mulo_rdy: out std_logic);
end entity;

architecture rtl of SinglePrecisionMultiplier is

  type parpro is array (0 to 23) of std_logic_vector(23 downto 0);


  signal rdy1,rdy2,rdy3,rdy4,rdy5,rdy6,rdy7,rdy8,rdy9,rdy10, rdy11: std_logic := '0';
  signal flag3,flag4,flag5,flag6,flag7,flag8,flag9,flag10: std_logic_vector(1 downto 0);
  signal fman10: std_logic_vector(22 downto 0);
  signal tag1,tag2,tag3,tag4,tag5,tag6,tag7,tag8,tag9,tag10: std_logic_vector(tag_width-1 downto 0);
  signal pipeline_stall: std_logic := '0';

  signal aman_1,aman_2,bman_1,bman_2: std_logic_vector(23 downto 0);
  signal anan1,bnan1,azero1,bzero1,ainf1,binf1,osgn1: std_logic := '0'; 
  signal aexp_s1,bexp_s1: std_logic_vector(7 downto 0);

  signal nocalc2,nocalc3,nocalc4,nocalc5,nocalc6,nocalc7,nocalc8,nocalc9,nocalc10: std_logic;-- := '0';
  signal output_s2,output_s23,output_s24,output_s25,output_s26,output_s27,output_s28,output_s29,output_s210: std_logic_vector(2 downto 0);
  signal int_exp: std_logic_vector(8 downto 0);

  signal fexp3,fexp4,fexp5,fexp6,fexp7,fexp8,fexp9,fexp10: std_logic_vector(7 downto 0);-- := X"00";

  signal pp: parpro;
  signal tr_400,tr_401,tr_402,tr_403,tr_404,tr_405,tr_406,tr_407,tr_408,tr_409,tr_410,tr_411: std_logic_vector(47 downto 0);

  signal tr51,tr52,tr53,tr54,tr55,tr56,tr61,tr62,tr63,tr7,tr_temp,tr9: std_logic_vector(47 downto 0);

  signal tr401,tr402,tr403,tr404,tr405,tr406,tr407,tr408,tr409,tr410,tr411,tr412: std_logic_vector(47 downto 0);-- := X"000000000000";
  signal tr413,tr414,tr415,tr416,tr417,tr418,tr419,tr420,tr421,tr422,tr423,tr424: std_logic_vector(47 downto 0);-- := X"000000000000";

begin

  stage_1: process(clk,reset)

    variable asgn,bsgn,osgn: std_logic := '0';
    variable aexp,bexp: std_logic_vector(7 downto 0);-- := X"00";
    variable aman,bman: std_logic_vector(23 downto 0);-- := "000000000000000000000000";
    variable anan,bnan,azero,bzero,ainf,binf: std_logic;-- := '0';

  begin
    if reset = '1' then
      rdy1 <= '0';
    else
      if clk'event and clk='1'then
	if env_rdy = '1' and pipeline_stall = '0' then

          aexp := INA(30 downto 23);
          bexp := INB(30 downto 23);
          aman := '1' & INA(22 downto 0);
          bman := '1' & INB(22 downto 0);

          if(aexp=X"FF") then
            if(unsigned(aman)=0) then
              ainf := '1';
              anan := '0';
              azero := '0';
            else
              anan := '1';
              azero := '0';
              ainf := '0';
            end if;
          elsif(aexp=X"00") then
            if unsigned(aman)=0 then
              azero := '1';
              ainf := '0';
              anan := '0';
            end if;
          else
            ainf := '0';
            anan := '0';
            azero := '0';
          end if;

          if(bexp=X"FF") then
            if(unsigned(bman)=0) then
              binf := '1';
              bnan := '0';
              bzero := '0';
            else
              bnan := '1';
              bzero := '0';
              binf := '0';
            end if;
          elsif(bexp=X"00") then
            if unsigned(bman)=0 then
              bzero := '1';
              binf := '0';
              bnan := '0';
            end if;
          else
            binf := '0';
            bnan := '0';
            bzero := '0';
          end if;

          osgn1 <= INA(31) xor INB(31);

          ainf1 <= ainf;
          binf1 <= binf;
          anan1 <= anan;
          bnan1 <= bnan;
          azero1 <= azero;
          bzero1 <= bzero;

          aexp_s1 <= aexp;
          bexp_s1 <= bexp;
          aman_1 <= aman;
          bman_1 <= bman;


          rdy1 <= '1';
          tag1 <= tag_in;

        elsif pipeline_stall = '1' then
        elsif env_rdy = '0' then
          rdy1 <= '0';
        end if;
      end if;
    end if;
  end process stage_1;





  stage_2: process(clk,reset)
  begin
    if reset = '1' then
      rdy2 <= '0';
    else
      if clk'event and clk='1'then
	if rdy1 = '1' and pipeline_stall = '0' then
          if (anan1 = '1' or bnan1 = '1') then
            output_s2 <= osgn1 & "10";
            nocalc2 <= '1';
          elsif (azero1 = '1' and binf1 = '1') or (ainf1 = '1' and bzero1 = '1') then
            output_s2 <= osgn1 & "10";
            nocalc2 <= '1';
          elsif azero1 = '1' or bzero1 = '1' then
            output_s2 <= osgn1 & "00";
            nocalc2 <= '1';
          elsif ainf1 = '1' or binf1 = '1' then
            output_s2 <= osgn1 & "11";
            nocalc2 <= '1';
          else
            int_exp <= std_logic_vector(unsigned('0' & aexp_s1) + unsigned('0' & bexp_s1));
            output_s2 <= osgn1 & "01";
            nocalc2 <= '0';
          end if;
          aman_2 <= aman_1;
          bman_2 <= bman_1;
          rdy2 <= '1';
          tag2 <= tag1;


	elsif pipeline_stall = '1' then
	elsif rdy1 = '0' then
          rdy2 <= '0';
	end if;
      end if;
    end if;
  end process stage_2;




  stage_3: process(clk,reset)

    variable exp3: unsigned(8 downto 0);

  begin
    if reset = '1' then
      rdy3 <= '0';
    else
      if clk'event and clk='1'then
	if rdy2 = '1' and pipeline_stall = '0' then
          if nocalc2 = '1' then
            nocalc3 <= '1';
            output_s23 <= output_s2;
            flag3 <= "00";
          elsif nocalc2 = '0' then
            exp3 := unsigned(int_exp);
            if(exp3 > 381) then
              output_s23 <= output_s2(2) & "11";
              nocalc3 <= '1';
              flag3 <= "10";
            elsif(exp3 < 127) then
              output_s23 <= output_s2(2) & "00";
              nocalc3 <= '1';
              flag3 <= "01";
            else
              exp3 := exp3 - 127;
              output_s23 <= output_s2(2) & "01";
              nocalc3 <= '0';
              flag3 <= "00";
            end if;	
          end if;
          fexp3 <= std_logic_vector(exp3(7 downto 0));
          rdy3 <= '1';
          tag3 <= tag2;

          for i in 0 to 23 loop
            for j in 0 to 23 loop
              pp(i)(j) <= aman_2(j) and bman_2(i);
            end loop;
          end loop;

	elsif pipeline_stall = '1' then
	elsif rdy2 = '0' then
          rdy3 <= '0';
	end if;
      end if;
    end if;
  end process stage_3;





  stage_4: process(clk,reset)
  begin
    if reset = '1' then
      rdy4 <= '0';
    else
      if clk'event and clk='1'then
	if rdy3 = '1' and pipeline_stall = '0' then
          if nocalc3 = '1' then
            nocalc4 <= '1';
          elsif nocalc3 = '0' then

            tr401 <= X"000000" & pp(0);
            tr402 <= X"00000" & "000" & pp(1) & '0';
            tr403 <= X"00000" & "00" & pp(2) & "00";
            tr404 <= X"00000" & '0' & pp(3) & "000";	

            tr405 <= X"00000" & pp(4) & X"0";
            tr406 <= X"0000" & "000" & pp(5) & X"0" & '0';
            tr407 <= X"0000" & "00" & pp(6) & X"0" & "00";
            tr408 <= X"0000" & '0' & pp(7) & X"0" & "000";

            tr409 <= X"0000" & pp(8) & X"00";
            tr410 <= X"000" & "000" & pp(9) & X"00" & '0';
            tr411 <= X"000" & "00" & pp(10) & X"00" & "00";
            tr412 <= X"000" & '0' & pp(11) & X"00" & "000";

            tr413 <= X"000" & pp(12) & X"000";
            tr414 <= X"00" & "000" & pp(13) & X"000" & '0';
            tr415 <= X"00" & "00" & pp(14) & X"000" & "00";
            tr416 <= X"00" & '0' & pp(15) & X"000" & "000";

            tr417 <= X"00" & pp(16) & X"0000";
            tr418 <= X"0" & "000" & pp(17) & X"0000" & '0';
            tr419 <= X"0" & "00" & pp(18) & X"0000" & "00";
            tr420 <= X"0" & '0' & pp(19) & X"0000" & "000";

            tr421 <= X"0" & pp(20) & X"00000";
            tr422 <= "000" & pp(21) & X"00000" & '0';
            tr423 <= "00" & pp(22) & X"00000" & "00";
            tr424 <= '0' & pp(23) & X"00000" & "000";

            nocalc4 <= '0';

          end if;


          output_s24 <= output_s23;
          fexp4 <= fexp3;
          flag4 <= flag3;
          rdy4 <= '1';
          tag4 <= tag3;

	elsif pipeline_stall = '1' then
	elsif rdy3 = '0' then
          rdy4 <= '0';
	end if;
      end if;
    end if;
  end process stage_4;


  stage_5: process(clk,reset)
  begin
    if reset = '1' then
      rdy5 <= '0';
    else
      if clk'event and clk='1'then
	if rdy4 = '1' and pipeline_stall = '0' then
          if nocalc4 = '1' then
            nocalc5 <= '1';
          elsif nocalc4 = '0' then

            tr_400 <= std_logic_vector(unsigned(tr401) + unsigned(tr402));
            tr_401 <= std_logic_vector(unsigned(tr403) + unsigned(tr404));
            tr_402 <= std_logic_vector(unsigned(tr405) + unsigned(tr406));
            tr_403 <= std_logic_vector(unsigned(tr407) + unsigned(tr408));
            tr_404 <= std_logic_vector(unsigned(tr409) + unsigned(tr410));
            tr_405 <= std_logic_vector(unsigned(tr411) + unsigned(tr412));
            tr_406 <= std_logic_vector(unsigned(tr413) + unsigned(tr414));
            tr_407 <= std_logic_vector(unsigned(tr415) + unsigned(tr416));
            tr_408 <= std_logic_vector(unsigned(tr417) + unsigned(tr418));
            tr_409 <= std_logic_vector(unsigned(tr419) + unsigned(tr420));
            tr_410 <= std_logic_vector(unsigned(tr421) + unsigned(tr422));
            tr_411 <= std_logic_vector(unsigned(tr423) + unsigned(tr424));

            nocalc5 <= '0';

          end if;


          output_s25 <= output_s24;
          fexp5 <= fexp4;
          flag5 <= flag4;
          rdy5 <= '1';
          tag5 <= tag4;

	elsif pipeline_stall = '1' then
	elsif rdy4 = '0' then
          rdy5 <= '0';
	end if;
      end if;
    end if;
  end process stage_5;



  stage_6: process(clk,reset)
  begin
    if reset = '1' then
      rdy6 <= '0';
    else
      if clk'event and clk='1'then
	if rdy5 = '1' and pipeline_stall = '0' then
          if nocalc5 = '1' then
            nocalc6 <= '1';
          else
            tr51 <= std_logic_vector(unsigned(tr_400) + unsigned(tr_401));
            tr52 <= std_logic_vector(unsigned(tr_402) + unsigned(tr_403));
            tr53 <= std_logic_vector(unsigned(tr_404) + unsigned(tr_405));
            tr54 <= std_logic_vector(unsigned(tr_406) + unsigned(tr_407));
            tr55 <= std_logic_vector(unsigned(tr_408) + unsigned(tr_409));
            tr56 <= std_logic_vector(unsigned(tr_410) + unsigned(tr_411));
            nocalc6 <= '0';
          end if;

          output_s26 <= output_s25;
          fexp6 <= fexp5;
          flag6 <= flag5;
          rdy6 <= '1';
          tag6 <= tag5;

	elsif pipeline_stall = '1' then
	elsif rdy5 = '0' then
          rdy6 <= '0';
	end if;
      end if;
    end if;
  end process stage_6;



  stage_7: process(clk,reset)
  begin
    if reset = '1' then
      rdy7 <= '0';
    else
      if clk'event and clk='1'then
	if rdy6 = '1' and pipeline_stall = '0' then
          if nocalc6 = '1' then
            nocalc7 <= '1';
          else
            tr61 <= std_logic_vector(unsigned(tr51) + unsigned(tr52));
            tr62 <= std_logic_vector(unsigned(tr53) + unsigned(tr54));
            tr63 <= std_logic_vector(unsigned(tr55) + unsigned(tr56));
            nocalc7 <= '0';
          end if;

          output_s27 <= output_s26;
          fexp7 <= fexp6;
          flag7 <= flag6;
          rdy7 <= '1';
          tag7 <= tag6;

	elsif pipeline_stall = '1' then
	elsif rdy6 = '0' then
          rdy7 <= '0';
	end if;
      end if;
    end if;
  end process stage_7;

  stage_8: process(clk,reset)
  begin
    if reset = '1' then
      rdy8 <= '0';
    else
      if clk'event and clk='1'then
	if rdy7 = '1' and pipeline_stall = '0' then
          if nocalc7 = '1' then
            nocalc8 <= '1';
          else
            tr7 <= std_logic_vector(unsigned(tr61) + unsigned(tr62));
            nocalc8 <= '0';
          end if;

          output_s28<= output_s27;
          fexp8 <= fexp7;
          flag8 <= flag7;
          rdy8 <= '1';
          tag8 <= tag7;
          tr_temp <= tr63;

	elsif pipeline_stall = '1' then
	elsif rdy7 = '0' then
          rdy8 <= '0';
	end if;
      end if;
    end if;
  end process stage_8;

  stage_9: process(clk,reset)
  begin
    if reset = '1' then
      rdy9 <= '0';
    else
      if clk'event and clk='1'then
	if rdy8 = '1' and pipeline_stall = '0' then
          if nocalc8 = '1' then
            nocalc9 <= '1';
          else
            tr9 <= std_logic_vector(unsigned(tr7) + unsigned(tr_temp));
            nocalc9 <= '0';
          end if;

          output_s29 <= output_s28;
          fexp9 <= fexp8;
          flag9 <= flag8;
          rdy9 <= '1';
          tag9 <= tag8;

	elsif pipeline_stall = '1' then
	elsif rdy8 = '0' then
          rdy9 <= '0';
	end if;
      end if;
    end if;
  end process stage_9;


  stage_10: process(clk,reset)
    variable man8: std_logic_vector(24 downto 0);
    variable exp8: unsigned(7 downto 0);
  begin
    if reset = '1' then
      rdy10 <= '0';
    else
      if clk'event and clk='1'then
	if rdy9 = '1' and pipeline_stall = '0' then
          if nocalc9 = '1' then
            nocalc10 <= '1';
            output_s210 <= output_s29;
            flag10 <= flag9;
          elsif nocalc9 = '0' then
            man8 := tr9(47 downto 23);
            exp8 := unsigned(fexp9);
            if man8(24) = '1' then
              if	exp8 = 254 then
                output_s210 <= output_s29(2) & "11";
                nocalc10 <= '1';
                flag10 <= "10";
              else
                exp8 := exp8 + 1;
                nocalc10 <= '0';
                fman10 <= man8(23 downto 1);
                output_s210 <= output_s29;
                flag10 <= flag9;
              end if;
            elsif exp8 = 0 then
              output_s210 <= output_s29(2) & "00";
              nocalc10 <= '1';
              flag10 <= "01";
            else
              fman10 <= man8(22 downto 0);
              output_s210 <= output_s29;
              nocalc10 <= '0';
              flag10 <= flag9;
            end if;
          end if;		
          rdy10 <= '1';
          tag10 <= tag9;
          fexp10 <= std_logic_vector(exp8);
        elsif pipeline_stall = '1' then
        elsif rdy9 = '0' then
          rdy10 <= '0';
        end if;
      end if;
    end if;
  end process stage_10;


  stage_11: process(clk,reset)
    variable temp: std_logic_vector(2 downto 0);
  begin
    if reset = '1' then
      rdy11 <= '0';
    else
      if clk'event and clk='1'then
	if rdy10 = '1' and pipeline_stall = '0' then
          rdy11 <= '1';
          temp := output_s210;
          if nocalc10 = '1' then
            case(temp(1 downto 0)) is
              when("00") => OUTM <= temp(2) & "000" & X"0000000"; NaN <= '0'; oflow <= '0'; uflow <= flag10(0);
            when("10") => OUTM <= temp(2) & X"FF" & "10000000000000000000000"; NaN <= '1'; oflow <= '0'; uflow <= '0';
            when("11") => OUTM <= temp(2) & X"FF" & "000" & X"00000"; NaN <= '0'; oflow <= flag10(1); uflow <= '0';
            when others => null; 
          end case;
          else
            OUTM <= temp(2) & fexp10 & fman10; NaN <= '0'; oflow <='0'; uflow <= '0';
          end if;
          tag_out <= tag10;
        else
          rdy11 <= '0';
        end if;
      end if;
    end if;
  end process stage_11;

  pipeline_stall <= (rdy11 and (not accept_rdy));
  muli_rdy <= not (rdy11 and (not accept_rdy));
  mulo_rdy <= rdy11;

end rtl;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- a basic unsigned adder..  if addition is specified, just
-- adds using a simple carry lookahead scheme.  if subtraction
-- is specified, takes the twos complement of the second operand
-- and adds the two numbers.  No overflow/negative checks
-- are performed.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;

entity AddSubCell  is
	generic ( operand_width: integer);
	port (A,B: in unsigned(operand_width-1 downto 0);
		Sum: out unsigned(operand_width-1 downto 0);
		BP,BG: out std_logic;
		stall: in std_logic;
		clk, reset: in std_logic);
end entity AddSubCell;

architecture Behave of AddSubCell is
begin
	process(clk, reset, A, B, stall)
		variable sumv: unsigned(operand_width-1 downto 0);
		variable prop, gen: std_logic;
	begin
		prop := '1';
		gen  := '0';

		sumv := A+B;

		for I in 0 to operand_width-1 loop
			prop := (prop and (A(I) or B(I)));
			gen  := (A(I) and B(I)) or (gen and (A(I) or B(I)));
		end loop;


		if(clk'event and clk = '1') then
		   if(stall = '0') then
			Sum <= sumv;
			BP <= prop;
			BG <= gen;
		   end if;
		end if;
	end process;
end Behave;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
entity UnsignedAdderSubtractor is
  
  generic (
    name: string;
    tag_width          : integer;
    operand_width      : integer;
    chunk_width        : integer
	);

  port (
    L            : in  unsigned(operand_width-1 downto 0);
    R            : in  unsigned(operand_width-1 downto 0);
    RESULT       : out unsigned(operand_width-1 downto 0);
    subtract_op  : in std_logic;
    clk, reset   : in  std_logic;
    in_rdy       : in  std_logic;
    out_rdy      : out std_logic;
    stall        : in std_logic;
    tag_in       : in std_logic_vector(tag_width-1 downto 0);
    tag_out      : out std_logic_vector(tag_width-1 downto 0));
end entity;


architecture Pipelined of UnsignedAdderSubtractor is
 
  constant num_chunks: integer := Ceil(operand_width, chunk_width);
  constant padded_operand_width: integer := num_chunks  * chunk_width;
  signal Lpadded, Rpadded, Resultpadded : unsigned(padded_operand_width-1 downto 0);

  constant pipe_depth : integer := 3;
  signal stage_active : std_logic_vector(0 to pipe_depth);


  type CWORD is array (natural range <>) of unsigned(chunk_width-1 downto 0);
  type TWORD is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);  
  signal stage_tags: TWORD(0 to pipe_depth);


  signal addsubcell_Sum, addsubcell_Sum_Delayed, 
			addsubcell_A, addsubcell_B, final_sums: CWord(0 to num_chunks-1);
  signal addsubcell_BP, addsubcell_BG : std_logic_vector(0 to num_chunks-1);
  signal addsubcell_Cin: std_logic_vector(0 to num_chunks);
  constant zero_Cin: std_logic_vector(0 to num_chunks) := (others => '0');


  signal block_carries: std_logic_vector(0 to num_chunks);
  signal subtract_op_1, subtract_op_2: std_logic;


  component AddSubCell  is
	generic ( operand_width: integer);
	port (A,B: in unsigned(operand_width-1 downto 0);
		Sum: out unsigned(operand_width-1 downto 0);
		BP,BG: out std_logic;
		stall: in std_logic;
		clk, reset: in std_logic);
  end component AddSubCell;
  
begin  -- Pipelined

  -- note: if subtract_op = '1', then complement R (see below) and add 1.
  process(subtract_op)
     variable TMP: std_logic_vector(0 to num_chunks);
  begin
     TMP := (others =>  '0');
     if (subtract_op = '1') then
       TMP(0) := '1';
     end if;
     addsubcell_Cin <= TMP;
  end process;

  stage_active(0) <= in_rdy;
  out_rdy <= stage_active(pipe_depth);
  stage_tags(0) <= tag_in;
  tag_out <= stage_tags(3);

  RESULT <= Resultpadded(operand_width-1 downto 0);


  -- pad. also if subtract_op = '1' then complement R and add 1 (addsubcell_Cin).
  process(L,R,subtract_op)
	variable ltmp, rtmp: unsigned(padded_operand_width-1 downto 0);
  begin
	ltmp := (others => '0'); ltmp(operand_width-1 downto 0) := L;
	rtmp := (others => '0'); rtmp(operand_width-1 downto 0) := R;
	Lpadded <= ltmp;

	if(subtract_op = '0') then
		Rpadded <= rtmp;
	else
		Rpadded <= not rtmp;
	end if;
  end process;

  Stage1:  for I in  0 to num_chunks-1 generate

	addsubCell_A(I) <= Lpadded(((I+1)*chunk_width)-1 downto (I*chunk_width));
	addsubCell_B(I) <= Rpadded(((I+1)*chunk_width)-1 downto (I*chunk_width));

	asCell: AddSubCell generic map(operand_width => chunk_width)
		port  map( A => addsubcell_A(I),
			   B => addsubcell_B(I),	
			   Sum => addsubcell_Sum(I),
			   BP => addsubcell_BP(I),
			   BG => addsubcell_BG(I),
			   stall => stall,
			   clk => clk,
			   reset => reset);
  end generate Stage1;

  process(clk)
  begin
	if(clk'event and clk = '1') then
		if(stall = '0') then
			stage_tags(1) <= stage_tags(0);
			subtract_op_1 <= subtract_op;
		end if;
		if(reset = '1') then
			stage_active(1) <= '0';
		elsif stall = '0' then
			stage_active(1) <= stage_active(0);
		end if;
	end if;
  end process;

  -- stage two: calculate the block carries.
  MoreThanOneChunk: if (num_chunks > 1) generate
     process(clk, reset, stall, stage_active, addsubcell_Cin, addsubcell_BP, addsubcell_BG)	
	variable cin: std_logic_vector(0 to num_chunks);
     begin
	cin := addsubcell_Cin;
	for I in 1 to num_chunks loop
		cin(I) := (cin(I-1) and addsubcell_BP(I-1))  or addsubcell_BG(I-1);
	end loop;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			stage_active(2) <= '0';
		elsif(stall = '0') then
			block_carries <= cin;
			stage_tags(2) <= stage_tags(1);
			addsubcell_Sum_Delayed <= addsubcell_Sum;
			subtract_op_2 <= subtract_op_1;
			stage_active(2) <= stage_active(1);
		end if;
	end if;
    end process;




  -- stage three: final sums
    process(clk)
	variable correction, tmp: unsigned(chunk_width-1 downto 0);
	variable is_negative: boolean;
    begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			stage_active(3) <= '0';
		elsif(stall = '0') then
			final_sums(0) <= addsubcell_Sum_Delayed(0);
			for I in 0 to num_chunks-1 loop
				correction := (others => '0');
				if(block_carries(I) = '1') then
					correction(0) := '1';
				end if;
				final_sums(I) <= addsubcell_Sum_Delayed(I) + correction;
			end loop;

			stage_tags(3) <= stage_tags(2);
			stage_active(3) <= stage_active(2);
		end if;
	end if;
    end process;

  end generate MoreThanOneChunk;

  OnlyOneChunk: if (num_chunks = 1) generate
     stage_tags(2) <= stage_tags(1);
     stage_active(2) <= stage_active(1);
     addsubcell_Sum_Delayed <= addsubcell_Sum;

     stage_tags(3) <= stage_tags(2);
     stage_active(3) <= stage_active(2);
     final_sums(0) <= addsubcell_Sum_Delayed(0) when (subtract_op = '0') else (addsubcell_Sum_Delayed(0) + 1);

  end generate OnlyOneChunk;

  -- collect final-sums into RESULT
  process(final_sums)
  begin
	for I in 0 to num_chunks-1 loop
		ResultPadded(((I+1)*chunk_width)-1 downto (I*chunk_width)) <= final_sums(I);
	end loop;
  end process;

end Pipelined;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- a basic unsigned multiplier.
--
-- for the moment, this just does a multiply and adds delay stages at
-- the end; presumably, the synthesis tool will retime things
-- appropriately..
--
-- TODO: pipeline this explicitly!
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity DelayCell is
   generic (operand_width: integer; delay: natural);
   port (Din: in unsigned(operand_width-1 downto 0);
	 Dout: out unsigned(operand_width-1 downto 0);
	 clk: in std_logic;
	 stall: in std_logic);
end entity DelayCell;

architecture Behave of DelayCell is
	type DArray is array (natural range <>) of unsigned(operand_width-1 downto 0);
	signal data_array: DArray(0 to delay);
begin

	data_array(0) <= Din;
	NonZeroDelay: if delay > 0 generate
	   SRgen: for I in 1 to delay generate
		process(clk)
		begin
			if(clk'event and clk = '1') then
				if(stall = '0') then
					data_array(I) <= data_array(I-1);
				end if;
			end if;
			
		end process;
	    end generate SRgen;
	end generate NonZeroDelay;
	
	Dout <= data_array(delay);
end Behave;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SumCell is
 	generic (operand_width: integer; ignore_diag: boolean; ignore_right: boolean);
	port (SU,SDiagIn: in unsigned(operand_width-1 downto 0);
              SR: in unsigned(1 downto 0);
	      SDiagOut: out unsigned(operand_width-1 downto 0);
	      SL: out unsigned(1 downto 0);
	      stall: in std_logic;
	      clk: in std_logic);
end entity SumCell;

architecture Behave of SumCell is
begin

	process(clk)
		variable x, y, z, sum: unsigned(operand_width+1 downto 0);
		variable t: unsigned(1 downto 0);
	begin

		if(clk'event and clk = '1') then
                        y := (others => '0');
			if(stall = '0') then
				x := "00" & SU;

				-- y := (1 => SR(1), 0 => SR(0), others => '0');
                                y(1) := SR(1);
                                y(0) := SR(0);

				z := "00" & SDiagIn;
		
				if(not (ignore_diag  or ignore_right)) then
					sum := x + y + z;
				elsif (ignore_diag and ignore_right) then
					sum := x;
				elsif (ignore_diag and (not ignore_right)) then
					sum := (x + y);
				else
					sum := (x + z);
				end if;
	
				t := sum(operand_width+1 downto operand_width);

				SDiagOut <= sum(operand_width-1 downto 0);
				SL <= t;
			end if;
		end if;
	end process;
end Behave;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MultiplierCell is
  generic (operand_width: integer);
  port (MT, MR, ST, DiagIn: in unsigned(operand_width-1 downto 0);
        ML, MD, SD, DiagOut: out unsigned(operand_width-1 downto 0);
        stall: in std_logic;
	clk: in std_logic);
end entity MultiplierCell;

architecture Simple of MultiplierCell is
	constant zero_const : unsigned(operand_width-2 downto 0) := (others => '0');
begin

	-- sent through without any delay.
	ML <= MR;

	process(clk)
		variable tmp,wext: unsigned((2*operand_width)-1 downto 0);
		variable u, v, w: unsigned(operand_width downto 0);
	begin
		if(clk'event and clk = '1') then
			if(stall = '0') then
				tmp := MT*MR;
		
				-- pad one bit to incoming summands.
				u :=  "0" & DiagIn;
                                v :=  "0" & ST;
		
				-- this is a operand_width+1 size addition
				w := (u + v);

				-- pad to 2*operand_width
				wext := zero_const & w;
		
				-- a full 2*operand_width addition.
				tmp := tmp + wext;

				-- send down the vertical operand
				-- with a cycle delay.
				MD <= MT;

				-- top half of result goes down to 
				-- next row (to be summed)
				SD <= tmp((2*operand_width)-1 downto operand_width);

				-- bottom half of the result goes out
				-- on the diagonal..
				DiagOut <= tmp(operand_width-1 downto 0);
			end if;
		end if;
	end process;
end Simple;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;

entity UnsignedMultiplier is
  
  generic (
    name: string;
    tag_width     : integer;
    operand_width : integer;
    chunk_width   : integer := 8);

  port (
    L, R       : in  unsigned(operand_width-1 downto 0);
    RESULT     : out unsigned((2*operand_width)-1 downto 0);
    clk, reset : in  std_logic;
    in_rdy     : in  std_logic;
    out_rdy    : out std_logic;
    stall      : in std_logic;
    tag_in     : in std_logic_vector(tag_width-1 downto 0);
    tag_out    : out std_logic_vector(tag_width-1 downto 0));
end entity;

architecture Pipelined of UnsignedMultiplier is

  constant pipe_depth : integer := operand_width/16;

  type RWORD is array (natural range <>) of unsigned((2*operand_width)-1 downto 0);
  type TWORD is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);  


  signal intermediate_results : RWORD(0 to pipe_depth);
  signal intermediate_tags : TWORD(0 to pipe_depth);  
  signal stage_active : std_logic_vector(0 to pipe_depth);
  
begin  -- Pipelined

  -- for now, just multiply..
  intermediate_results(0) <= L*R;


  -- I/O
  intermediate_tags(0) <= tag_in;
  stage_active(0) <= in_rdy;
  out_rdy <= stage_active(pipe_depth);
  tag_out <= intermediate_tags(pipe_depth);
  RESULT <= intermediate_results(pipe_depth);
  
  -- for now, just add stages after the multiply
  -- the synthesis tool should retime.  Later
  -- we'll get around to doing the array multiplier
  -- right.
  Pipeline: for STAGE in 1 to pipe_depth generate

    process(clk)
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          stage_active(STAGE) <= '0';
        elsif(stall = '0') then
          stage_active(STAGE) <= stage_active(STAGE-1);
        end if;

        if(stall = '0') then
          intermediate_results(STAGE) <= intermediate_results(STAGE-1);
          intermediate_tags(STAGE) <= intermediate_tags(STAGE-1);
        end if;
        
      end if;
    end process;
    
  end generate Pipeline;
end Pipelined;


 
architecture ArrayMul of UnsignedMultiplier is

	constant NumChunks : integer := Ceil(operand_width, chunk_width);

	constant padded_operand_width: integer  := NumChunks*chunk_width;
	signal Lpadded, Rpadded: unsigned(padded_operand_width-1 downto 0);
	signal RESULTpadded: unsigned((2*padded_operand_width)-1 downto 0);

	type TwoDTagArray is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);
	signal tag_array: TwoDTagArray(0 to 2*NumChunks);

	type TwoDChunkArray is array (natural range <>, natural range <>) of unsigned(chunk_width-1 downto 0);
	signal MT, ML, ST, DiagIn, SD, MR, MD, DiagOut: TwoDChunkArray(0 to NumChunks-1, 0 to NumChunks-1);



	signal rdy_array: std_logic_vector(0 to 2*NumChunks);

        -- the multiplier cells are arranged in a NumChunk X NumChunk array.
        -- Cell (I,J) receives R(I) (MT),  L(J) (MR) and a partial sum from above (ST).
	-- Cell (I,J) receives an incoming diagonal sum from Cell (I-1,J+1) and
        -- passes on its sum to the diagonal block Cell (I+1,J-1).
	--
	component DelayCell 
   		generic (operand_width: integer; delay: natural);
   		port (Din: in unsigned(operand_width-1 downto 0);
	 		Dout: out unsigned(operand_width-1 downto 0);
	 		clk: in std_logic;
	 		stall: in std_logic);
	end component DelayCell;

	component MultiplierCell is
  		generic (operand_width: integer);
  		port (MT, MR, ST, DiagIn: in unsigned(operand_width-1 downto 0);
        		ML, MD, SD, DiagOut: out unsigned(operand_width-1 downto 0);
        		stall: in std_logic;
			clk: in std_logic);
	end component MultiplierCell;

	component SumCell is
 		generic (operand_width: integer; ignore_diag: boolean; ignore_right: boolean);
		port (SU,SDiagIn: in unsigned(operand_width-1 downto 0);
              		SR: in unsigned(1 downto 0);
	      		SDiagOut: out unsigned(operand_width-1 downto 0);
	      		SL: out unsigned(1 downto 0);
	      		stall: in std_logic;
	      		clk: in std_logic);
	end component SumCell;

	type OneDChunkArray is array (natural range <>) of unsigned(chunk_width-1 downto 0);
	signal SU,SDiagIn,SDiagOut: OneDChunkArray(0 to NumChunks-1);

	type OneD2BitArray is array (natural range <>) of unsigned(1 downto 0);
        signal SR,SL: OneD2BitArray(0 to NumChunks-1);

	signal result_array : OneDChunkArray(0 to (2*NumChunks)-1);
begin

	process(L)
		variable lpad : unsigned(padded_operand_width-1 downto 0);
	begin
		lpad := (others => '0');
		lpad(operand_width-1 downto 0) := L;
		Lpadded <= lpad;
	end process;

	process(R)
		variable rpad : unsigned(padded_operand_width-1 downto 0);
	begin
		rpad := (others => '0');
		rpad(operand_width-1 downto 0) := R;
		Rpadded <= rpad;
	end process;

	RESULT <= RESULTpadded((2*operand_width)-1 downto 0);

	tag_array(0) <= tag_in;
	rdy_array(0) <= in_rdy;
	
	Tags: for ROW in 1 to (2*NumChunks) generate
		process(clk)
		begin
			if(clk'event and clk = '1') then
				if(reset = '1') then
					rdy_array(ROW) <= '0';
					tag_array(ROW) <= (others => '0');
				elsif(stall = '0') then
					tag_array(ROW) <= tag_array(ROW-1);
					rdy_array(ROW) <= rdy_array(ROW-1);
				end if;
			end if;
		end process;
	end generate Tags;
	tag_out <= tag_array(2*NumChunks);
	out_rdy <= rdy_array(2*NumChunks);

	Rows: for ROW in 0 to NumChunks-1 generate
		Cols: for COL in 0 to NumChunks-1 generate

			-- incoming  L values get into MT(0,-).
			ROWBC: if ROW = 0 generate
                                MT(ROW,COL) <= Lpadded(((COL+1)*chunk_width)-1 downto (COL*chunk_width));

				-- incoming signals to top row are 0.
				DiagIn(ROW,COL) <= (others => '0');
				ST(ROW,COL) <= (others => '0');

			end generate ROWBC;

		        COLBC: if COL=NumChunks-1 and ROW>0 generate
				-- left border column has incoming diagonals 0
				DiagIn(ROW,COL) <= (others => '0');
			end generate COLBC;

			-- from the right, R values enter with each row 
			-- getting an appropriate delay.
			COLBC2: if COL = 0 generate
				delInst: DelayCell generic map(operand_width => chunk_width,
								delay => ROW)
					port map(Din => Rpadded(((ROW+1)*chunk_width)-1 downto (ROW*chunk_width)),
						 Dout => MR(ROW,COL),
						 clk => clk,
						 stall => stall);
			end generate COLBC2;

			-- passing from right to left.
			Cols1: if COL > 0 generate
				MR(ROW,COL) <= ML(ROW,COL-1);
			end generate Cols1;

			ConnectArray: if ROW>0 generate

				-- from top to bottom
				MT(ROW,COL) <= MD(ROW-1,COL);
				ST(ROW,COL) <= SD(ROW-1,COL);
				
				-- diagonally.
				Cols2: if COL < NumChunks-1 generate
					DiagIn(ROW,COL) <= DiagOut(ROW-1,COL+1);
				end generate Cols2;
			end generate ConnectArray;

			mulCell: MultiplierCell generic map(operand_width => chunk_width)
				port map(MT => MT(ROW,COL),
					 ML => ML(ROW,COL),
					 ST => ST(ROW,COL),
					 DiagIn => DiagIn(ROW,COL),
					 SD => SD(ROW,COL),
					 MR => MR(ROW,COL),
					 MD => MD(ROW,COL),
					 stall => stall,
					 DiagOut => DiagOut(ROW,COL),
					 clk => clk);
		end generate Cols;
	end generate Rows;


	--  instantiate an array of sum cells to take
	--  care of the SD correction.
	sumArray: for Cols in 0 to NumChunks-1 generate
	
		scell: SumCell generic map (operand_width => chunk_width,
						ignore_diag => (Cols = NumChunks-1),
						ignore_right => (Cols = 0))
			port map(SU => SU(Cols),
				 SDiagIn => SDiagIn(Cols),
				 SR => SR(Cols),
				 SDiagOut => SDiagOut(Cols),
				 SL => SL(Cols),
				 stall => stall,
				 clk => clk);

		BR: if(Cols = 0) generate
			-- 0s from the right at the right boundary
			SR(Cols) <= (others => '0');
		end generate BR;
				
		BL: if(Cols = NumChunks-1) generate
			-- 0s from the diagonal at the left boundary.
			SDiagIn(Cols) <= (others => '0');
		end generate BL;

		--   inputs to the cells are delayed to match the sum
		--   propagation.

		--  sum coming down..
		dSU: DelayCell generic map(operand_width => chunk_width, delay => Cols)
			port map(Din => SD(NumChunks-1,Cols),
				 Dout => SU(Cols),
				 clk => clk,
				 stall => stall);
		
		Cntr1: if(Cols > 0) generate
			SR(Cols) <= SL(Cols-1);
		end generate Cntr1;
		
		Cntr2: if (Cols < NumChunks-1) generate
			-- diagonal coming in..  the leftmost cell has no incoming diagonal.
			dSDiagIn: DelayCell generic map(operand_width => chunk_width, delay => Cols)
				port map(Din => DiagOut(NumChunks-1,Cols+1),
				 Dout => SDiagIn(Cols),
				 clk => clk,
				 stall => stall);
		end generate Cntr2;
		
	end generate sumArray;


	--       instantiate delay elements to match delays
        --       inserted due to sum-cell array.


	-- the right column has 2*N-1 delays inserted.
	RightColumn:  for Rows in 0 to NumChunks-1 generate
		dRc: DelayCell generic map(operand_width => chunk_width, delay => ((2*NumChunks)-1) - Rows)
			port map(Din => DiagOut(Rows,0),
				 Dout => result_array(Rows),
				 stall => stall,
				 clk => clk);
	end generate RightColumn;

	-- the bottom row has N-C delays inserted as C goes from 0 to N-2
	BottomRow: for Cols in 0 to NumChunks-2 generate
		dBr: DelayCell generic map(operand_width => chunk_width, delay => NumChunks-(Cols+1))
			port map(Din => SDiagOut(Cols),
				 Dout => result_array(Cols+NumChunks),
				 stall => stall,
				 clk => clk);
		
	end generate BottomRow;

	-- leftmost element has no delays inserted.
	result_array((2*NumChunks)-1) <= SDiagOut(NumChunks-1);


	-- result: pack the diagonals into the result vector.
	process(result_array)
	begin
		for I in 0 to (2*NumChunks)-1 loop
			RESULTpadded(((I+1)*chunk_width)-1 downto (I*chunk_width))
				<= result_array(I);
		end loop;
	end process;

end ArrayMul;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- a basic unsigned shifter.
--
-- for the moment, this just does a shift and adds delay stages at
-- the end; presumably, the synthesis tool will retime things
-- appropriately..
--
-- TODO: pipeline this explicitly!
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Utilities.all;


entity UnsignedShifter is
  
  generic (
    name:string;
    shift_right_flag   : boolean;
    tag_width          : integer;
    operand_width      : integer;
    shift_amount_width : integer);

  port (
    L       : in  unsigned(operand_width-1 downto 0);
    R       : in  unsigned(shift_amount_width-1 downto 0);
    RESULT     : out unsigned(operand_width-1 downto 0);
    clk, reset : in  std_logic;
    in_rdy     : in  std_logic;
    out_rdy    : out std_logic;
    stall      : in std_logic;
    tag_in     : in std_logic_vector(tag_width-1 downto 0);
    tag_out    : out std_logic_vector(tag_width-1 downto 0));
end entity;


architecture Pipelined of UnsignedShifter is

  constant phases_per_stage: integer := 8;
  constant num_sig_bits: integer := Maximum(1,Minimum(shift_amount_width, Ceil_Log2(operand_width)));
  constant pipe_depth : integer := Ceil(num_sig_bits,phases_per_stage);

  type RWORD is array (natural range <>) of unsigned(operand_width-1 downto 0);
  type TWORD is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);  
  type SWORD is array (natural range <>) of unsigned(num_sig_bits-1 downto 0);  


  signal intermediate_results : RWORD(0 to pipe_depth);
  signal intermediate_tags : TWORD(0 to pipe_depth);  
  signal intermediate_shift_amount : SWORD(0 to pipe_depth);  
  signal stage_active : std_logic_vector(0 to pipe_depth);

  
  constant debug_flag: boolean := global_debug_flag;
begin  -- Pipelined

  Debug: if debug_flag  generate
	
	DebugBlock: block
		signal pipe_depth_sig, num_sig_bits_sig, tmp_sig, tmp_sig_2: integer;
	begin
		pipe_depth_sig <= pipe_depth;
		num_sig_bits_sig <= num_sig_bits;
		tmp_sig <= Ceil(num_sig_bits,phases_per_stage);
		tmp_sig_2 <= (num_sig_bits/phases_per_stage);
	end block;

  end generate debug;

   
  TrivOp: if operand_width = 1 generate
	intermediate_results(0) <= (others => '0') when R(0) = '1' else L;
  end generate TrivOp;
  

  NonTrivOp: if operand_width > 1 generate



        genStages: for STAGE in 1 to pipe_depth generate
  		process(clk, reset, stall, stage_active, intermediate_results, intermediate_shift_amount)
			variable shifted_L: unsigned(operand_width-1 downto 0);
			variable shift_amount: unsigned(num_sig_bits-1 downto 0);
  		begin
			shifted_L := intermediate_results(STAGE-1);
			shift_amount := intermediate_shift_amount(STAGE-1);

			for I in ((STAGE-1)*phases_per_stage) to 
					Minimum(num_sig_bits-1,(STAGE*phases_per_stage)-1) loop  
				if(shift_amount(I) = '1') then
					if(shift_right_flag) then
						shifted_L :=  shift_right(shifted_L, 2**I);
					else
						shifted_L :=  shift_left(shifted_L, 2**I);
					end if;
				end if;
			end loop;

			if(clk'event and clk='1') then

                                if(reset = '1') then
					stage_active(STAGE) <=  '0';
				elsif stall = '0' then
					stage_active(STAGE) <= stage_active(STAGE-1);
  					intermediate_results(STAGE) <= shifted_L;
  					intermediate_tags(STAGE) <= intermediate_tags(STAGE-1);
					intermediate_shift_amount(STAGE) <= 
							intermediate_shift_amount(STAGE-1);
				end if;
			end if;
  		end process;
	end generate genStages;

  end generate NonTrivOp;


  -- I/O
  intermediate_results(0) <=  L;
  intermediate_tags(0) <= tag_in;
  intermediate_shift_amount(0) <= R(num_sig_bits-1 downto 0);
  stage_active(0) <= in_rdy;
  out_rdy <= stage_active(pipe_depth);
  tag_out <= intermediate_tags(pipe_depth);
  RESULT <= intermediate_results(pipe_depth);
  
end Pipelined;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity CounterBase is 
	generic(name: string; data_width : integer);
	port(clk, reset: in std_logic; count_out: out std_logic_vector(data_width-1 downto 0));
end CounterBase;


architecture Behave of CounterBase is
	signal counter_sig: unsigned(data_width-1 downto 0);
begin
	process(clk)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				counter_sig <= (others => '0');
			else
				counter_sig <= counter_sig + 1;
			end if;
		end if;
	end process;

	count_out <= std_logic_vector(counter_sig);
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity InputMuxWithBuffering is
  generic (name: string;
	   iwidth: integer := 10;
	   owidth: integer := 10;
	   twidth: integer := 3;
	   nreqs: integer := 1;
	   buffering: IntegerArray;
	   no_arbitration: Boolean := false;
	   registered_output: Boolean := true;
	   full_rate: boolean);
  port (
    -- req/ack follow pulse protocol
    reqL                 : in  BooleanArray(nreqs-1 downto 0);
    ackL                 : out BooleanArray(nreqs-1 downto 0);
    dataL                : in  std_logic_vector(iwidth-1 downto 0);
    -- output side req/ack level protocol
    reqR                 : out std_logic;
    ackR                 : in  std_logic;
    dataR                : out std_logic_vector(owidth-1 downto 0);
    -- tag specifies the requester index 
    tagR                : out std_logic_vector(twidth-1 downto 0);
    clk, reset          : in std_logic);
end InputMuxWithBuffering;


architecture Behave of InputMuxWithBuffering is

  type WordArray is array (natural range <>) of std_logic_vector(owidth-1 downto 0);
  signal rx_data_in, rx_data_out : WordArray(nreqs-1 downto 0);

  signal reqFromRx, ackToRx: std_logic_vector(nreqs-1 downto 0);
  signal fairReqs, fairAcks: std_logic_vector(nreqs-1 downto 0);
  signal reqP, ackP: std_logic_vector(nreqs-1 downto 0);
  signal reqFair, ackFair: std_logic_vector(nreqs-1 downto 0);

  signal kill_zero: std_logic;
  signal reqR_sig, ackR_sig: std_logic;
  signal dataR_sig: std_logic_vector(owidth-1 downto 0);
  signal tagR_sig                : std_logic_vector(twidth-1 downto 0);
  signal oq_data_in : std_logic_vector((twidth + owidth)-1 downto 0);
  signal oq_data_out : std_logic_vector((twidth + owidth)-1 downto 0);

  --alias cbuffering: IntegerArray(nreqs-1 downto 0) is buffering;

begin  -- Behave

   kill_zero <= '0';


  assert(iwidth = owidth*nreqs) report "mismatched i/o widths in InputMuxBase" severity error;

  -----------------------------------------------------------------------------
  -- first stage: receive buffers.
  -----------------------------------------------------------------------------
  RxGen: for I in 0 to nreqs-1 generate 
     process(dataL)
        --variable regv : std_logic_vector(owidth-1 downto 0);
     begin
        -- Extract(dataL,I,regv);
        rx_data_in(I) <= dataL(((I+1)*owidth)-1 downto I*owidth);
     end process;


     rxBuf: ReceiveBuffer generic map(name => name & "-rxBuf-" & Convert_To_String(I),
					buffer_size =>  buffering(I),
					data_width => owidth,
					full_rate => full_rate)
		port map (write_req => reqL(I),
			  write_ack => ackL(I),
			  write_data => rx_data_in(I),
			  -------------------------
			  -- note: cross-over.
			  read_req => ackToRx(I),
			  read_ack => reqFromRx(I),
			  -------------------------
			  read_data => rx_data_out(I),
			  clk => clk, reset => reset);
					
  end generate RxGen;

  -----------------------------------------------------------------------------
  -- second-stage "fairify" the level-reqs (to avoid starvation).
  -----------------------------------------------------------------------------
  fairify: NobodyLeftBehind generic map (name => name & "-fairify", num_reqs => nreqs)
		port map (clk => clk, reset => reset, reqIn => reqFromRx, ackOut => ackToRx,
					reqOut => reqFair, ackIn => ackFair);


  -----------------------------------------------------------------------------
  -- priority encoding or pass through
  -----------------------------------------------------------------------------
  NoArbitration: if no_arbitration generate
    reqP <= reqFair;
    reqR_sig <= OrReduce(reqP);
    ackFair <= reqP when ackR_sig = '1' else (others => '0');
  end generate NoArbitration;

  Arbitration: if not no_arbitration generate
    reqP <= PriorityEncode(reqFair);
    reqR_sig <= OrReduce(reqP);
    ackFair <= reqP when ackR_sig = '1' else (others => '0');
  end generate Arbitration;

  -----------------------------------------------------------------------------
  -- data multiplexor
  -----------------------------------------------------------------------------
  process(reqP,rx_data_out)
  begin
    dataR_sig <= (others => '0');
    for J in 0 to nreqs-1 loop
      if(reqP(J) = '1') then
        dataR_sig <= rx_data_out(J);
        exit;
      end if;
    end loop;
  end process;    

  -----------------------------------------------------------------------------
  -- tag generation
  -----------------------------------------------------------------------------
  taggen : BinaryEncoder generic map (
    name => name & "-taggen",
    iwidth => nreqs,
    owidth => twidth)
    port map (
      din  => reqP,
      dout => tagR_sig);

  -----------------------------------------------------------------------------
  -- output queue.. data and tag passed out of mux. 
  -- TODO: link the output queue to the input muxing to save
  --       one stage?
  -----------------------------------------------------------------------------
  ifReg: if registered_output generate
        
      oqueue : QueueBase generic map (
	name => name & "-oqueue",
        queue_depth => 2,
        data_width  => twidth + owidth)
        port map (
          clk      => clk,
          reset    => reset,
          data_in  => oq_data_in,
          push_req => reqR_sig,
          push_ack => ackR_sig,
          data_out => oq_data_out,
          pop_ack  => reqR,
          pop_req  => ackR);
      
  end generate ifReg;

  ifNoReg: if (not registered_output) generate
     oq_data_out <= oq_data_in;
     reqR <= reqR_sig;
     ackR_sig <= ackR;
  end generate ifNoReg;

  oq_data_in <= dataR_sig & tagR_sig;
  dataR <= oq_data_out((twidth+owidth)-1 downto twidth);
  tagR  <= oq_data_out(twidth-1 downto 0);

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Components.all;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

--
-- a full-rate input port.  The assumption here
-- is that a data item is picked up from the
-- input port for every req pulse.  The production
-- of a new output data-item is indicated by an
-- ack pulse.
--
entity InputPortRevised is
  generic (name : string;
	   num_reqs: integer;
	   data_width: integer;
	   output_buffering: IntegerArray;
	   nonblocking_read_flag: boolean := false;
	   no_arbitration: boolean := false);
  port (
    -- pulse interface with the data-path
    sample_req        : in  BooleanArray(num_reqs-1 downto 0); -- sacrificial.
    sample_ack        : out BooleanArray(num_reqs-1 downto 0); -- sacrificial.
    update_req        : in  BooleanArray(num_reqs-1 downto 0);
    update_ack        : out BooleanArray(num_reqs-1 downto 0);
    data              : out std_logic_vector((num_reqs*data_width)-1 downto 0);
    -- ready/ready interface with outside world
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : in  std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
end entity;


architecture Base of InputPortRevised is

  --alias outBUFs: IntegerArray(num_reqs-1 downto 0) is output_buffering;
  signal has_room, write_enable : std_logic_vector(num_reqs-1 downto 0);

  type   IPWArray is array(integer range <>) of std_logic_vector(data_width-1 downto 0);
  signal write_data, read_data: IPWArray(num_reqs-1 downto 0);

  signal demux_data : std_logic_vector((num_reqs*data_width)-1 downto 0);

  signal ack_raw: BooleanArray(num_reqs-1 downto 0);
  
  type FsmState is (Idle, Waiting);
   
  -- to deal with nonblocking case..
  signal oreq_qualified       : std_logic;
  signal oack_qualified       : std_logic;
  signal odata_qualified      : std_logic_vector(data_width-1 downto 0);

  constant c_d_0      : std_logic_vector(data_width-1 downto 0) := (others => '0');

  -- bypass if there is only one requester.
  constant bypass_flag : boolean := (num_reqs = 1);

begin

  -----------------------------------------------------------------------------
  -- non-block/block qualification.. no need to do it here since nonblock
  -- functionality is present in UnloadRegister.
  -----------------------------------------------------------------------------
  oreq <= oreq_qualified;
  oack_qualified <= oack;
  odata_qualified <= odata;


  -----------------------------------------------------------------------------
  -- data register for every requester.
  -----------------------------------------------------------------------------
  ProTx : for I in 0 to num_reqs-1 generate

    --
    -- Note: for correct functioning of this input port
    --   external dependencies on the control-path side
    --   must be correctly setup.
    --     sr->sa->cr->ca chain
    --     ca -o-> sr  (0-delay) dependency.
    --
    sample_ack(I) <= sample_req(I); -- to maintain illusion of split protocol.

    -- the unload-register..
    ulreg: UnloadRegister
		generic map (name => name & "-unload-reg",
				data_width => data_width,
				bypass_flag => bypass_flag,
				nonblocking_read_flag => nonblocking_read_flag)	
		port map (write_req => write_enable(I),
				write_ack => has_room(I),
				  write_data => write_data(I),
				unload_req => update_req(I),
				  unload_ack => update_ack(I),
				   read_data => read_data(I),
				     clk => clk, reset => reset);
  end generate ProTx;

  demux : InputPortLevel generic map (
    name => name & "-demux",
    num_reqs       => num_reqs,
    data_width     => data_width,
    no_arbitration => no_arbitration)
    port map (
      req => has_room,
      ack => write_enable,
      data => demux_data,
      oreq => oreq_qualified,
      odata => odata_qualified,
      oack => oack_qualified,
      clk => clk,
      reset => reset);

  -----------------------------------------------------------------------------
  -- data handling
  -----------------------------------------------------------------------------
  process(read_data)
    variable ldata: std_logic_vector((num_reqs*data_width)-1 downto 0);
  begin
    for J in num_reqs-1 downto 0 loop
      ldata(((J+1)*data_width)-1 downto J*data_width) := read_data(J);
    end loop;
    data <= ldata;
  end process;

  gen : for I in num_reqs-1 downto 0 generate
    write_data(I) <= demux_data(((I+1)*data_width)-1 downto I*data_width); 
  end generate gen;

end Base;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity InterlockBuffer is
  generic (name: string; buffer_size: integer := 2; 
  	in_data_width : integer := 32;
  	out_data_width : integer := 32;
  	flow_through: boolean := false;
	cut_through : boolean := false;
  	bypass_flag : boolean := false);
  port (write_req: in boolean;
        write_ack: out boolean;
        write_data: in std_logic_vector(in_data_width-1 downto 0);
        read_req: in boolean;
        read_ack: out boolean;
        read_data: out std_logic_vector(out_data_width-1 downto 0);
        clk : in std_logic;
        reset: in std_logic);
end InterlockBuffer;

architecture default_arch of InterlockBuffer is

  constant data_width: integer := Minimum(in_data_width,out_data_width);

  signal buf_write_req, buf_write_ack: std_logic;
  signal buf_write_data, buf_read_data:  std_logic_vector(data_width-1 downto 0);

  type LoadFsmState is (l_idle, l_busy);
  signal l_fsm_state : LoadFsmState;

  signal has_data: std_logic;

  -- Don't F-around with this.
  constant use_unload_register : boolean := 
		((not global_use_optimized_unload_buffer) and (not cut_through))
		or (global_use_optimized_unload_buffer and (not cut_through) and (buffer_size /= 2));

  --
  -- Do not slow down the interlock buffer!
  --
  constant use_simple_ilock_implementation :boolean 
			:= global_use_optimized_unload_buffer and
					(not flow_through) and  (buffer_size = 1) and
						(not bypass_flag); 
			
  
-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- default_arch

  -- interlock buffer must have buffer-size > 0
  assert buffer_size > 0 report " interlock buffer size must be > 0 " severity failure;
  
  flowThrough: if flow_through generate

    write_ack <= write_req;
    read_ack <= read_req;

    inSmaller: if in_data_width <= out_data_width generate
      process(write_data)
        variable rvar : std_logic_vector(out_data_width-1 downto 0);
      begin
        rvar := (others => '0');
        rvar(in_data_width-1 downto 0) := write_data;
        read_data <= rvar;
      end process;
    end generate inSmaller;

    outSmaller: if out_data_width < in_data_width generate
      read_data <= write_data(out_data_width-1 downto 0);
    end generate outSmaller;

  end generate flowThrough;

  NoFlowThrough: if (not flow_through) generate


    interlockBuf: if (buffer_size > 0) generate
      inSmaller: if in_data_width <= out_data_width generate
        buf_write_data <= write_data;
  
        process(buf_read_data)
          begin
          read_data <= (others => '0');
          read_data(data_width-1 downto 0)  <= buf_read_data;
        end process;
      end generate inSmaller;
  
      outSmaller: if out_data_width < in_data_width generate
        buf_write_data <= write_data(data_width-1 downto 0);
        read_data  <= buf_read_data;
      end generate outSmaller;
      
      SimpleImplGen: if use_simple_ilock_implementation  generate
         sb: block
             signal joined_sig: boolean;
         begin

		cj: join2 generic map (bypass => true, name => "simpleImplGen:join2")
			port map (pred0 => write_req, pred1 => read_req, 
					symbol_out => joined_sig, 
						clk => clk, reset => reset);

		write_ack <= joined_sig;
		process(clk, reset, joined_sig, buf_write_data)
		begin
			if (clk'event and (clk = '1')) then 
				if(reset = '1') then
					read_ack <= false;
				else
					if(joined_sig) then
						buf_read_data <= buf_write_data;
					end if;
					read_ack <= joined_sig;
				end if;
			 end if;	
		end process;
         end block sb;
      end generate SimpleImplGen;

      ulbImplGen: if (not use_simple_ilock_implementation) generate
         -- write FSM to pipe.
         process(clk,reset, l_fsm_state, buf_write_ack, write_req)
           variable nstate : LoadFsmState;
         begin
           nstate := l_fsm_state;
           buf_write_req <= '0';
           write_ack <= false;
           if(l_fsm_state = l_idle) then
	     if(write_req) then
               buf_write_req <= '1';
               if(buf_write_ack = '1') then
                 write_ack <= true;
               else
                 nstate := l_busy;
               end if;
	     end if;
           else
	     buf_write_req <= '1';
	     if(buf_write_ack = '1') then
               nstate := l_idle;
               write_ack <= true;
	     end if;
           end if;
     
           if(clk'event and clk = '1') then
	     if(reset = '1') then
               l_fsm_state <= l_idle;
	     else
               l_fsm_state <= nstate;
	     end if;
           end if;
         end process;
     
         -- the unload buffer.
         buf : UnloadBuffer generic map (
           name =>  name & " buffer ",
           data_width => data_width,
           buffer_size => buffer_size, 
	   use_unload_register => use_unload_register,
           bypass_flag => bypass_flag)
           port map (
             write_req   => buf_write_req,
             write_ack   => buf_write_ack,
             write_data  => buf_write_data,
             unload_req  => read_req,
             unload_ack  => read_ack,
             read_data   => buf_read_data,
 	     has_data => has_data,
             clk         => clk,
             reset       => reset);
  
	end generate ulbImplGen; 
       end generate interlockBuf;
     end generate NoFlowThrough;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;


-- a simple multiplexor with output
-- queue.
entity LevelMux is
  generic(name:string;
	  num_reqs: integer;
	  data_width: integer;
	  no_arbitration: boolean := true);
  port (
    write_req       : in  std_logic_vector(num_reqs-1 downto 0);
    write_ack       : out std_logic_vector(num_reqs-1 downto 0);
    write_data      : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
    read_req        : in  std_logic;
    read_ack        : out std_logic;
    read_data       : out std_logic_vector(data_width-1 downto 0);
    clk, reset      : in  std_logic);
end entity;

architecture Base of LevelMux is
  
  type OPWArray is array(integer range <>) of std_logic_vector(data_width-1 downto 0);
  signal data_array : OPWArray(num_reqs-1 downto 0);
  signal req_active, ack_sig , fair_reqs, fair_acks : std_logic_vector(num_reqs-1 downto 0);
  
  signal q_data_in,q_data_out  : std_logic_vector(data_width-1 downto 0);
  signal q_push_req, q_push_ack, q_pop_req, q_pop_ack: std_logic;
begin

  -- input arbitration.
  fairify: NobodyLeftBehind generic map(name => name & "-fairify", num_reqs => num_reqs)
		port map(clk => clk, reset => reset,
				reqIn => write_req,
				ackOut => write_ack,
				reqOut => fair_reqs,
				ackIn => fair_acks);
  
  NoArb: if no_arbitration generate
     req_active <= fair_reqs;
  end generate NoArb;

  Arb: if not no_arbitration generate
     req_active <= PriorityEncode(fair_reqs);
  end generate Arb;


  -- combinational multiplexor (AND-OR form).
  -- AND
  gen: for I in num_reqs-1 downto 0 generate

       ack_sig(I) <= req_active(I) and q_push_ack; 
       fair_acks(I) <= ack_sig(I);

       process(write_data,req_active(I))
         variable target: std_logic_vector(data_width-1 downto 0);
       begin
          if(req_active(I) = '1') then
		-- Extract(write_data,I,target);
		target := write_data(((I+1)*data_width)-1 downto I*data_width);
	  else
		target := (others => '0');
	  end if;	
       	  data_array(I) <= target;
       end process;
  end generate gen;

  -- OR
  process (data_array)
    variable var_odata : std_logic_vector(data_width-1 downto 0) := (others => '0');
  begin  -- process
    var_odata := (others => '0');
    for I in 0 to num_reqs-1 loop
      var_odata := data_array(I) or var_odata;
    end loop;  -- I
    q_data_in <= var_odata;
  end process;


  -- output queue (2 stage).
  q_push_req <= OrReduce(req_active);
  q_pop_req  <= read_req;
  read_ack   <= q_pop_ack;
  read_data  <= q_data_out;
  oQ:  QueueBase generic map(name => "-oQ", queue_depth => 2, data_width => data_width)
	port map( clk => clk, reset => reset,
			data_in => q_data_in,
			push_req => q_push_req,
			push_ack => q_push_ack,
			data_out => q_data_out,
			pop_req => q_pop_req,
			pop_ack => q_pop_ack);
end Base;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;

--
-- at the input side, introduce a receive
-- buffer into which the input data is concatenated
-- with a tag and a time-stamp.
--
-- The receive buffers are muxed using a merge
-- tree that compares the time-stamps.
-- From the output of the merge-tree, the data
-- and tag are separated to produce maddr, mtag.
--
entity LoadReqSharedWithInputBuffers is
  generic
    (
	name : string;
	addr_width: integer := 8;
      	num_reqs : integer := 1; -- how many requesters?
	tag_length: integer := 1;
	no_arbitration: Boolean := false;
        min_clock_period: Boolean := true;
	input_buffering: IntegerArray;
	time_stamp_width: integer := 0
    );
  port (
    -- req/ack follow pulse protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    -- concatenated address corresponding to access
    dataL                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
    -- address to memory
    maddr                   : out std_logic_vector((addr_width)-1 downto 0);
    mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);

    mreq                    : out std_logic;
    mack                    : in std_logic;
    -- clock, reset (active high)
    clk, reset              : in std_logic);
end LoadReqSharedWithInputBuffers;

architecture Vanilla of LoadReqSharedWithInputBuffers is

  constant iwidth: integer := addr_width*num_reqs;
  constant owidth: integer := addr_width;

  constant debug_flag : boolean := global_debug_flag;

  -- must register..  ack implies that address has been sampled.
  constant registered_output : boolean := true; 

  type TagWordArray is array (natural range <>) of unsigned(tag_length-1 downto 0);
  signal rx_tag_in: TagWordArray(num_reqs-1 downto 0);

  constant rx_word_length: integer := addr_width + tag_length + time_stamp_width;
  type RxBufWordArray is array (natural range <>) of std_logic_vector(addr_width + tag_length + time_stamp_width-1 downto 0);

  signal rx_data_in, rx_data_out : RxBufWordArray(num_reqs-1 downto 0);
  signal kill_sig : std_logic;

  signal imux_data_in_accept,  imux_data_in_valid: std_logic_vector(num_reqs-1 downto 0);
  signal imux_data_in: std_logic_vector((rx_word_length*num_reqs)-1 downto 0);

  signal imux_data_out_accept,  imux_data_out_valid: std_logic;
  signal imux_data_out: std_logic_vector(rx_word_length-1 downto 0);
  
  --alias IBUFs: IntegerArray(num_reqs-1 downto 0) is input_buffering;
begin  -- Behave

  assert(tag_length >= Ceil_Log2(num_reqs)) report "insufficient tag width" severity error;
 
  kill_sig <= '0'; -- no killing!

  tagGen: for I in 0 to num_reqs-1 generate
	rx_tag_in(I) <= To_Unsigned(I,tag_length);	
  end generate tagGen;


  TstampGen: if time_stamp_width > 0 generate
	Tsb: block 
		signal time_stamp: std_logic_vector(time_stamp_width-1 downto 0);
	begin
		tsc: CounterBase generic map(name => name & "-TstampGen-Tsb", data_width => time_stamp_width)
			port map(clk => clk, reset => reset, count_out => time_stamp);

		rxInDataGen: for I in 0 to num_reqs-1 generate
			rx_data_in(I) <= dataL(((I+1)*addr_width)-1 downto I*addr_width) & std_logic_vector(rx_tag_in(I)) & time_stamp;
		end generate rxInDataGen;
	end block Tsb;
  end generate TstampGen;

  NoTstampGen: if time_stamp_width < 1 generate
	rxInDataGen: for I in 0 to num_reqs-1 generate
		rx_data_in(I) <= dataL(((I+1)*addr_width)-1 downto I*addr_width) & std_logic_vector(rx_tag_in(I));
	end generate rxInDataGen;
  end generate NoTstampGen;

  -- receive buffers.
  RxGen: for I in 0 to num_reqs-1 generate
	rb: ReceiveBuffer generic map(name => name & "-RxGen-rb-" & Convert_To_String(I),
					buffer_size => Maximum(2,input_buffering(I)),
					data_width => rx_word_length,
					full_rate => false) -- Load-data-path will be double buffered.
		port map(write_req => reqL(I), 
			 write_ack => ackL(I), 
			 write_data => rx_data_in(I), 
			 read_req => imux_data_in_accept(I), 
			 read_ack => imux_data_in_valid(I), 
                         read_data => rx_data_out(I),
			 clk => clk, 
			 reset => reset);

  end generate RxGen;

  -- 2D to 1D array conversion.
  process(rx_data_out)
  begin
	for I in 0 to num_reqs-1 loop
		imux_data_in(((I+1)*rx_word_length)-1 downto (I*rx_word_length))
			<= rx_data_out(I);
        end loop;
  end process;

  -- the multiplexor.
  NonTrivTstamp: if time_stamp_width > 0 generate
  	imux: merge_tree
    	   generic map(name => name & "-NonTrivTstamp-imux",
		g_number_of_inputs => num_reqs,
		g_data_width => rx_word_length,
                g_time_stamp_width => time_stamp_width, 
                g_tag_width => tag_length,
		g_mux_degree => 4096, -- some large number.. allow big muxes.
		g_num_stages => 1,    -- with single stage delay 
		g_port_id_width => 0)
           port map(merge_data_in => imux_data_in,
	            merge_req_in  => imux_data_in_valid,
	            merge_ack_out => imux_data_in_accept,
	            merge_data_out => imux_data_out,
                    merge_req_out => imux_data_out_valid,
	            merge_ack_in  => imux_data_out_accept,
      	            clock        => clk,
      	            reset      => reset);
  end generate NonTrivTstamp;

  TrivTstamp: if time_stamp_width < 1 generate
	imux: LevelMux generic map (name => name & "-TrivTstamp-imux",
				num_reqs => num_reqs, data_width => rx_word_length, no_arbitration => false)
		port map(write_req => imux_data_in_valid,
			 write_ack => imux_data_in_accept,
			 write_data => imux_data_in,
			 read_req => imux_data_out_accept,
		         read_ack => imux_data_out_valid,
			 read_data => imux_data_out,
			 clk => clk, reset => reset);
  end generate TrivTstamp;


  -- outgoing tag, address.
  mreq <= imux_data_out_valid;
  imux_data_out_accept <= mack;
  maddr <= imux_data_out(rx_word_length-1 downto (tag_length + time_stamp_width));
  mtag <= imux_data_out(tag_length+time_stamp_width-1 downto 0);
  

end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- uses an aggressive pulse-to-level translation
-- that allows back-to-back transfers to an output
-- port.  The combinational paths are a bit longer
-- but cant have everything..
--
-- added full_rate flag to indicate that throughput is paramount.
entity OutputPortRevised is
  generic(name : string;
	  num_reqs: integer;
	  data_width: integer;
	  no_arbitration: boolean := false;
	  input_buffering: IntegerArray;
	  full_rate: boolean);
  port (
    sample_req        : in  BooleanArray(num_reqs-1 downto 0);
    sample_ack        : out BooleanArray(num_reqs-1 downto 0);
    update_req        : in  BooleanArray(num_reqs-1 downto 0); -- sacrificial.
    update_ack        : out BooleanArray(num_reqs-1 downto 0); -- sacrificial.
    data       : in  std_logic_vector((num_reqs*data_width)-1 downto 0);
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : out std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
end entity;

architecture Base of OutputPortRevised is

  signal reqR, ackR : std_logic_vector(num_reqs-1 downto 0);

  signal omux_data_in       : std_logic_vector((num_reqs*data_width)-1 downto 0);

  type   OPWArray is array(integer range <>) of std_logic_vector(data_width-1 downto 0);
  signal in_data_array, out_data_array : OPWArray(num_reqs-1 downto 0);
  
  constant input_buf_sizes: IntegerArray(num_reqs-1 downto 0) :=  input_buffering;

  signal zero_sig: std_logic;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

  zero_sig <= '0';

  -----------------------------------------------------------------------------
  -- protocol conversion
  -----------------------------------------------------------------------------
  BufGen : for I in 0 to num_reqs-1 generate
	
	in_data_array(I) <= data(((I+1)*data_width)-1 downto (I*data_width));
	
	--  
	-- update ack..
        --   Note: to prevent runaway,  the following dependencies must be
	--    imposed in the control path.
        --  
        --   sa -> cr
        --   ca -o-> sr (0-delay)
        --
	process(clk,reset)
        begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				update_ack(I) <= false;
			else
				update_ack(I) <= update_req(I); -- sacrificial.. to maintain pretense of split protocol.
			end if;
		end if;
	end process;

	rxB: ReceiveBuffer 
		generic map( name => name & "-rxB" & Convert_To_String(I),
				buffer_size => input_buf_sizes(I),
				data_width => data_width,
				full_rate => full_rate)
		port map(write_req => sample_req(I),
		 	write_ack => sample_ack(I),
		 	write_data => in_data_array(I),
		 	-- note: cross-over
		 	read_req =>  ackR(I),
		 	read_ack => reqR(I), 
	         	read_data => out_data_array(I),	
		 	clk => clk, reset => reset);

  end generate BufGen;

  process(out_data_array)
  begin
	for J in  0 to num_reqs-1 loop
		omux_data_in(((J+1)*data_width)-1 downto J*data_width) <= out_data_array(J);
	end loop;
  end process;


  mux : OutputPortLevel generic map (
    name => name & "-mux",
    num_reqs       => num_reqs,
    data_width     => data_width,
    no_arbitration => no_arbitration)
    port map (
      req   => reqR,
      ack   => ackR,
      data  => omux_data_in,
      oreq  => oreq,
      oack  => oack,
      odata => odata,
      clk   => clk,
      reset => reset);
end Base;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

--
-- a safe register with no combinational paths
-- from input to output or vice-versa.
--
entity PipelineRegister is
  generic (name : string; data_width: integer);
  port (
    read_req       : in  std_logic;
    read_ack       : out std_logic;
    read_data      : out std_logic_vector(data_width-1 downto 0);
    write_req       : in  std_logic;
    write_ack       : out std_logic;
    write_data      : in std_logic_vector((data_width-1) downto 0);
    clk, reset : in  std_logic);
  
end PipelineRegister;

architecture default_arch of PipelineRegister is

   type FsmState is (Empty, Full);
   signal fsm_state : FsmState;
   signal data_reg : std_logic_vector(data_width-1 downto 0);
  
begin  -- default_arch

	process(clk, reset, write_req, read_req, write_data, fsm_state)
		variable next_state : FsmState;
		variable read_ack_v, write_ack_v, latch_v : std_logic;
	begin
		next_state := fsm_state;
		read_ack_v := '0';
		write_ack_v := '0';
		latch_v := '0';
	
		case fsm_state is 
			when Empty =>
				write_ack_v := '1';
				if(write_req = '1') then
					next_state := Full;
					latch_v := '1';
				end if;
			when Full =>
				read_ack_v := '1';
				if(read_req = '1') then
					next_state := Empty;
				end if;
		end case;
					
		write_ack <= write_ack_v;
		read_ack  <= read_ack_v;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= Empty;
			else
				fsm_state <= next_state;
			end if;

			if(latch_v = '1') then
				data_reg <= write_data;
			end if;
		end if;
	end process;

	read_data <=  data_reg;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
--   re-engineered Queue core implementation to improve LUT count and critical path!
--   Why didn't I think of this before?
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity QueueBaseCore is
  generic(name : string := "Anon"; 
		queue_depth: integer := 3; 
		reverse_bypass_flag: boolean := false;
		data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       empty, full: out std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity QueueBaseCore;

architecture behave of QueueBaseCore is

  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin  -- SimModel

 pDZero:  if(queue_depth = 0) generate

	empty <= '1';
	full  <= '1';

	data_out <= data_in;

	push_ack <= pop_req;
	pop_ack  <= push_req;

 end generate pDZero;

 pDEq1: if (queue_depth = 1) generate
    bbb1: block
	signal qsize: std_logic;
	signal push_ack_sig, pop_ack_sig: std_logic;
    begin
   

     	rbpGen1: if (reverse_bypass_flag) generate
		push_ack_sig <= '1' when (qsize = '0') or (pop_req = '1') else '0';
     	end generate rbpGen1;

     	noRbpGen1: if (not reverse_bypass_flag) generate
		push_ack_sig <= '1' when (qsize = '0') else '0';
     	end generate noRbpGen1;
		
	pop_ack_sig  <= '1' when (qsize = '1') else '0';

	full  <= not push_ack_sig;
	empty <= not pop_ack_sig;

	push_ack <= push_ack_sig;
	pop_ack <= pop_ack_sig;
     	ob: block
        	signal queue_data: std_logic_vector(data_width-1 downto 0);
     	begin
		
		process(clk, reset, data_in, push_req, push_ack_sig, pop_req, pop_ack_sig, qsize, queue_data)
        		variable next_queue_data: std_logic_vector(data_width-1 downto 0);
			variable next_qsize: std_logic;
			variable push, pop: boolean;
		begin 
		 	next_qsize := qsize;
			next_queue_data := queue_data;

			push := (push_req = '1') and (push_ack_sig = '1');
			pop := (pop_req = '1') and (pop_ack_sig = '1');

			if (push and (not pop)) then
				next_qsize := '1';
			elsif (pop and (not push)) then
				next_qsize := '0';
			end if;

			if(push) then
				next_queue_data := data_in;
			end if;

			if(clk'event and (clk = '1')) then
				if(reset = '1') then
					qsize <= '0';
					queue_data <= (others => '0');
				else
					qsize <= next_qsize;
					queue_data <= next_queue_data;
				end if;
			end if;
		end process;

		data_out <= queue_data;
     	end block ob;
    end block bbb1;
 end generate pDEq1;
 
 pDGOne: if (queue_depth > 1) generate

     lb: block
     	signal queue_data: QueueArray (0 to queue_depth-1); 
        signal state_vector: std_logic_vector(queue_depth-1 downto 0);
        signal reverse_bypass_applicable : boolean;
	signal push_ack_sig, pop_ack_sig: std_logic;
	constant Zstatus: std_logic_vector(queue_depth-1 downto 0) := (others => '1');
     begin


	empty <= (not pop_ack_sig);
	full  <= (not push_ack_sig);
	
     	rbpGen: if (reverse_bypass_flag) generate

     		push_ack_sig <= '1' when ((state_vector(queue_depth-1) = '0') or reverse_bypass_applicable) else '0';
		reverse_bypass_applicable <= (state_vector = Zstatus) and (pop_req = '1');
     	end generate rbpGen;
	
     	noRbpGen: if (not reverse_bypass_flag) generate
     		push_ack_sig <= '1' when (state_vector(queue_depth-1) = '0')  else '0';
		reverse_bypass_applicable <= false;
     	end generate noRbpGen;
	push_ack <= push_ack_sig;

     	pop_ack_sig <= '1' when state_vector(0) = '1' else '0';
	pop_ack <= pop_ack_sig;

     	data_out <= queue_data(0);

	-- sequence of stages
	--   Each stage has the following inputs
	--        push pop  status(k+1) status(k) status(k-1)
	--   and performs actions as follows:
	--  -------------------------------------------------------------------
	--   status(k+1) status(k) status(k-1)   Action
	--  -------------------------------------------------------------------
	--      0           0            0        No action.
	--      0           0            1        If push.(~pop), then load din 
	--                                        into stage, set status(k) = 1
	--                                        Else, nothing.
	--      0           1            1        If push.pop then load din into
	--                                        stage, status stays the same.
	--                                        If (~push).pop set status(k) = 0
	--                                        Else nothing.
	--      1           1             1       If pop load data(k+1) into
	--                                        stage, keep status(k) = 1
	--                                        Else nothing.
	--  -------------------------------------------------------------------
	stageGen: for K in queue_depth-1 downto 0 generate 
		sb: block
		   -- signals
		   signal data_kp1: std_logic_vector(data_width-1 downto 0);
                   signal status_kp1, status_k, status_km1: std_logic;
		   signal stat_3 : std_logic_vector(2 downto 0); 
		   signal push, pop: boolean;
		begin
			push <= (push_req = '1') and (push_ack_sig = '1');
			pop  <= (pop_req = '1')  and (pop_ack_sig  = '1');

			stat_3 (1) <= state_vector(K);

			topGen: if (K = (queue_depth - 1)) generate
			    cb: block
                            begin
				stat_3 (2) <= '0';
				stat_3 (0) <= state_vector(K-1);
				data_kp1 <= (others => '0');
                            end block cb;
			end generate topGen;

			midGen: if (K < (queue_depth-1)) and (K > 0) generate 
			    cb: block
                            begin
				stat_3 (2) <= state_vector(K+1);
				stat_3 (0) <= state_vector(K-1);
				data_kp1 <= queue_data(K+1);
                            end block cb;
			end generate midGen;

			botGen: if (K = 0) generate
			    cb: block
                            begin
				stat_3 (2) <= state_vector(K+1);
				stat_3 (0) <= '1';
				data_kp1 <= queue_data(K+1);
                            end block cb;
			end generate botGen;
		
			status_k <= state_vector(K);

			process(clk, reset)
                   		variable next_status_k_var: std_logic;
				variable next_stage_data_var: std_logic_vector(data_width-1 downto 0);
			begin
				next_status_k_var := status_k;
				next_stage_data_var := queue_data(K);
				
				case stat_3 is
					when "001" =>
						if(push and (not pop)) then
							next_stage_data_var := data_in;
							next_status_k_var   := '1';
						end if;
					when "011" =>
						if (push and pop) then
							next_stage_data_var := data_in;
							next_status_k_var := '1';
						elsif ((not push) and pop) then
							next_status_k_var := '0';
						end if;
					when "111" =>
						if pop then
							next_stage_data_var := data_kp1;
						end if;
					when others => null;
				end case;	
			
				if(clk'event and (clk = '1')) then
					if(reset = '1') then
						state_vector(K) <= '0';
						queue_data(K) <= (others => '0');
					else
						state_vector(K) <= next_status_k_var;
						queue_data(K) <= next_stage_data_var;
					end if;
				end if;
			end process;
		end block sb;
	end generate stageGen;
     end block lb;
 end generate pDGOne;


end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


-- Save a slot, introduce a pop_req -> push_ack path.
entity QueueBaseSaveSlot is
  generic(name : string; queue_depth: integer := 2; data_width: integer := 32;
		save_one_slot: boolean := false);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity QueueBaseSaveSlot;

architecture behave of QueueBaseSaveSlot is



  constant physical_queue_depth: integer := queue_depth-1;
  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);
  function Incr(x: integer; M: integer) return integer is
  begin
    if(x < M) then
      return(x + 1);
    else
      return(0);
    end if;
  end Incr;


begin  -- SimModel

  assert (queue_depth > 0) report "QueueBaseSaveSlot " & name & " must have at least one slot"
			severity error;

 --
 -- 0-depth queue is just a set of wires.
 --
 triv: if physical_queue_depth = 0 generate
	push_ack <= pop_req;
	pop_ack  <= push_req;
	data_out <= data_in;
 end generate triv;



 qDGt0: if physical_queue_depth > 0 generate 
  NTB: block 
  	signal queue_array : QueueArray(physical_queue_depth-1 downto 0);
  	signal read_pointer, write_pointer : integer range 0 to physical_queue_depth-1;
  	signal incr_write_pointer, incr_read_pointer : integer range 0 to physical_queue_depth-1;
  	signal queue_size : integer range 0 to physical_queue_depth;
  begin
 
    assert (queue_size < physical_queue_depth) report "Queue " & name & " is full." severity note;
    assert (queue_size < (3*physical_queue_depth/4)) report "Queue " & name & " is three-quarters-full." severity note;
    assert (queue_size < (physical_queue_depth/2)) report "Queue " & name & " is half-full." severity note;
    assert (queue_size < (physical_queue_depth/4)) report "Queue " & name & " is quarter-full." severity note;

    qD1: if (physical_queue_depth = 1) generate
     incr_read_pointer <= read_pointer;
     incr_write_pointer <= write_pointer;
    end generate qD1;

    qDG1: if (physical_queue_depth > 1) generate
     incr_read_pointer <= Incr(read_pointer, physical_queue_depth-1);
     incr_write_pointer <= Incr(write_pointer, physical_queue_depth-1);
    end generate qDG1;

    push_ack <= '1' when (queue_size < physical_queue_depth) or (pop_req = '1') else '0';
    pop_ack  <= '1' when (queue_size > 0) else '0';

    -- bottom pointer gives the data in FIFO mode..
    data_out <= queue_array(read_pointer);
  
    -- single process
    process(clk, reset, read_pointer, write_pointer, incr_read_pointer, incr_write_pointer, queue_size, push_req, pop_req)
      variable qsize : integer range 0 to physical_queue_depth;
      variable push,pop : boolean;
      variable next_read_ptr,next_write_ptr : integer range 0 to physical_queue_depth-1;
    begin

      qsize := queue_size;
      push  := false;
      pop   := false;
      next_read_ptr := read_pointer;
      next_write_ptr := write_pointer;
      
      if (((pop_req = '1') or (qsize < physical_queue_depth)) and push_req = '1') then
          push := true;
      end if;
  
      if((qsize > 0) and pop_req = '1') then
          pop := true;
      end if;
  
  
      if(push) then
          next_write_ptr := incr_write_pointer;
      end if;
  
      if(pop) then
          next_read_ptr := incr_read_pointer;
      end if;
  
  
      if(pop and (not push)) then
          qsize := qsize - 1;
      elsif(push and (not pop)) then
          qsize := qsize + 1;
      end if;
        
  
      if(clk'event and clk = '1') then
        
	if(reset = '1') then
           queue_size <= 0;
           read_pointer <= 0;
           write_pointer <= 0;
           queue_array(0) <= (others => '0'); -- initially 0.
	else
           if(push) then
          	queue_array(write_pointer) <= data_in;
           end if;
        
           queue_size <= qsize;
           read_pointer <= next_read_ptr;
           write_pointer <= next_write_ptr;

        end if;
      end if;

    end process;
   end block NTB;
  end generate qDGt0;
  

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity QueueBaseWithBypass is
  generic(name : string; queue_depth: integer := 1; data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity QueueBaseWithBypass;

architecture behave of QueueBaseWithBypass  is

  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);
  function Incr(x: integer; M: integer) return integer is
  begin
    if(x < M) then
      return(x + 1);
    else
      return(0);
    end if;
  end Incr;

begin  -- SimModel

 --
 -- 0-depth queue is just a set of wires.
 --
 triv: if queue_depth = 0 generate
	push_ack <= pop_req;
	pop_ack  <= push_req;
	data_out <= data_in;
 end generate triv;


 nontriv: if queue_depth > 0 generate 
  NTB: block 
  	signal queue_array : QueueArray(queue_depth-1 downto 0);
  	signal read_pointer, write_pointer : integer range 0 to queue_depth-1;
  	signal queue_size : integer range 0 to queue_depth;
        signal data_out_from_queue : std_logic_vector(data_width-1 downto 0);
        signal bypass_signal: Boolean;
  begin
 
    assert (queue_size < queue_depth) report "Queue " & name & " is full." severity note;

    push_ack <= '1' when (bypass_signal or (queue_size < queue_depth)) else '0';
    pop_ack  <= '1' when (bypass_signal or (queue_size > 0)) else '0';

    -- bottom pointer gives the data in FIFO mode..
    data_out_from_queue <= queue_array(read_pointer);

    --
    -- if queue size = 0, and if push-req is true, then data is
    -- presented to data-out through the bypass path.
    --
    data_out <= data_in when bypass_signal else data_out_from_queue;

  
    -- single process
    process(clk, queue_size, push_req, pop_req, write_pointer, read_pointer)
      variable qsize : integer range 0 to queue_depth;
      variable push,pop : boolean;
      variable next_read_ptr,next_write_ptr : integer range 0 to queue_depth-1;
      variable bypass: boolean;
    begin

      qsize := queue_size;
      push  := false;
      pop   := false;
      next_read_ptr := read_pointer;
      next_write_ptr := write_pointer;

      bypass := ((qsize = 0) and  (push_req = '1') and (pop_req = '1'));
      bypass_signal <= bypass;
      
      if((qsize < queue_depth) and (push_req = '1') and (not bypass)) then
          push := true;
      end if;
  
      if((qsize > 0) and (pop_req = '1') and (not bypass)) then
          pop := true;
      end if;
  
  
      if(push) then
          next_write_ptr := Incr(next_write_ptr,queue_depth-1);
      end if;
  
      if(pop) then
         next_read_ptr := Incr(next_read_ptr,queue_depth-1);
      end if;
  
      if(pop and (not push)) then
         qsize := qsize - 1;
      elsif(push and (not pop)) then
         qsize := qsize + 1;
      end if;
        
  
      if(clk'event and clk = '1') then
        if(reset = '1') then
		queue_size <= 0;
		read_pointer <= 0;
		write_pointer <= 0;
	else
        	if(push) then
          		queue_array(write_pointer) <= data_in;
        	end if;
        	
        	queue_size <= qsize;
        	read_pointer <= next_read_ptr;
        	write_pointer <= next_write_ptr;
	end if;
      end if;
      
    end process;
   end block NTB;
  end generate nontriv;
  

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- TODO: add bypass path to the receive buffer.
--       this will reduce buffering requirements
--       by a factor of two (for full pipelining).
--
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity ReceiveBuffer  is
  generic (name: string; buffer_size: integer ; data_width : integer ; full_rate: boolean);
  port ( write_req: in boolean;
         write_ack: out boolean;
         write_data: in std_logic_vector(data_width-1 downto 0);
         read_req: in std_logic;
         read_ack: out std_logic;
         read_data: out std_logic_vector(data_width-1 downto 0);
         clk : in std_logic;
         reset: in std_logic);
end ReceiveBuffer;

architecture default_arch of ReceiveBuffer is

  signal push_req, push_ack, pop_req, pop_ack: std_logic_vector(0 downto 0);
  signal pipe_data_in:  std_logic_vector(data_width-1 downto 0);

  constant use_full_rate_repeater : boolean := (full_rate and (buffer_size = 1));

  type RxBufFsmState is (idle, busy);
  signal fsm_state : RxBufFsmState;

-- see comment above..
--##decl_synopsys_sync_set_reset##



begin  -- default_arch

  -- the output pipe.
  notFRR: if not use_full_rate_repeater generate
    bufPipe : PipeBase 
    generic map (
      name =>  name & "-bufPipe",
      num_reads  => 1,
      num_writes => 1,
      data_width => data_width,
      lifo_mode  => false,
      shift_register_mode => false,
      depth      => buffer_size,
      full_rate  => full_rate)
    port map (
        read_req   => pop_req,
        read_ack   => pop_ack,
        read_data  => read_data,
        write_req  => push_req,
        write_ack  => push_ack,
        write_data => write_data,
        clk        => clk,
        reset      => reset);
  end generate notFRR;

  FRR: if use_full_rate_repeater generate
    bufRptr: FullRateRepeater
    generic map (
      name =>  name & "-frrptr",
      data_width => data_width)
    port map ( clk => clk,reset => reset,
		data_in => write_data,
		data_out => read_data,
		push_req => push_req(0),
		pop_req => pop_req(0),
		push_ack => push_ack(0),
		pop_ack => pop_ack(0));
  end generate FRR;

  read_ack <= pop_ack(0);
  pop_req(0) <= read_req;

  -- FSM
  process(clk,reset, fsm_state, write_req, push_ack)
	variable nstate : RxBufFsmState;
	variable pushreqv: std_logic;
	variable decr: boolean;
	variable wackv : boolean;
  begin
	wackv := false;
	pushreqv := '0'; 

	nstate := fsm_state;
	case fsm_state is
		when idle => 
			if(write_req) then
				pushreqv := '1';
				if(push_ack(0) = '1') then 
					wackv := true;
				else
					nstate := busy;	
				end if;
			end if;
		when busy => 
			pushreqv := '1';
			if (push_ack(0) = '1') then
				nstate := idle;
				wackv := true;
			end if;
	end case;

	push_req(0) <= pushreqv;
	write_ack <= wackv;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			fsm_state <= idle;
		else
			fsm_state <= nstate;
		end if;
	end if;
		
  end process;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;

entity SelectSplitProtocol is
  generic(name: string; 
	  data_width: integer; 
	  buffering: integer; 
	  flow_through: boolean := false; 
	  full_rate: boolean );
  port(x,y: in std_logic_vector(data_width-1 downto 0);
       sel: in std_logic_vector(0 downto 0);
       z : out std_logic_vector(data_width-1 downto 0);
       sample_req: in boolean;
       sample_ack: out boolean;
       update_req: in boolean;
       update_ack: out boolean;
       clk,reset: in std_logic);
end SelectSplitProtocol;


architecture arch of SelectSplitProtocol is 
   signal ilb_data_in: std_logic_vector(data_width-1 downto 0);
begin

    
     -- if mux select is X during normal operations then we
     -- have a problem.
     -- assert (not (sample_req and clk'event  and (clk = '1') and (reset = '0')) 
		-- or (not is_x(sel(0)))) report "mux " & name & " select is X" severity error;

     ilb_data_in <=  x when (sel(0) = '1') else y;

     noFlowThrough: if (not flow_through) generate
    	ilb: InterlockBuffer 
		generic map(name => name & "-ilb",
				buffer_size => buffering,
				in_data_width => data_width,
				out_data_width => data_width)
		port map(write_req => sample_req,
			 write_ack => sample_ack,
			 write_data => ilb_data_in,
			 read_req  => update_req,
			 read_ack => update_ack,
			 read_data => z,
			 clk => clk, reset => reset);
     end generate noFlowThrough;

	-- like a combinational circuit..
	-- the control path must worry about all
	-- sequencing issues.
     flowThrough: if (flow_through) generate
	z <= ilb_data_in;
    	sample_ack <= sample_req;
    	update_ack <= update_req;

     end generate flowThrough;
end arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- Assumption: guard-interface will not change until
-- sr_in -> sa_out sequence has completed.
--
entity SgiSampleFsm is
	generic (name: string);
	port (sr_in: in Boolean;
		sr_in_q: out Boolean;
		push_req: out std_logic;
		push_ack: in std_logic;
		clk, reset: in std_logic);
end entity;

architecture BehaviouralFsm of SgiSampleFsm is
	type SrInState is (Idle, WaitOnPushAck);
	signal sr_in_state: SrInState;

	signal sr_in_q_sig: Boolean;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

	sr_in_q <= sr_in_q_sig;

	process(sr_in_state, sr_in, push_ack, clk, reset)
		variable next_sr_in_state: SrInState;
		variable sr_in_q_var: Boolean;
		variable push_req_var: std_logic;
	begin
		sr_in_q_var := false;
		next_sr_in_state := sr_in_state;
		push_req_var := '0';

		case sr_in_state is
			when Idle =>
				if (sr_in) then
					push_req_var := '1';
					if(push_ack = '1') then
						sr_in_q_var := true;
					else
						next_sr_in_state := WaitOnPushAck;
					end if;
				end if;
			when WaitOnPushAck =>
				push_req_var := '1';
				if(push_ack = '1') then
					sr_in_q_var := true;
					next_sr_in_state := Idle;
				end if;
		end case;

		push_req <= push_req_var;
		sr_in_q_sig  <= sr_in_q_var;

		if (clk'event and clk = '1') then
			if(reset = '1') then
				sr_in_state <= Idle;
			else
				sr_in_state <= next_sr_in_state;
			end if;
		end if;
	end process;
end BehaviouralFsm;
	
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.Types.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- Assumption: guard-interface will not change until
-- sr_in -> sa_out sequence has completed.
--
entity SgiUpdateFsm is
	generic (name: string);
	port (cr_in: in Boolean;
		cr_out: out Boolean;
		ca_in: in Boolean;
		ca_out: out Boolean;
		pop_req: out std_logic;
		pop_ack: in std_logic;
		pop_data: in std_logic_vector(0 downto 0);
		clk, reset: in std_logic);
end entity;

architecture BehaviouralFsm of SgiUpdateFsm is

	type UpdateFsmState is (UpdateFsmRun, UpdateFsmWaitPop, UpdateFsmWaitCain);
	signal update_fsm_state: UpdateFsmState;

	signal ca_out_d, ca_out_u: boolean;

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

	process(clk, reset, pop_ack, cr_in, ca_in, pop_data, update_fsm_state)
		variable next_update_fsm_state_var: UpdateFsmState;
		variable pop_req_var : std_logic;
		variable cr_out_var, ca_out_d_var, ca_out_u_var: boolean;
	begin
		next_update_fsm_state_var := update_fsm_state;
		pop_req_var := '0';
		cr_out_var := false;
		ca_out_d_var := false;
		ca_out_u_var := false;

		case update_fsm_state is
			when UpdateFsmRun =>
				if(cr_in) then
					pop_req_var := '1';
					if(pop_ack = '1') then
						if(pop_data(0) = '0') then
							ca_out_d_var := true;
						else
							cr_out_var := true;
							next_update_fsm_state_var := UpdateFsmWaitCain;
						end if;
					else
						next_update_fsm_state_var := UpdateFsmWaitPop;
					end if;
				end if;
			when UpdateFsmWaitPop =>
				pop_req_var := '1';
				if(pop_ack = '1') then
					if(pop_data(0) = '0') then
						ca_out_d_var := true;
						next_update_fsm_state_var := UpdateFsmRun;
					else
						cr_out_var := true;
						next_update_fsm_state_var := UpdateFsmWaitCain;
					end if;
				end if;
			when UpdateFsmWaitCain =>
				if(ca_in) then
					ca_out_u_var := true;
					if(cr_in) then 
						pop_req_var := '1';
						if(pop_ack = '1') then
							if(pop_data(0) = '0') then
								ca_out_d_var := true;
								next_update_fsm_state_var := UpdateFsmRun;
							else
								cr_out_var := true;
							end if;
						else
							next_update_fsm_state_var := UpdateFsmWaitPop;
						end if;
					else
						next_update_fsm_state_var := UpdateFsmRun;
					end if;
				end if;
		end case;

		ca_out_u <= ca_out_u_var;
		cr_out   <= cr_out_var;
		pop_req  <= pop_req_var;

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				ca_out_d <= false;
				update_fsm_state <= UpdateFsmRun;
			else
				ca_out_d <= ca_out_d_var;
				update_fsm_state <= next_update_fsm_state_var;
			end if;
		end if;
	end process;

	ca_out <= ca_out_d or ca_out_u;
end BehaviouralFsm;
	
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

--
-- base Pipe.
--  in all cases, we will go for an implementation which
--  gives a throughput of one word/cycle.
--

entity SignalBase is
  generic (name : string;
	   volatile_flag: boolean := false;
           num_writes: integer;
           data_width: integer);
  port (
    read_data      : out std_logic_vector(data_width-1 downto 0);
    write_req       : in  std_logic_vector(num_writes-1 downto 0);
    write_ack       : out std_logic_vector(num_writes-1 downto 0);
    write_data      : in std_logic_vector((num_writes*data_width)-1 downto 0);
    clk, reset : in  std_logic);
  
end SignalBase;

architecture default_arch of SignalBase is

  signal pipe_data, read_data_reg: std_logic_vector(data_width-1 downto 0);
  signal pipe_req, pipe_ack: std_logic;
  
begin  -- default_arch


  manyWriters: if (num_writes > 1) generate
    wmux : OutputPortLevel generic map (
      name => name & "-wmux",
      num_reqs       => num_writes,
      data_width     => data_width,
      no_arbitration => false)
      port map (
        req   => write_req,
        ack   => write_ack,
        data  => write_data,
        oreq  => pipe_req,                -- no cross-over, drives req
        oack  => pipe_ack,                -- no cross-over, receives ack
        odata => pipe_data,
        clk   => clk,
        reset => reset);
  end generate manyWriters;

  singleWriter: if (num_writes = 1) generate
    pipe_req <= write_req(0);
    write_ack(0) <= pipe_ack;
    pipe_data <= write_data;
  end generate singleWriter;
 
  -- in signal mode, the pipe is just a flag
  -- write always succeeds.
  pipe_ack <= '1';

  -- in volatile-mode, the signal follws the input
  -- as long as the request is maintained else
  -- it shows a blank (0)
  VolatileGen: if volatile_flag generate
	read_data <= pipe_data when pipe_req = '1' else (others => '0');
  end generate VolatileGen;

  -- in non-volatile mode, the signal is a flag, 
  -- set by pipe-reg.
  nonVolatileGen: if not volatile_flag generate
     process(clk,reset) 
     begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			read_data_reg <= (others => '0');	
		else
			if(pipe_req = '1') then
				read_data_reg <= pipe_data;
			end if;
		end if;
	end if;
     end process;

     read_data <= read_data_reg;
  end generate nonVolatileGen;


end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library ahir;
use ahir.Utilities.all;
use ahir.SubPrograms.all;

--
-- a special purpose queue which keeps a 1-bit data value.
--
entity SingleBitQueueBase is
  generic(name : string; queue_depth: integer := 1; bypass_flag: boolean := false);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(0 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(0 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity SingleBitQueueBase;

architecture behave of SingleBitQueueBase is

  function rotate_left(x: std_logic_vector) return std_logic_vector is
	alias lx: std_logic_vector(1 to x'length) is x;
	variable ret_val : std_logic_vector(1 to x'length);
  begin
	ret_val(1 to x'length-1)  := lx(2 to x'length);
	ret_val (x'length) := lx(1);
	return(ret_val);
  end rotate_left;


begin  -- SimModel

 --
 -- 0-depth queue is just a set of wires.
 --
 triv: if queue_depth = 0 generate
	push_ack <= pop_req;
	pop_ack  <= push_req;
	data_out <= data_in;
 end generate triv;



 qDGt0: if queue_depth > 0 generate 
  NTB: block 
  	signal queue_vector: std_logic_vector(queue_depth-1 downto 0);
  	signal write_pointer, incr_write_pointer: std_logic_vector(queue_depth-1 downto 0);
  	signal read_pointer, incr_read_pointer: std_logic_vector(queue_depth-1 downto 0);
     	signal queue_size : unsigned ((Ceil_Log2(queue_depth+1))-1 downto 0);
	signal empty_flag, bypass_active : boolean := false;
	signal actual_push_req: std_logic;
  begin

 
    assert (queue_size < queue_depth) report "Queue " & name & " is full." severity note;
    assert (queue_size < (3*queue_depth/4)) report "Queue " & name & " is three-quarters-full." severity note;
    assert (queue_size < (queue_depth/2)) report "Queue " & name & " is half-full." severity note;
    assert (queue_size < (queue_depth/4)) report "Queue " & name & " is quarter-full." severity note;

    qD1: if (queue_depth = 1) generate
     incr_read_pointer <= read_pointer;
     incr_write_pointer <= write_pointer;
    end generate qD1;

    byp_gen: if bypass_flag generate

	empty_flag <= (queue_size = 0);
	bypass_active <= (empty_flag and (push_req = '1'));

	actual_push_req <= '0' when (bypass_active and (pop_req = '1')) else push_req;
    	pop_ack  <= '1' when ((queue_size > 0) or bypass_active) else '0';

    	data_out(0) <= data_in(0) when bypass_active else
				OrReduce (queue_vector and read_pointer);
    end generate byp_gen;

    no_byp_gen: if not bypass_flag generate

	bypass_active <= false;
	actual_push_req <= push_req;
    	pop_ack  <= '1' when (queue_size > 0) else '0';
    
	-- bottom pointer gives the data in FIFO mode..
    	data_out(0) <= OrReduce (queue_vector and read_pointer);

    end generate no_byp_gen;

    qDG1: if (queue_depth > 1) generate
     incr_read_pointer <= rotate_left(read_pointer);
     incr_write_pointer <= rotate_left(write_pointer);
    end generate qDG1;

    push_ack <= '1' when (queue_size < queue_depth) else '0';

  
    -- single process
    process(clk, reset, read_pointer, write_pointer, incr_read_pointer, incr_write_pointer, queue_size, 
			actual_push_req, pop_req)
      variable qsize : unsigned ((Ceil_Log2(queue_depth+1))-1 downto 0);
      variable push,pop : boolean;
      variable next_read_ptr,next_write_ptr : std_logic_vector(queue_depth-1 downto 0);
    begin

      qsize := queue_size;
      push  := false;
      pop   := false;
      next_read_ptr := read_pointer;
      next_write_ptr := write_pointer;
      
      if((qsize < queue_depth) and (actual_push_req = '1')) then
          push := true;
      end if;
  
      if((qsize > 0) and (pop_req = '1') and (not bypass_active)) then
          pop := true;
      end if;
  
  
      if(push) then
          next_write_ptr := incr_write_pointer;
      end if;
  
      if(pop) then
          next_read_ptr := incr_read_pointer;
      end if;
  
  
      -- queue size modified only in non-bypass case
      if(pop and (not push)) then
          qsize := qsize - 1;
      elsif(push and (not pop)) then
          qsize := qsize + 1;
      end if;
        
  
      if(clk'event and clk = '1') then
        
	if(reset = '1') then
           queue_size <= (others => '0');
           read_pointer <= (0 => '1', others => '0');
           write_pointer <= (0 => '1', others => '0');
           queue_vector <= (others => '0'); -- initially 0.
	else
           if(push) then
		if(data_in(0) = '1') then
			queue_vector <= queue_vector or write_pointer;
		else
			queue_vector <= queue_vector and (not write_pointer);
		end if;
           end if;
        
           queue_size <= qsize;
           read_pointer <= next_read_ptr;
           write_pointer <= next_write_ptr;

        end if;
      end if;

    end process;
   end block NTB;
  end generate qDGt0;
  

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.Utilities.all;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;

-- a simple slicing element.
entity SliceSplitProtocol is
  generic(name: string; 
	in_data_width : integer; 
	high_index: integer; 
	low_index : integer; 
	buffering : integer;
	flow_through: boolean := false;
	full_rate: boolean := false
	);
  port(din: in std_logic_vector(in_data_width-1 downto 0);
       dout: out std_logic_vector(high_index-low_index downto 0);
       sample_req: in boolean;
       sample_ack: out boolean;
       update_req: in boolean;
       update_ack: out boolean;
       clk,reset: in std_logic);
end SliceSplitProtocol;


architecture arch of SliceSplitProtocol is
   signal ilb_data_in: std_logic_vector(high_index-low_index downto 0);
begin

  assert ((high_index < in_data_width) and (low_index >= 0) and (high_index >= low_index))
    report "inconsistent slice parameters" severity failure;
  
  noFlowThrough: if (not flow_through) generate

    ilb_data_in <= din(high_index downto low_index);
    ilb: InterlockBuffer 
		generic map(name => name & "-ilb",
				buffer_size => buffering,
				in_data_width => (high_index - low_index) + 1,
				out_data_width => (high_index - low_index) + 1)
		port map(write_req => sample_req,
			 write_ack => sample_ack,
			 write_data => ilb_data_in,
			 read_req  => update_req,
			 read_ack => update_ack,
			 read_data => dout,
			 clk => clk, reset => reset);

  end generate noFlowThrough;

  flowThrough: if flow_through generate
    dout <= din(high_index downto low_index);
    sample_ack <= sample_req;
    update_ack <= update_req;
  end generate flowThrough;
  
end arch;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##


-- a guard-interface to conform with the split protocol.
-- With this interface, the guard at the time of initiation
-- of the operation will be remembered (using a queue) 
-- and the remembered value will be used to generate the
-- completion protocol.
-- 
-- The benefit is that the guard-expression can be reevaluated
-- as soon as the operation starts (instead of waiting
-- for the operation to finish...).  This helps pipelining.
--
-- Assumptions
--   1. sr_in -> sr_in without intervening sa_out is not possible.
--   2. cr_in -> cr_in without intervening ca_out is not possible.
--
entity SplitGuardInterfaceBase is
	generic (name: string; buffering:integer);
	port (sr_in: in Boolean;
	      sa_out: out Boolean;
	      sr_out: out Boolean;
	      sa_in: in Boolean;
	      cr_in: in Boolean;
	      ca_out: out Boolean;
	      cr_out: out Boolean;
	      ca_in: in Boolean;
	      guard_interface: in std_logic;
	      clk: in std_logic;
	      reset: in std_logic);
end entity;


architecture Behave of SplitGuardInterfaceBase is
  signal push, push_ack, pop, pop_ack: std_logic;
  signal qdata_in, qdata : std_logic_vector(0 downto 0);

  type RhsState is (r_Idle, r_Wait_On_Ack_In, r_Wait_On_Queue);
  signal rhs_state: RhsState;

  -- for debug purposes only
  signal s_counter, c_counter: integer;

  -- number of stages!  This will cause
  -- the minimum latency of sr -> ca to
  -- increase to this number...  Be careful..
  constant g_queue_number_of_stages : integer := Ceil(buffering, max_single_bit_queue_depth_per_stage);

  -- constant g_queue_number_of_stages : integer := 1;
 
  signal sr_in_q : Boolean;
  signal guard_interface_sustained, guard_interface_registered: std_logic;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin
	qdata_in(0) <= guard_interface;

	qI: ShiftRegisterSingleBitQueue  -- bypass to maintain delays
		generic map(name => name & "-qI", 
					queue_depth => buffering, 
					number_of_stages => g_queue_number_of_stages,
					bypass_flag => true
			   )
		port map(clk => clk, reset => reset,
				data_in => qdata_in,
				push_req => push,
				push_ack => push_ack,
				data_out => qdata,
				pop_req => pop,
				pop_ack => pop_ack);

	-----------------------------------------------------------------------------------------------
	-- sample side logic.
	-----------------------------------------------------------------------------------------------
	sampleFsm: SgiSampleFsm
			generic map (name => name & "-sample-fsm")
			port map (clk => clk, reset => reset,
					sr_in => sr_in, sr_in_q => sr_in_q,
					push_req => push, push_ack => push_ack);


	-- Race condition in PHI statements can be an issue!
	process(clk, reset, guard_interface, sr_in)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				guard_interface_registered <= '0';
			elsif(sr_in) then
				guard_interface_registered <= guard_interface;
			end if;
		end if;
	end process;
	guard_interface_sustained <= guard_interface when sr_in else guard_interface_registered;

	-- sr_out
	sr_out <= sr_in_q when (guard_interface_sustained = '1') else false;
	
	-- sa_out
	sa_out <= sr_in_q when (guard_interface_sustained = '0') else sa_in;

	-----------------------------------------------------------------------------------------------
	-- update side logic.
	-----------------------------------------------------------------------------------------------
	updateFsm: SgiUpdateFsm
			generic map 
				 (name => name & "-update-fsm")
			port map (clk => clk,
					reset => reset,
					cr_in => cr_in,
					cr_out => cr_out,
					ca_in => ca_in,
					ca_out => ca_out,
					pop_req => pop,
					pop_ack => pop_ack,
					pop_data => qdata);

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity SplitGuardInterface is
	generic (name: string; nreqs: integer; buffering:IntegerArray; use_guards: BooleanArray; 
			sample_only: Boolean; update_only: Boolean);
	port (sr_in: in BooleanArray(nreqs-1 downto 0);
	      sa_out: out BooleanArray(nreqs-1 downto 0); 
	      sr_out: out BooleanArray(nreqs-1 downto 0);
	      sa_in: in BooleanArray(nreqs-1 downto 0); 
	      cr_in: in BooleanArray(nreqs-1 downto 0);
	      ca_out: out BooleanArray(nreqs-1 downto 0); 
	      cr_out: out BooleanArray(nreqs-1 downto 0);
	      ca_in: in BooleanArray(nreqs-1 downto 0); 
	      guards: in std_logic_vector(nreqs-1 downto 0);
	      clk: in std_logic;
	      reset: in std_logic);
end entity;


architecture Behave of SplitGuardInterface is
	constant gFlags: BooleanArray(nreqs-1 downto 0) := use_guards;
	constant gBufs: IntegerArray(nreqs-1 downto 0) := buffering;
begin
	BaseGen: for I in nreqs-1 downto 0 generate

	     gCase: if gFlags(I) generate
		SampleOnly: if sample_only generate
		   sgis: SplitSampleGuardInterfaceBase
			generic map (name => name & "-gCase-SampleOnly-sgis-" & Convert_To_String(I), buffering => gBufs(I))
			port map(sr_in => sr_in(I),
				 sr_out => sr_out(I),
				 sa_in => sa_in(I),
				 sa_out => sa_out(I),
				 cr_in => cr_in(I),
				 cr_out => cr_out(I),
				 ca_in => ca_in(I),
				 ca_out => ca_out(I),
				 guard_interface => guards(I),
				 clk => clk, reset => reset);
		end generate SampleOnly;

		UpdateOnly: if update_only generate
		   sgiu: SplitUpdateGuardInterfaceBase
			generic map (name => name & "-gCase-UpdateOnly-sgiu-" & Convert_To_String(I), buffering => gBufs(I))
			port map(sr_in => sr_in(I),
				 sr_out => sr_out(I),
				 sa_in => sa_in(I),
				 sa_out => sa_out(I),
				 cr_in => cr_in(I),
				 cr_out => cr_out(I),
				 ca_in => ca_in(I),
				 ca_out => ca_out(I),
				 guard_interface => guards(I),
				 clk => clk, reset => reset);
		end generate UpdateOnly;

		SampleAndUpdate: if (not (sample_only or update_only)) generate
		   sgi: SplitGuardInterfaceBase
			generic map (name => name & "-gCase-SampleAndUpdate-sgiu-" & Convert_To_String(I), buffering => gBufs(I))
			port map(sr_in => sr_in(I),
				 sr_out => sr_out(I),
				 sa_in => sa_in(I),
				 sa_out => sa_out(I),
				 cr_in => cr_in(I),
				 cr_out => cr_out(I),
				 ca_in => ca_in(I),
				 ca_out => ca_out(I),
				 guard_interface => guards(I),
				 clk => clk, reset => reset);
		end generate SampleAndUpdate;

              end generate gCase;
	   
 	      noG: if not gFlags(I) generate
		 sr_out(I) <= sr_in(I);
		 sa_out(I) <= sa_in(I);
		 cr_out(I) <= cr_in(I);
		 ca_out(I) <= ca_in(I);
              end generate noG;
        end generate;

end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- A half guard interface which forwards only
-- the sample.  (used on output ports).
--  Madhav P. Desai.
entity SplitSampleGuardInterfaceBase is
	generic (name: string; buffering:integer);
	port (sr_in: in Boolean;
	      sa_out: out Boolean;
	      sr_out: out Boolean;
	      sa_in: in Boolean;
	      cr_in: in Boolean;
	      ca_out: out Boolean;
	      cr_out: out Boolean;
	      ca_in: in Boolean;
	      guard_interface: in std_logic;
	      clk: in std_logic;
	      reset: in std_logic);
end entity;


architecture Behave of SplitSampleGuardInterfaceBase is
	Type FsmState is (Idle, Busy);
	signal fsm_state: FsmState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

	-- cr/ca interface is a dummy... no need to forward to the
	-- operator which does not care anyway.
	cr_out <= false;
	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				ca_out <= false;
			else
				ca_out <= cr_in;
			end if;
		end if;
	end process;


	-- sample guard FSM.
	process(clk, guard_interface, fsm_state, sr_in, sa_in)
		variable next_state : FsmState;
		variable sr_out_var, sa_out_var: Boolean;
	begin
		next_state := fsm_state;
		sr_out_var := false;
		sa_out_var := false;
		case fsm_state is
			when Idle =>
				if(sr_in) then
					if(guard_interface  = '1') then
						sr_out_var := true;
						if(sa_in) then
							sa_out_var := true;
						else
							next_state := Busy;
						end if;
					else
						-- give ack, since guard is 0.
						sa_out_var := true;	
					end if;
				end if;
			when Busy => 
				if(sa_in) then
					next_state := Idle;
					sa_out_var := true;
				end if;
		end case;
		
		sr_out <= sr_out_var;
		sa_out <= sa_out_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= Idle;
			else 
				fsm_state <= next_state;
			end if;
		end if;
	end process;	
	
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##


-- A half guard interface which forwards only
-- the update.  (used on input ports).
--  Madhav P. Desai.
entity SplitUpdateGuardInterfaceBase is
	generic (name: string; buffering:integer);
	port (sr_in: in Boolean;
	      sa_out: out Boolean;
	      sr_out: out Boolean;
	      sa_in: in Boolean;
	      cr_in: in Boolean;
	      ca_out: out Boolean;
	      cr_out: out Boolean;
	      ca_in: in Boolean;
	      guard_interface: in std_logic;
	      clk: in std_logic;
	      reset: in std_logic);
end entity;


architecture Behave of SplitUpdateGuardInterfaceBase is
	Type FsmState is (Idle, Busy);
	signal fsm_state: FsmState;
	signal ca_out_u, ca_out_d: Boolean;
	signal guard_interface_reg, sampled_guard_interface: std_logic;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin
	sa_out <= sr_in;
	sr_out <= false;
		
	-- sr/sa interface is a dummy... no need to forward to the
	process (clk, reset, sr_in)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				guard_interface_reg <= '0';
			elsif sr_in then
				guard_interface_reg <= guard_interface;
			end if;
		end if;
	end process;
	sampled_guard_interface <= guard_interface when sr_in else guard_interface_reg;


	-- update guard FSM.
	process(clk, sampled_guard_interface, fsm_state, cr_in, ca_in)
		variable next_state : FsmState;
		variable cr_out_var, ca_out_var_d, ca_out_var_u: Boolean;
	begin
		next_state := fsm_state;
		cr_out_var := false;
		ca_out_var_u := false;
		ca_out_var_d := false;
		case fsm_state is
			when Idle =>
				if(cr_in) then
					if(sampled_guard_interface  = '1') then
						cr_out_var := true;
						next_state := Busy;
					else
						-- give delayed ack, since guard is 0.
						ca_out_var_d := true;	
					end if;
				end if;
			when Busy => 
				if(ca_in) then
					ca_out_var_u := true;
					if(cr_in) then
						if(sampled_guard_interface = '1') then
							cr_out_var := true;
						else
							ca_out_var_d := true;
							next_state := Idle;
						end if;
					else
						next_state := Idle;
					end if;
				end if;
		end case;
		
		cr_out <= cr_out_var;
		ca_out_u <= ca_out_var_u;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= Idle;
				ca_out_d <= false;
			else 
				fsm_state <= next_state;
				ca_out_d <= ca_out_var_d;
			end if;
		end if;
	end process;	
	ca_out <= ca_out_u or ca_out_d;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;

entity StoreReqSharedWithInputBuffers is
    generic
    (
	name : string;
	addr_width: integer;
	data_width : integer;
	time_stamp_width : integer;
      	num_reqs : integer; -- how many requesters?
	tag_length: integer;
	no_arbitration: Boolean := false;
        min_clock_period: Boolean := true;
	input_buffering: IntegerArray
    );
  port (
    -- req/ack follow pulse protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    -- address corresponding to access
    addr                    : in std_logic_vector((addr_width*num_reqs)-1 downto 0);
    data                    : in std_logic_vector((data_width*num_reqs)-1 downto 0);
    -- address to memory
    maddr                   : out std_logic_vector(addr_width-1 downto 0);
    mdata                   : out std_logic_vector(data_width-1 downto 0);
    mtag                    : out std_logic_vector(tag_length+time_stamp_width-1 downto 0);
    mreq                    : out std_logic;
    mack                    : in std_logic;
    -- clock, reset (active high)
    clk, reset              : in std_logic);
end StoreReqSharedWithInputBuffers;

architecture Vanilla of StoreReqSharedWithInputBuffers is

  constant iwidth: integer := addr_width*num_reqs;
  constant owidth: integer := addr_width;

  constant debug_flag : boolean := global_debug_flag;

  -- must register..  ack implies that address has been sampled.
  constant registered_output : boolean := true; 

  type TagWordArray is array (natural range <>) of unsigned(tag_length-1 downto 0);
  signal rx_tag_in: TagWordArray(num_reqs-1 downto 0);

  constant rx_word_length: integer := addr_width + data_width + tag_length + time_stamp_width;
  type RxBufWordArray is array (natural range <>) of std_logic_vector(rx_word_length-1 downto 0);

  signal rx_data_in, rx_data_out : RxBufWordArray(num_reqs-1 downto 0);

  signal imux_data_in_accept,  imux_data_in_valid: std_logic_vector(num_reqs-1 downto 0);
  signal imux_data_in: std_logic_vector((rx_word_length*num_reqs)-1 downto 0);

  signal imux_data_out_accept,  imux_data_out_valid: std_logic;
  signal imux_data_out: std_logic_vector(rx_word_length-1 downto 0);
  
  -- alias IBUFs: IntegerArray(num_reqs-1 downto 0) is input_buffering;
begin  -- Behave
  assert(tag_length >= Ceil_Log2(num_reqs)) report "insufficient tag width" severity error;
 

  tagGen: for I in 0 to num_reqs-1 generate
	rx_tag_in(I) <= To_Unsigned(I,tag_length);	
  end generate tagGen;


  TstampGen: if time_stamp_width > 0 generate
	Tsb: block 
		signal time_stamp: std_logic_vector(time_stamp_width-1 downto 0);
	begin
		tsc: CounterBase generic map(name => name & "-TstampGen->Tsb-tsc", data_width => time_stamp_width)
			port map(clk => clk, reset => reset, count_out => time_stamp);

		rxInDataGen: for I in 0 to num_reqs-1 generate
			rx_data_in(I) <= addr(((I+1)*addr_width)-1 downto I*addr_width) &
					 data(((I+1)*data_width)-1 downto I*data_width)  &  std_logic_vector(rx_tag_in(I)) & time_stamp;
		end generate rxInDataGen;
	end block Tsb;
  end generate TstampGen;

  NoTstampGen: if time_stamp_width < 1 generate
	rxInDataGen: for I in 0 to num_reqs-1 generate
		rx_data_in(I) <= addr(((I+1)*addr_width)-1 downto I*addr_width)  &
					 data(((I+1)*data_width)-1 downto I*data_width) & std_logic_vector(rx_tag_in(I));
	end generate rxInDataGen;
  end generate NoTstampGen;

  -- receive buffers.
  RxGen: for I in 0 to num_reqs-1 generate
	rb: ReceiveBuffer generic map(name => name & "-rb " & Convert_To_String(I),
					buffer_size => Maximum(2,input_buffering(I)),
					data_width => rx_word_length,
					full_rate => false) -- double buffered.. automatically full-rate.
		port map(write_req => reqL(I), 
			 write_ack => ackL(I), 
			 write_data => rx_data_in(I), 
			 read_req => imux_data_in_accept(I), 
			 read_ack => imux_data_in_valid(I), 
                         read_data => rx_data_out(I),
			 clk => clk, 
			 reset => reset);

  end generate RxGen;

  -- data for input mux.
  process(rx_data_out)
  begin
	for I in 0 to num_reqs-1 loop
		imux_data_in(((I+1)*rx_word_length)-1 downto (I*rx_word_length))
			<= rx_data_out(I);
	end loop;
  end process;

  -- the multiplexor.
  NonTrivTstamp: if time_stamp_width > 0 generate
  	imux: merge_tree
    	   generic map(name => name & "-NonTrivTstamp-imux", g_number_of_inputs => num_reqs,
		g_data_width => rx_word_length,
                g_time_stamp_width => time_stamp_width, 
                g_tag_width => tag_length,
		g_mux_degree => 4096, -- some large number.. allow big muxes.
		g_num_stages => 1,    -- with single stage delay 
		g_port_id_width => 0)
           port map(merge_data_in => imux_data_in,
	            merge_req_in  => imux_data_in_valid,
	            merge_ack_out => imux_data_in_accept,
	            merge_data_out => imux_data_out,
                    merge_req_out => imux_data_out_valid,
	            merge_ack_in  => imux_data_out_accept,
      	            clock        => clk,
      	            reset      => reset);
  end generate NonTrivTstamp;

  TrivTstamp: if time_stamp_width < 1 generate
	imux: LevelMux generic map (name => name & "-TrivTstamp-imux", 
				num_reqs => num_reqs, data_width => rx_word_length, no_arbitration => false)
		port map(write_req => imux_data_in_valid,
			 write_ack => imux_data_in_accept,
			 write_data => imux_data_in,
			 read_req => imux_data_out_accept,
		         read_ack => imux_data_out_valid,
			 read_data => imux_data_out,
			 clk => clk, reset => reset);
  end generate TrivTstamp;


  -- outgoing tag, address, data
  mreq <= imux_data_out_valid;
  imux_data_out_accept <= mack;
  maddr <= imux_data_out(rx_word_length-1 downto (data_width + tag_length + time_stamp_width));
  mdata <= imux_data_out((rx_word_length - addr_width)-1 downto (tag_length + time_stamp_width));
  mtag <= imux_data_out(tag_length+time_stamp_width-1 downto 0);

end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- 
--  whatever appears at in_data is
--  read by whoever wishes to read it.
--
--
entity SystemInPort is
   generic (name : string;
	    num_reads: integer;
	    in_data_width: integer;
            out_data_width : integer; 
	    full_rate: boolean);
   port (read_req : in std_logic_vector(num_reads-1 downto 0);
         read_ack : out std_logic_vector(num_reads-1 downto 0);
         read_data: out std_logic_vector((num_reads*out_data_width)-1 downto 0);
         in_data  : in std_logic_vector(in_data_width-1 downto 0);
	 clk : in std_logic;
	 reset : in std_logic);
end entity;

architecture Mixed of SystemInPort is

    constant min_width : integer := Minimum(in_data_width, out_data_width);
    signal data_reg, tr_p_in_data: std_logic_vector(min_width-1 downto 0);
    signal tr_data : std_logic_vector(out_data_width-1 downto 0);
    signal valid_data : std_logic;
begin

    -- stored data will be of minimum width.
    TruncateOrPad(in_data, tr_p_in_data); 
    process(clk)
    begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			data_reg <= (others => '0');
			valid_data <= '0';
		else
			data_reg <= tr_p_in_data;
			valid_data <= '1';
		end if;
	end if;
    end process;


    -- pad out data_reg..
    TruncateOrPad(data_reg, tr_data);

    -- padded data is broadcast to all readers.
    ReadGen: for I in 0 to num_reads-1 generate

      read_ack(I) <= valid_data;
      process(tr_data)
      begin
	read_data(((I+1)*out_data_width)-1 downto I*out_data_width) <= tr_data;
      end process;
    end generate ReadGen;
end Mixed;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

--
-- Last successful write wins.
--
entity SystemOutPort is
   generic (name : string;
	    num_writes: integer;
	    in_data_width: integer;
            out_data_width : integer;
	    full_rate: boolean := false); 
   port (write_req : in std_logic_vector(num_writes-1 downto 0);
         write_ack : out std_logic_vector(num_writes-1 downto 0);
         write_data: in std_logic_vector((num_writes*in_data_width)-1 downto 0);
         out_data  : out std_logic_vector(out_data_width-1 downto 0);
	 clk : in std_logic;
	 reset : in std_logic);
end entity;

architecture Mixed of SystemOutPort is
    constant min_width : integer := Minimum(in_data_width, out_data_width);
    
    signal read_req, read_ack: std_logic_vector(0 downto 0);
    signal pipe_data_in: std_logic_vector((num_writes*min_width)-1 downto 0);
    signal pipe_data_out: std_logic_vector(min_width-1 downto 0);
    signal out_reg: std_logic_vector(min_width-1 downto 0);
    
begin

    -- keep only the necessary bits of write_data.
    wPadTrunc: for I in 0 to num_writes-1 generate
		-- signal arguments.
	TruncateOrPad(write_data(((I+1)*in_data_width)-1 downto I*in_data_width), 
					pipe_data_in((I+1)*min_width-1 downto I*min_width));
    end generate wPadTrunc;

    read_req(0) <= '1';

    -- data coming from pipe..
    TruncateOrPad(pipe_data_out, out_data);

    --
    -- pipe.. to provide interlock so only one writer succeeds at a time.
    --
    opipe: PipeBase generic map(name => name & "-opipe", 
				    num_reads => 1,
					num_writes => num_writes, data_width => min_width,
						lifo_mode => false, signal_mode => true, depth => 1, full_rate => full_rate)
		port map(read_req => read_req, read_ack => read_ack,
				read_data => pipe_data_out,
					write_req => write_req, write_ack => write_ack,
						write_data => pipe_data_in,
							clk => clk, reset => reset);

end Mixed;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;
-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

--  
--
-- A more "optimized" version of the old UnloadBuffer.
-- tries to avoid the use of an extra register.  Use
-- when buffer-size > 1.
--  
--
entity UnloadBufferRevisedNonblocking is

  generic (name: string; 
		buffer_size: integer ; 
		data_width : integer ; 
		bypass_flag: boolean );

  port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);

end UnloadBufferRevisedNonblocking;

architecture default_arch of UnloadBufferRevisedNonblocking is

  signal pop_req, pop_ack, push_req, push_ack: std_logic_vector(0 downto 0);

  signal pipe_data_out, ufsm_bypass_write_data, ufsm_write_data:  std_logic_vector(data_width-1 downto 0);
  signal pipe_has_data: boolean;


  signal write_to_pipe: boolean;
  signal unload_from_pipe : boolean;

  signal empty, full: std_logic;
  signal ufsm_write_req, ufsm_write_ack: std_logic;
  signal ufsm_bypass_write_req, ufsm_bypass_write_ack: std_logic;

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch

	ufsm_write_data <= pipe_data_out;
	ufsm_write_req  <= pop_ack(0);
	pop_req(0) <= ufsm_write_ack;

	push_req(0) <= write_req;
	write_ack   <= push_ack(0);

	ufsm: UnloadFsmNoblock generic map (name => name & ":ufsm", data_width => data_width)
		port map (
			   write_req => ufsm_write_req,
			   write_ack => ufsm_write_ack,
			   unload_req => unload_req,
			   unload_ack => unload_ack,
			   data_in => ufsm_write_data,
			   data_out => read_data,
			   clk => clk, reset => reset);

  	pipe_has_data <= (empty = '0');
  	has_data <= '1' when pipe_has_data else '0';


  	bufPipe : QueueBaseWithEmptyFull generic map (
        	name =>  name & "-blocking_read-bufPipe",
        	data_width => data_width,
		reverse_bypass_flag => bypass_flag,
        	queue_depth      => buffer_size)
      	port map (
        	pop_req   => pop_req(0),
        	pop_ack   => pop_ack(0),
        	data_out  => pipe_data_out,
        	push_req  => push_req(0),
        	push_ack  => push_ack(0),
        	data_in => write_data,
		empty => empty,
		full => full,
        	clk        => clk,
        	reset      => reset);

	
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.GlobalConstants.all;
-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

--  
--
-- A more "optimized" version of the old UnloadBuffer.
-- tries to avoid the use of an extra register.  Use
-- when buffer-size > 1.
--  
--
entity UnloadBufferRevised is

  generic (name: string; 
		buffer_size: integer ; 
		data_width : integer ; 
		bypass_flag: boolean );

  port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
	has_data: out std_logic;
        clk : in std_logic;
        reset: in std_logic);

end UnloadBufferRevised;

architecture default_arch of UnloadBufferRevised is

  signal pop_req, pop_ack, push_req, push_ack: std_logic_vector(0 downto 0);

  signal pipe_data_out, ufsm_bypass_write_data, ufsm_write_data:  std_logic_vector(data_width-1 downto 0);
  signal pipe_has_data: boolean;


  signal write_to_pipe: boolean;
  signal unload_from_pipe : boolean;

  signal empty, full: std_logic;
  signal ufsm_write_req, ufsm_write_ack: std_logic;
  signal ufsm_bypass_write_req, ufsm_bypass_write_ack: std_logic;

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch

	ufsm_write_data <= pipe_data_out;
	ufsm_write_req  <= pop_ack(0);
	pop_req(0) <= ufsm_write_ack;

	push_req(0) <= write_req;
	write_ack   <= push_ack(0);

	ufsm: UnloadFsm generic map (name => name & ":ufsm", data_width => data_width)
		port map (
			   write_req => ufsm_write_req,
			   write_ack => ufsm_write_ack,
			   unload_req => unload_req,
			   unload_ack => unload_ack,
			   data_in => ufsm_write_data,
			   data_out => read_data,
			   clk => clk, reset => reset);

  	pipe_has_data <= (empty = '0');
  	has_data <= '1' when pipe_has_data else '0';


  	bufPipe : QueueBaseWithEmptyFull generic map (
        	name =>  name & "-blocking_read-bufPipe",
        	data_width => data_width,
		reverse_bypass_flag => bypass_flag,
        	queue_depth      => buffer_size)
      	port map (
        	pop_req   => pop_req(0),
        	pop_ack   => pop_ack(0),
        	data_out  => pipe_data_out,
        	push_req  => push_req(0),
        	push_ack  => push_ack(0),
        	data_in => write_data,
		empty => empty,
		full => full,
        	clk        => clk,
        	reset      => reset);

	
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

--  A non-blocking version of the state machine for
--  handling the revised case of the unload-buffer.
--
-- BUG ALERT:  there is something wrong about this 
--             which causes incorrect behaviour. 
--             Am stymied for the moment (MPD)
--
entity UnloadFsmNoBlock is
  generic (name: string; data_width: integer);
  port ( 
	 write_req: in std_logic;
         write_ack: out std_logic;
         unload_req: in boolean;
         unload_ack: out boolean;
	 data_in :  in std_logic_vector(data_width-1 downto 0);
	 data_out :  out std_logic_vector(data_width-1 downto 0);
         clk : in std_logic;
         reset: in std_logic
	);
end UnloadFsmNoBlock;

architecture default_arch of UnloadFsmNoBlock is
	signal unload_ack_sig : boolean;
	signal unload_ack_d_sig : boolean;

	signal write_ack_sig: std_logic;

	type FsmState is (Idle, WhatWillItBe, DataValid, ZeroData);
	signal fsm_state : FsmState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch

	process(fsm_state, write_req, data_in,  unload_req, clk, reset)
		variable next_fsm_state_var : FsmState;
		variable unload_ack_d_var: boolean;
		variable write_ack_var : std_logic;

		variable data_out_var: std_logic_vector(data_width-1 downto 0);

	begin
		unload_ack_d_var := false;

		write_ack_var  := '0';
		next_fsm_state_var := fsm_state;

		data_out_var := data_in;

		case fsm_state is 
			-- reset state, nothing seen so far.
			when Idle =>
				if(unload_req) then
					unload_ack_d_var := true;
					next_fsm_state_var := WhatWillItBe;
				end if;
			when ZeroData => 
				-- Acked state, hold until next unload-req
				-- hold 0 data until next unload-req.
				data_out_var := (others => '0');
				if(unload_req) then
					unload_ack_d_var := true;
					next_fsm_state_var := WhatWillItBe;
				end if;
			when DataValid =>
				-- Acked state, hold until next unload-req
				-- write_req is '1' here... 
				if(unload_req) then
					unload_ack_d_var := true;

					-------------------------------
					-- ack it here..
					-------------------------------
					write_ack_var    := '1';
					-------------------------------

					-- what will we see next?
					next_fsm_state_var := WhatWillItBe;
				end if;
			when WhatWillItBe =>
				-- 
				-- Acked state, but data will be determined
				-- in this state.
				--
				if(write_req = '0') then

					-- zero data..
					data_out_var := (others => '0');
					

					if(unload_req) then
						unload_ack_d_var := true;
					else
						-- hold zero data.	
						next_fsm_state_var := ZeroData;
					end if;
				else 
					-- valid data, must hold until next
					-- unload-req.
						

					if(unload_req) then
						unload_ack_d_var := true;

						-------------------------------
						-- ack it here..
						-------------------------------
						write_ack_var    := '1';
						-------------------------------
					else
						next_fsm_state_var := DataValid;
					end if;
				end if;
		end case;

		write_ack_sig <= write_ack_var;
		data_out <= data_out_var;

		if(clk'event and clk='1') then
			if(reset = '1') then
				fsm_state <= Idle;
				unload_ack_d_sig <= false;
			else
				fsm_state <= next_fsm_state_var;
				unload_ack_d_sig <= unload_ack_d_var;
			end if;
		end if;
	end process;

	unload_ack <= unload_ack_d_sig;
	write_ack  <= write_ack_sig;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity UnloadFsm is
  generic (name: string; data_width: integer);
  port ( 
	 write_req: in std_logic;
         write_ack: out std_logic;
         unload_req: in boolean;
         unload_ack: out boolean;
	 data_in :  in std_logic_vector(data_width-1 downto 0);
	 data_out :  out std_logic_vector(data_width-1 downto 0);
         clk : in std_logic;
         reset: in std_logic
	);
end UnloadFsm;

architecture default_arch of UnloadFsm is
	signal unload_ack_sig : boolean;
	signal unload_ack_d_sig : boolean;

	signal write_ack_sig: std_logic;

	type FsmState is (Idle, DataValid, WaitOnData);
	signal fsm_state : FsmState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch

	process(fsm_state, write_req, data_in,  unload_req, clk, reset)
		variable next_fsm_state_var : FsmState;
		variable unload_ack_var: boolean;
		variable unload_ack_d_var: boolean;
		variable write_ack_var : std_logic;

		variable data_out_var: std_logic_vector(data_width-1 downto 0);

	begin
		unload_ack_var := false;
		unload_ack_d_var := false;

		write_ack_var  := '0';
		next_fsm_state_var := fsm_state;

		data_out_var := data_in;

		case fsm_state is 
			-- reset state, nothing seen so far.
			when Idle =>
				if(unload_req) then
					if(write_req = '1') then
						next_fsm_state_var := DataValid;
						unload_ack_d_var := true;
					else
						next_fsm_state_var := WaitOnData;
					end if;
				end if;
			when DataValid =>
				-- write_req = '1' got you here.  Suppress the
				-- write ack until the next unload req.
				if(unload_req) then
					-- pop!
					-- ack the writer, go to wait on data.
					write_ack_var := '1';

					-- we don't know if the next cycle will
					-- have data or not.
					next_fsm_state_var := WaitOnData;
				end if;
			when WaitOnData  =>
				-- This is the "fast" state.
				if (write_req = '1') then
					unload_ack_var := true;

					if(unload_req) then
						write_ack_var := '1';
						-- stay in this state..
					else
						next_fsm_state_var := DataValid;
					end if;
				end if;
		end case;

		unload_ack_sig <= unload_ack_var;
		write_ack_sig <= write_ack_var;
		data_out <= data_out_var;

		if(clk'event and clk='1') then
			if(reset = '1') then
				fsm_state <= Idle;
				unload_ack_d_sig <= false;
			else
				fsm_state <= next_fsm_state_var;
				unload_ack_d_sig <= unload_ack_d_var;
			end if;
		end if;
	end process;

	unload_ack <= unload_ack_sig or unload_ack_d_sig;
	write_ack  <= write_ack_sig;

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity UnloadRegister is
  generic (name: string; 
		data_width : integer ; 
		bypass_flag: boolean := false;  -- if specified, bypasses in->out if possible.
		nonblocking_read_flag : boolean := false);
  port ( write_req: in std_logic;
        write_ack: out std_logic;
        write_data: in std_logic_vector(data_width-1 downto 0);
        unload_req: in boolean;
        unload_ack: out boolean;
        read_data: out std_logic_vector(data_width-1 downto 0);
        clk : in std_logic;
        reset: in std_logic);
end UnloadRegister;

architecture default_arch of UnloadRegister is
	signal unload_ack_sig : boolean;
	signal write_req_nonblockified : std_logic;
	signal write_data_nonblockified: std_logic_vector(data_width-1 downto 0);
	type FsmState is (Idle, Waiting);
	signal fsm_state : FsmState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- default_arch


    noBypass: if not bypass_flag generate 
	-- FSM
  	--   Two states: Idle, Waiting
  	process(clk, reset, fsm_state, unload_req, write_req, write_data)
     		variable nstate: FsmState;
     		variable load_v : boolean;
		variable write_ack_v : std_logic;
		variable data_v : std_logic_vector(data_width-1 downto 0);
        begin
     		nstate :=  fsm_state;
		write_ack_v := '0';
     		load_v := false;
		data_v := write_data;
  		
     		case fsm_state is
         		when Idle => 
               			if(unload_req) then
					write_ack_v := '1';
					if (write_req = '1') then
						load_v := true;
					elsif nonblocking_read_flag then
						load_v := true;
						data_v := (others => '0'); -- non-blocking!
					else
						nstate := Waiting;
					end if;
				end if;
	 		when Waiting =>
				write_ack_v := '1';
				if(write_req = '1') then
					load_v := true;
					nstate := Idle;
				end if;
     		end case;
 
		write_ack <= write_ack_v;
		
     		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= idle;
				unload_ack <= false;
           			read_data <= (others => '0');
			else
				fsm_state <= nstate;
				unload_ack <= load_v;
				if(load_v) then
           				read_data <= data_v;
        			end if;
			end if;
		
     		end if;
  	end process;
   end generate noBypass;

  --
  -- buffer_size = 0 means we want a fast write_data->read_data path
  -- with the UnloadBuffer just doing protocol conversion.
  --
  yesBypassNonBlocking: if bypass_flag and nonblocking_read_flag generate
     bypassBlock: block
        signal bypass_reg_flag: Boolean;
	signal write_data_reg, write_data_prereg: std_logic_vector(data_width-1 downto 0);

        -- delayed and immediate versions of unload-ack
	-- corresponding to the two possible unload scenarios.
	signal unload_ack_sig: boolean;
     begin
    
	-- FSM
  	--   Two states: Idle, Waiting
  	process(clk,fsm_state, unload_req, write_req, write_data)
     		variable nstate: FsmState;
     		variable loadv : boolean;
     		variable write_ackv: std_logic;
     		variable datav: std_logic_vector(data_width-1 downto 0);
        begin
     		nstate :=  fsm_state;
     		write_ackv := '0';

     		loadv := false;
     		datav := (others => '0');
  		
     		case fsm_state is
         		when idle => 
               			if(unload_req) then
					nstate := Waiting;
               			end if;
	 		when Waiting =>
		    		write_ackv := '1';
				loadv   := true;

				-- write-data is 0 unless write-reg='1'.
				if(write_req = '1') then
		    			datav := write_data;
				end if;


				if(not unload_req) then
					nstate := Idle;
				end if;
     		end case;
 
     		write_ack <= write_ackv;
                unload_ack_sig <= loadv;
		write_data_prereg <= datav;
		
     		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= idle;
           			write_data_reg <= (others => '0');
			else
				fsm_state <= nstate;
				if(loadv) then
           				write_data_reg <= datav;
        			end if;
			end if;
     		end if;
  	end process;
        read_data <= write_data_prereg when unload_ack_sig else write_data_reg;
	unload_ack <= unload_ack_sig;
    end block;
  end generate yesBypassNonBlocking;

  yesBypassBlocking: if bypass_flag and (not nonblocking_read_flag) generate
     bypassBlock: block
	type FsmStateBypass is (Idle, Waiting_1, Waiting_2);
        signal bypass_reg_flag: Boolean;
	signal write_data_reg, write_data_prereg: std_logic_vector(data_width-1 downto 0);

        -- delayed and immediate versions of unload-ack
	-- corresponding to the two possible unload scenarios.
	signal unload_ack_sig: boolean;
	signal fsm_state_bypass : FsmStateBypass;
     begin
    
	-- FSM
  	--   Three states: Idle, Waiting_1, Waiting_2.. Not clear
	--     why we need Waiting_1 and Waiting_2?  I thought I
	--     had a reason for this.. Let the synthesis tool 
	--     optimize this one.
	--
	-- creates a forward path from write_req to unload_ack..
	-- 
  	process(clk,fsm_state_bypass, unload_req, write_req, write_data)
     		variable nstate: FsmStateBypass;
     		variable loadv : boolean;
     		variable write_ackv: std_logic;
     		variable datav: std_logic_vector(data_width-1 downto 0);
        begin
     		nstate :=  fsm_state_bypass;
     		write_ackv := '0';

     		loadv := false;
		datav := write_data;
  		
     		case fsm_state_bypass is
         		when idle => 
               			if(unload_req) then
					nstate := Waiting_1;
               			end if;
	 		when Waiting_1 =>
				-- unload-req observed in previous cycle, wait for write-req.
		    		write_ackv := '1';

				if (write_req = '1') then
					loadv   := true;
					if(not unload_req) then
						-- no unload-req? go to idle..
						-- else stay here..
						nstate := Idle;
					end if;
				else
					nstate := Waiting_2;
				end if;
			when Waiting_2 =>
				-- unload req observed.. but not immediately
				-- previous cycle.  Idle and Waiting_2 are 
				-- distinguished by the fact that when we
				-- are in Waiting_2, we have a pending unload.
		    		write_ackv := '1';
				if(write_req = '1') then
					loadv := true;
					if(unload_req) then
						nstate := Waiting_1;
					else
						nstate := Idle;
					end if;
				end if;
     		end case;
 
     		write_ack <= write_ackv;
                unload_ack_sig <= loadv;
		write_data_prereg <= datav;
		
     		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state_bypass <= Idle;
           			write_data_reg <= (others => '0');
			else
				fsm_state_bypass <= nstate;
				if(loadv) then
           				write_data_reg <= datav;
        			end if;
			end if;
     		end if;
  	end process;
	-- note bypass..
        read_data <= write_data_prereg when unload_ack_sig else write_data_reg;
	unload_ack <= unload_ack_sig;
    end block;
  end generate yesBypassBlocking;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- TODO: add bypass generic to create a flow-through
--       trivial operator (to save clock-cycles!)
--
-- The unshared operator uses a split protocol.
--    reqL/ackL  for sampling the inputs
--    reqR/ackR  for updating the outputs.
-- The two pairs should be used independently,
-- that is, there should be NO DEPENDENCY between
-- ackL and reqR!
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.OperatorPackage.all;
use ahir.BaseComponents.all;
use ahir.FloatOperatorPackage.all;

entity UnsharedOperatorWithBuffering is
  generic
    (
      name   : string;
      operator_id   : string;          -- operator id
      input1_is_int : Boolean := true; -- false means float
      input1_characteristic_width : integer := 0; -- characteristic width if input1 is float
      input1_mantissa_width       : integer := 0; -- mantissa width if input1 is float
      iwidth_1      : integer;    -- width of input1
      input2_is_int : Boolean := true; -- false means float
      input2_characteristic_width : integer := 0; -- characteristic width if input2 is float
      input2_mantissa_width       : integer := 0; -- mantissa width if input2 is float
      iwidth_2      : integer;    -- width of input2
      num_inputs    : integer := 2;    -- can be 1 or 2.
      output_is_int : Boolean := true;  -- false means that the output is a float
      output_characteristic_width : integer := 0;
      output_mantissa_width       : integer := 0;
      owidth        : integer;          -- width of output.
      constant_operand : std_logic_vector; -- constant operand.. (it is always the second operand)
      constant_width : integer;
      buffering      : integer;
      use_constant  : boolean := false;
      flow_through  : boolean := false;
      full_rate: boolean 
      );
  port (
    -- req -> ack follow pulse protocol
    reqL:  in Boolean;
    ackL : out Boolean;
    reqR : in Boolean;
    ackR:  out Boolean;
    -- operands.
    dataL      : in  std_logic_vector(iwidth_1 + iwidth_2 - 1 downto 0);
    dataR      : out std_logic_vector(owidth-1 downto 0);
    clk, reset : in  std_logic);
end UnsharedOperatorWithBuffering;


architecture Vanilla of UnsharedOperatorWithBuffering is
  signal   result: std_logic_vector(owidth-1 downto 0);
  constant iwidth : integer := iwidth_1  + iwidth_2;
  
  -- joined req, and joint ack.
  signal fReq,fAck: boolean;
 

begin  -- Behave

  assert((num_inputs = 1) or (num_inputs = 2)) report "either 1 or 2 inputs" severity failure;
  -----------------------------------------------------------------------------
  -- combinational block..
  -----------------------------------------------------------------------------
  comb_block: GenericCombinationalOperator
    generic map (
      name => name & "-comb_block",
      operator_id                 => operator_id,
      input1_is_int               => input1_is_int,
      input1_characteristic_width => input1_characteristic_width,
      input1_mantissa_width       => input1_mantissa_width,
      iwidth_1                    => iwidth_1,
      input2_is_int               => input2_is_int,
      input2_characteristic_width => input2_characteristic_width,
      input2_mantissa_width       => input2_mantissa_width,
      iwidth_2                    => iwidth_2,
      num_inputs                  => num_inputs,
      output_is_int               => output_is_int,
      output_characteristic_width => output_characteristic_width,
      output_mantissa_width       => output_mantissa_width,
      owidth                      => owidth,
      constant_operand            => constant_operand,
      constant_width              => constant_width,
      use_constant                => use_constant)
    port map (data_in => dataL, result  => result);


  noFlowThrough: if not flow_through generate
    -----------------------------------------------------------------------------
    -- output interlock buffer
    -----------------------------------------------------------------------------
    ilb: InterlockBuffer 

	  generic map(name => name & "-ilb",
			  buffer_size => buffering,
			  in_data_width => owidth,
			  out_data_width => owidth) 

	  port map(write_req => reqL, write_ack => ackL, write_data => result,
			  read_req => reqR, read_ack => ackR, read_data => dataR,
				  clk => clk, reset => reset);
  end generate noFlowThrough;

  flowThrough: if flow_through generate
		-- in the flow-through case, the operator looks just like
		-- a combinational circuit.  
                -- NOTE that there is no bypass register for the data.
                -- Control sequencing must be handled entirely by the
		-- control-path which uses this operator.

		ackL <= reqL;
		ackR <= reqR;
		dataR <= result;

  end generate flowThrough;

end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.Types.all;
use ahir.Utilities.all;
use ahir.Subprograms.all;

entity BypassRegister  is
	generic (data_width: integer; bypass: boolean);
	port (clk, reset: in std_logic; enable: in boolean; 
			din: in std_logic_vector(data_width-1 downto 0);
			q: out std_logic_vector(data_width-1 downto 0));
end entity;

architecture Behaveee of  BypassRegister is
   signal din_reg: std_logic_vector(data_width-1 downto 0);
begin
	process(clk,reset, enable)
	begin
		if(clk'event and clk = '1') then
			if reset = '1' then
				din_reg <= (others => '0');
			elsif enable then
				din_reg <= din;
			end if;
		end if;
	end process;
   ifByp: if bypass generate
	q <= din when enable else din_reg;
   end generate ifByp;
   ifNoByp: if not bypass generate
	q <= din_reg;
   end generate ifNoByp;
end Behaveee;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Components.all;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.GlobalConstants.all;

--  input port specialized for P2P ports.
entity InputPort_P2P is
  generic (name : string;
	   data_width: integer;
	   queue_depth: integer;
	   bypass_flag: boolean := false;
	   barrier_flag: boolean := false;
	   nonblocking_read_flag: boolean);
  port (
    -- pulse interface with the data-path
    sample_req        : in  Boolean; -- sacrificial.
    sample_ack        : out Boolean; -- sacrificial.
    update_req        : in  Boolean;
    update_ack        : out Boolean;
    data              : out std_logic_vector(data_width-1 downto 0);
    -- ready/ready interface with outside world
    oreq       : out std_logic;
    oack       : in  std_logic;
    odata      : in  std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
end entity;


architecture Base of InputPort_P2P is
  signal noblock_update_req, noblock_update_ack: boolean;
  signal noblock_data : std_logic_vector(data_width-1 downto 0);
  type SampleFsmState is (IDLE, WAITING);
  signal fsm_state: SampleFsmState;
  signal has_data: std_logic;

  -- Don't f-around with this.
  constant use_unload_register :boolean :=  (not global_use_optimized_unload_buffer) or bypass_flag;

begin

    noBarrier: if (not barrier_flag) or nonblocking_read_flag generate
	sample_ack <= sample_req;
    end generate noBarrier; 

    withBarrier: if (barrier_flag and (not nonblocking_read_flag)) generate
     -- sample ack when there is something at the 
     -- input of the port.  This is useful in 
     -- setting up barriers.
       process(clk, reset, fsm_state, sample_req, oack)
       	variable next_fsm_state: SampleFsmState;
       begin
	next_fsm_state := fsm_state;
	sample_ack <= false;
	case fsm_state is
		when IDLE => 
			if ((oack = '1') or (has_data = '1')) then
				sample_ack <= sample_req;
			elsif sample_req then
				next_fsm_state := WAITING;
			end if;
		when WAITING => 
			if (has_data = '1') or (oack = '1') then
				sample_ack <= true;
				next_fsm_state := IDLE;
			end if;
	end case;
	if(clk'event and clk = '1') then
		if(reset = '1') then
			fsm_state <= IDLE;
		else
			fsm_state <= next_fsm_state;
		end if;
	end if;
       end process;
     end generate withBarrier;
	
     ub: UnloadBuffer
	generic map (name => name & "-ub", 
				data_width => data_width,
				   buffer_size => queue_depth, 
					bypass_flag => bypass_flag,  
						use_unload_register => use_unload_register,
							nonblocking_read_flag => nonblocking_read_flag)
	port map (write_req => oack, write_ack => oreq, 
					write_data => odata,
				unload_req => update_req,
				unload_ack => update_ack,
				has_data => has_data,
				read_data =>  data, clk => clk, reset => reset);
end Base;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity PipeJoin is
  generic (name : string; data_width_0, data_width_1: integer);
  port (
    write_req_0   : in std_logic;
    write_ack_0   : out std_logic;
    write_data_0   : in std_logic_vector(data_width_0-1 downto 0);
    write_req_1   : in std_logic;
    write_ack_1   : out std_logic;
    write_data_1   : in std_logic_vector(data_width_1-1 downto 0);
    read_req      : in  std_logic;
    read_ack       : out std_logic;
    read_data     : out std_logic_vector((data_width_1 + data_width_0)-1 downto 0);
    clk, reset : in  std_logic);
end PipeJoin;

architecture default_arch of PipeJoin is
begin  -- default_arch
   assert false report "NOT IMPLEMENTED" severity ERROR;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity PipeMerge is
  generic (name : string; data_width_0, data_width_1: integer);
  port (
    write_req_0   : in std_logic;
    write_ack_0   : out std_logic;
    write_data_0   : in std_logic_vector(data_width_0-1 downto 0);
    write_req_1   : in std_logic;
    write_ack_1   : out std_logic;
    write_data_1   : in std_logic_vector(data_width_1-1 downto 0);
    read_req      : in  std_logic;
    read_ack       : out std_logic;
    read_data     : out std_logic_vector((data_width_1 + data_width_0)-1 downto 0);
    clk, reset : in  std_logic);
end PipeMerge;

architecture default_arch of PipeMerge is
begin  -- default_arch
   assert false report "NOT IMPLEMENTED" severity ERROR;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity PipeMux is
  generic (name : string; data_width: integer);
  port (
    write_req_0   : in std_logic;
    write_ack_0   : out std_logic;
    write_data_0   : in std_logic_vector(data_width-1 downto 0);
    write_req_1   : in std_logic;
    write_ack_1   : out std_logic;
    write_data_1   : in std_logic_vector(data_width-1 downto 0);
    read_req      : in  std_logic;
    read_ack       : out std_logic;
    read_data     : out std_logic_vector(data_width-1 downto 0);
    clk, reset : in  std_logic);
end PipeMux;

architecture default_arch of PipeMux is

   signal priority_flag: std_logic;
  
begin  -- default_arch
   assert false report "NOT IMPLEMENTED" severity ERROR;
end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;

entity PipeSizeMonitor is
  generic (name : string; depth: integer);
  port (
    write_req   : in  std_logic;
    write_ack   : in  std_logic;
    read_req    : in  std_logic;
    read_ack    : in  std_logic;
    has_data    : out Boolean;
    clk, reset  : in  std_logic);
end PipeSizeMonitor;

architecture default_arch of PipeSizeMonitor is
  signal number_of_elements_in_pipe: unsigned ((Ceil_Log2(depth+2))-1 downto 0); 
begin  -- default_arch
		-- count number of elements in pipe.
	process(clk, reset)
  	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				number_of_elements_in_pipe <= (others => '0');
			else
				if((read_req = '1') and (read_ack = '1')) then
					if(not ((write_req = '1') and (write_ack = '1'))) then
				          number_of_elements_in_pipe <= (number_of_elements_in_pipe -1);
					end if;
				elsif((write_req = '1') and (write_ack = '1')) then
					number_of_elements_in_pipe <= (number_of_elements_in_pipe + 1);
				end if;
			end if;
		end if;
  	end process;
	
  	has_data <= (number_of_elements_in_pipe > 0);

end default_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.Utilities.all;

--
-- higher in->out latency, but distributed in space (think ASIC, ASIC).
-- often good enough.
--
entity ShiftRegisterQueue is
  generic(name : string; queue_depth: integer := 1; data_width: integer := 32);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(data_width-1 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(data_width-1 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity ShiftRegisterQueue;

architecture behave of ShiftRegisterQueue is

  type QueueArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);
  constant n_stages : integer := (queue_depth + 1)/2;
  signal intermediate_data: QueueArray(0 to n_stages);
  signal intermediate_lr_req: std_logic_vector(0 to n_stages);
  signal intermediate_lr_ack: std_logic_vector(0 to n_stages);

begin  -- SimModel

     intermediate_data(0) <= data_in;
     intermediate_lr_req(0) <= push_req;
     push_ack <= intermediate_lr_ack(0);

     stageGen: for I in 0 to n_stages-1 generate
	qinst: QueueBase 
		generic map (name => name & "-stageGen-qinst-" & Convert_To_String(I),
				queue_depth => 2, data_width => data_width)
		port map ( reset => reset, clk => clk, 
			data_in => intermediate_data(I),
			push_req => intermediate_lr_req(I),
			push_ack => intermediate_lr_ack(I),
			pop_req  => intermediate_lr_ack(I+1), -- cross-over
			pop_ack => intermediate_lr_req(I+1), -- cross-over
			data_out => intermediate_data(I+1));
     end generate stageGen;

     data_out <= intermediate_data(n_stages);
     intermediate_lr_ack(n_stages) <= pop_req;
     pop_ack <= intermediate_lr_req(n_stages);

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.Utilities.all;
use ahir.GlobalConstants.all;

--
-- higher in->out latency, but distributed in space (think ASIC, ASIC).
-- often good enough.
--
entity ShiftRegisterSingleBitQueue is
  generic(name : string; queue_depth: integer; number_of_stages: integer; bypass_flag: boolean := false);
  port(clk: in std_logic;
       reset: in std_logic;
       data_in: in std_logic_vector(0 downto 0);
       push_req: in std_logic;
       push_ack: out std_logic;
       data_out: out std_logic_vector(0 downto 0);
       pop_ack : out std_logic;
       pop_req: in std_logic);
end entity ShiftRegisterSingleBitQueue;

architecture behave of ShiftRegisterSingleBitQueue is

  constant stage_depth : integer := Ceil(queue_depth, number_of_stages);

  signal intermediate_data:   std_logic_vector(0 to number_of_stages);
  signal intermediate_lr_req: std_logic_vector(0 to number_of_stages);
  signal intermediate_lr_ack: std_logic_vector(0 to number_of_stages);

begin  -- SimModel

	assert(number_of_stages > 0) report "In " & name & " number of stages must be > 0 " severity failure;

     intermediate_data(0) <= data_in(0);
     intermediate_lr_req(0) <= push_req;
     push_ack <= intermediate_lr_ack(0);

     stageGen: for I in 0 to number_of_stages-1 generate
	qinst: SingleBitQueueBase 
		generic map (name => name & "-stageGen-qinst-" & Convert_To_String(I),
				queue_depth => stage_depth, bypass_flag => bypass_flag)
		port map ( reset => reset, clk => clk, 
				data_in => intermediate_data(I to I),
				push_req => intermediate_lr_req(I),
				push_ack => intermediate_lr_ack(I),
				pop_req  => intermediate_lr_ack(I+1), -- cross-over
				pop_ack => intermediate_lr_req(I+1), -- cross-over
				data_out => intermediate_data((I+1) to (I+1)));
     end generate stageGen;

     data_out(0) <= intermediate_data(number_of_stages);
     intermediate_lr_ack(number_of_stages) <= pop_req;
     pop_ack <= intermediate_lr_req(number_of_stages);

end behave;
library ieee;
use ieee.std_logic_1164.all;

entity SingleCycleStartFinFsm is
	port (clk, reset, start_req, fin_req : in std_logic;
		enable, start_ack, fin_ack: out std_logic) ;
end entity SingleCycleStartFinFsm;

architecture BehaveProcess of SingleCycleStartFinFsm is
       signal fin_ack_sig: std_logic;
begin
	fin_ack <= fin_ack_sig;

	process(clk,reset, fin_req, start_req, fin_ack_sig)
		variable next_fin_ack_sig: std_logic;
		variable enable_var : std_logic;
	begin
		next_fin_ack_sig := fin_ack_sig;
		enable_var := '0';

		case fin_ack_sig is
			when '0' =>
				if(start_req = '1') then
					enable_var := '1';
					next_fin_ack_sig := '1';
				end if;
			when '1' =>
				if((fin_req = '1') and (start_req  = '1')) then
					enable_var := '1';
				elsif (fin_req = '1') then
					next_fin_ack_sig := '0';
				end if;
			when others => 
				null;
		end case;

		enable <= enable_var;
                start_ack <= enable_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fin_ack_sig <= '0';
			else
				fin_ack_sig <= next_fin_ack_sig;
			end if;
		end if;
	end process;
end BehaveProcess; 
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

entity LevelRepeater is
    generic(name: string; g_data_width: integer := 32; g_depth : integer := 1);
    port(clk: in std_logic;
       		reset: in std_logic;
		enable: in std_logic;
       		data_in: in std_logic_vector(g_data_width-1 downto 0);
       		valid_in: in std_logic;
       		data_out: out std_logic_vector(g_data_width-1 downto 0);
       		valid_out : out std_logic;
       		stall: in std_logic);
end entity LevelRepeater;

architecture behave of LevelRepeater is
	signal ivalids: std_logic_vector(0 to g_depth);
	type DwordArray is array (natural range <>) of std_logic_vector (g_data_width-1 downto 0);
	signal data_regs: DwordArray(0 to g_depth);
begin  -- SimModel

        assert (g_depth > 0) report "LevelRepeater:" & name & " depth must be > 0" severity error;

	ivalids(0) <= valid_in;
	-- if enable is low, we stuff the data-in else we stuff in the
	-- last data seen..  (repeat it..)
 	nontriv: if (g_depth > 0) generate
        	data_regs(0) <= data_in when (enable = '1') else data_regs(1);
	end generate nontriv;
 	triv: if (g_depth = 0) generate
        	data_regs(0) <= data_in;
	end generate triv;

	valid_out  <= ivalids(g_depth);
        data_out   <= data_regs(g_depth);

        genSR: for I in 1 to g_depth generate 
	  process(clk, reset)
	  begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				ivalids(I) <= '0';
			elsif (stall = '0') then
				ivalids(I) <= ivalids(I-1);
				data_regs(I)  <= data_regs(I-1);
			end if;
		end if;
   	   end process;
        end generate genSR;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

-- Forget the fancy name. This is a shift register in which
-- the decision to shift at each stage is determined by a 
-- stall-vector.  The enable re-inserts that last inserted value into
-- the shift register.
entity SquashLevelRepeater is
    generic(name: string; g_data_width: integer := 32; g_depth : integer := 1);
    port(clk: in std_logic;
       		reset: in std_logic;
		enable: in std_logic;
       		data_in: in std_logic_vector(g_data_width-1 downto 0);
       		data_out: out std_logic_vector(g_data_width-1 downto 0);
       		stall_vector: in std_logic_vector(1 to g_depth));
end entity SquashLevelRepeater;

architecture behave of SquashLevelRepeater is
	type DwordArray is array (natural range <>) of std_logic_vector (g_data_width-1 downto 0);
	signal data_regs: DwordArray(0 to g_depth);
begin  -- SimModel

        assert (g_depth > 0) report "SquashLevelRepeater:" & name & " depth must be > 0" severity error;

	-- if enable is high, we stuff the data-in else we stuff in the
	-- last data seen..  (ie, hold it.)
 	nontriv: if (g_depth > 0) generate
        	data_regs(0) <= data_in when (enable = '1') else data_regs(1);
	end generate nontriv;
 	triv: if (g_depth = 0) generate
        	data_regs(0) <= data_in;
	end generate triv;

        data_out   <= data_regs(g_depth);

        genSR: for I in 1 to g_depth generate 
	  process(clk)
	  begin
		if(clk'event and clk = '1') then
			if (stall_vector(I) = '0') then
				data_regs(I)  <= data_regs(I-1);
			end if;
		end if;
   	   end process;
        end generate genSR;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

-- a stall protocol to pulse translator used at the
-- output end of a data-path operator in order
-- to interface to the control path.
-- Madhav Desai.
entity Stall_To_Pulse_Translate_Entity is
  generic (name : string);
  port(
	stall_out : out std_logic;
        rR : in  boolean;
        valid_in : in std_logic;
        aR : out boolean;
        clk : in std_logic;
        reset : in std_logic);
end entity;

architecture Behave of Stall_To_Pulse_Translate_Entity is
  type S2PState is (Idle, WaitForValid, HoldValue);
  signal s2p_state : S2PState;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin  -- Behave

  process(clk, reset, valid_in, rR, s2p_state)
    variable nstate : S2PState;
    variable stall_out_var: std_logic;
  begin
    nstate := s2p_state;
    stall_out_var := '1';
    aR <= false;

    case s2p_state is
        when Idle =>
	  stall_out_var :=  valid_in; -- if valid is observed, start stalling.
          if(rR) then
              nstate := WaitForValid;
          end if;
        when WaitForValid => -- rR has been observed, we are waiting for valid-in.
          stall_out_var := valid_in;  -- stall if valid is observed.
          if(valid_in = '1') then
            aR <= true;
	    if(not rR) then
	      nstate := HoldValue;  -- hold value until rR.
	    else
	      stall_out_var := '0'; -- rR seen, no need to hold, move the pipeline forward.
	    end if;
          end if; 
        when HoldValue =>  -- hold the value until the next rR;
          stall_out_var := '1';  -- keep stalling until rR...
	  if (rR) then
	     nstate := WaitForValid;
             stall_out_var := '0'; -- quit stalling, no need to hold value..
	  end if;
    end case;

    stall_out <= stall_out_var;

    if(clk'event and clk = '1') then
	if reset = '1' then
		s2p_state <= Idle;
	else
      		s2p_state <= nstate;
	end if;
    end if;
  end process;
end Behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

--
-- stall_in is used to stall the stages in a shift-register pipeline.
-- A stage is stalled only if its successor is non-empty and has stalled.
--
entity ValidPropagator is
    generic(name: string; g_depth : integer := 1);
    port(clk: in std_logic;
       		reset: in std_logic;
       		stall_in: in std_logic;
       		valid_in: in std_logic;
       		valid_out : out std_logic;
       		stall_vector: out std_logic_vector(1 to  g_depth));
end entity ValidPropagator;

architecture behave of ValidPropagator is
	-- output of th kth stage is valid... 0 is the
	-- input.
	signal ivalids: std_logic_vector(0 to g_depth);

	-- kth stage has stalled.
	signal stalls:  std_logic_vector(1 to (g_depth+1));
begin  -- SimModel

        assert (g_depth > 0) report "ValidPropagator:" & name & " depth must be > 0" severity error;

	ivalids(0) <= valid_in;
	valid_out  <= ivalids(g_depth);

	stalls(g_depth+1) <=  stall_in;
	stall_vector <= stalls(1 to g_depth);

        genSR: for I in 1 to g_depth generate 
	  stalls(I) <= (ivalids(I) and stalls(I+1));

	  process(clk, reset)
	  begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				ivalids(I) <= '0';
			elsif (stalls(I) = '0') then
				ivalids(I) <= ivalids(I-1);
			end if;
		end if;
   	   end process;
        end generate genSR;

end behave;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;


entity fpadd32 is -- 
    generic (name: string := "fpadd32"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpadd32;

architecture Struct of fpadd32 is
begin

   adder: GenericFloatingPointAdderSubtractor
		generic map(name => name & "-adder",
				tag_width => tag_length,
				exponent_width => 8,
				fraction_width => 23,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true,
				use_as_subtractor => false)
		port map(INA => L, INB => R,
				OUTADD => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				addi_rdy => start_ack, addo_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;


entity fpadd64 is -- 
    generic (name: string:= "fpadd64"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpadd64;

architecture Struct of fpadd64 is
begin

   adder: GenericFloatingPointAdderSubtractor
		generic map(name => name & "-adder", tag_width => tag_length,
				exponent_width => 11,
				fraction_width => 52,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true,
				use_as_subtractor => false)
		port map(INA => L, INB => R,
				OUTADD => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				addi_rdy => start_ack, addo_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;


entity fpmul32 is -- 
    generic (name: string:= "fpmul32"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpmul32;

architecture Struct of fpmul32 is
begin

   mul: GenericFloatingPointMultiplier
		generic map(name => name & "-mul", tag_width => tag_length,
				exponent_width => 8,
				fraction_width => 23,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true)
		port map(INA => L, INB => R,
				OUTMUL => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				muli_rdy => start_ack, mulo_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;


entity fpmul64 is -- 
    generic (name: string:= "fpmul64"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpmul64;

architecture Struct of fpmul64 is
begin

   mul: GenericFloatingPointMultiplier
		generic map(name => name & "-mul", tag_width => tag_length,
				exponent_width => 11,
				fraction_width => 52,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true)
		port map(INA => L, INB => R,
				OUTMUL => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				muli_rdy => start_ack, mulo_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;


entity fpsub32 is -- 
    generic (name: string := "fpsub32"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpsub32;

architecture Struct of fpsub32 is
begin

   sub: GenericFloatingPointAdderSubtractor
		generic map(name => name & "-sub", tag_width => tag_length,
				exponent_width => 8,
				fraction_width => 23,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true,
				use_as_subtractor => true)
		port map(INA => L, INB => R,
				OUTADD => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				addi_rdy => start_ack, addo_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;


entity fpsub64 is -- 
    generic (name: string := "fpsub64"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpsub64;

architecture Struct of fpsub64 is
begin

   sub: GenericFloatingPointAdderSubtractor
		generic map(name => name & "-sub", tag_width => tag_length,
				exponent_width => 11,
				fraction_width => 52,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true,
				use_as_subtractor => true)
		port map(INA => L, INB => R,
				OUTADD => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				addi_rdy => start_ack, addo_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;


entity fpu32 is -- 
    generic (name: string := "fpu32"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      OP_ID : in std_logic_vector(7 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpu32;

architecture Struct of fpu32 is
      signal OUTADD, OUTMUL, addsub_L, addsub_R : std_logic_vector(31 downto 0);
      signal req_to_omux, ack_from_omux: std_logic_vector(1 downto 0);

      signal data_to_omux: std_logic_vector((2*(32+tag_length))-1 downto 0);
      signal data_from_omux: std_logic_vector((32+tag_length)-1 downto 0);
      signal reqi_omux: std_logic_vector(1 downto 0);
      signal acki_omux: std_logic_vector(1 downto 0);
       
      signal mul_tag_out, addsub_tag_out: std_logic_vector(tag_length-1 downto 0);

      signal muli_req, addsubi_req: std_logic;
      signal muli_ack, addsubi_ack: std_logic;
      signal mulo_req, addsubo_req: std_logic;
      signal mulo_ack, addsubo_ack: std_logic;


      
begin

   muli_req <= start_req when (OP_ID = "00000010") else '0';
   addsubi_req <= start_req when ((OP_ID="00000001") or (OP_ID = "00000000")) else '0';
   start_ack <= muli_ack when (OP_ID = "00000010") else addsubi_ack when 
			((OP_ID="00000001") or (OP_ID = "00000000")) else '0';

   addsub_L <= L;
   process(R, OP_ID)
	variable X: std_logic_vector(31 downto 0);
   begin
	X(30 downto 0) := R(30 downto 0);
	if(OP_ID = "00000001") then
		X(31) := not R(31);
	else
		X(31) := R(31);
	end if;
	addsub_R <= X;
   end process;

   addsub: GenericFloatingPointAdderSubtractor
		generic map(name => name & "-addsub", tag_width => tag_length,
				exponent_width => 8,
				fraction_width => 23,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true,
				use_as_subtractor => false)
		port map(INA => addsub_L, INB => addsub_R,
				OUTADD => OUTADD,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => addsub_tag_out,
				env_rdy => addsubi_req, accept_rdy => addsubo_req,
				addi_rdy => addsubi_ack, addo_rdy => addsubo_ack);

   mul: GenericFloatingPointMultiplier
		generic map(name => name & "-mul", tag_width => tag_length,
				exponent_width => 8,
				fraction_width => 23,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true)
		port map(INA => L, INB => R,
				OUTMUL => OUTMUL,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => mul_tag_out,
				env_rdy => muli_req, accept_rdy => mulo_req,
				muli_rdy => muli_ack, mulo_rdy => mulo_ack);

   data_to_omux <= OUTADD & addsub_tag_out & OUTMUL & mul_tag_out;
   reqi_omux(1) <= addsubo_ack;
   reqi_omux(0) <= mulo_ack;
   addsubo_req <= acki_omux(1);
   mulo_req <= acki_omux(0);


   omux:  OutputPortLevel generic map(name => name & "-omux", num_reqs => 2,
					data_width => data_from_omux'length,
					no_arbitration => false)
			port map(req => reqi_omux,
				ack => acki_omux,
				data => data_to_omux,
				oreq => fin_ack,
				oack => fin_req,
				odata => data_from_omux,
				clk => clk,
				reset => reset);

   ret_val_x_x <= data_from_omux(31+tag_length downto tag_length);
   tag_out <= data_from_omux(tag_length-1 downto 0);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.float_pkg.all;
use aHiR_ieee_proposed.math_utility_pkg.all;


entity fpu64 is -- 
    generic (name: string := "fpu64"; tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(63 downto 0);
      R : in  std_logic_vector(63 downto 0);
      OP_ID : in std_logic_vector(7 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity fpu64;

architecture Struct of fpu64 is
      signal OUTADD, OUTMUL, addsub_L, addsub_R : std_logic_vector(63 downto 0);
      signal req_to_omux, ack_from_omux: std_logic_vector(1 downto 0);

      signal data_to_omux: std_logic_vector((2*(64+tag_length))-1 downto 0);
      signal data_from_omux: std_logic_vector((64+tag_length)-1 downto 0);
      signal reqi_omux: std_logic_vector(1 downto 0);
      signal acki_omux: std_logic_vector(1 downto 0);
       
      signal mul_tag_out, addsub_tag_out: std_logic_vector(tag_length-1 downto 0);

      signal muli_req, addsubi_req: std_logic;
      signal muli_ack, addsubi_ack: std_logic;
      signal mulo_req, addsubo_req: std_logic;
      signal mulo_ack, addsubo_ack: std_logic;


      
begin

   muli_req <= start_req when (OP_ID = "00000010") else '0';
   addsubi_req <= start_req when ((OP_ID="00000001") or (OP_ID = "00000000")) else '0';
   start_ack <= muli_ack when (OP_ID = "00000010") else addsubi_ack when 
			((OP_ID="00000001") or (OP_ID = "00000000")) else '0';

   addsub_L <= L;
   process(R, OP_ID)
	variable X: std_logic_vector(63 downto 0);
   begin
	X := R;
	if(OP_ID = "00000001") then
		X(63) := not R(63);
	end if;
	addsub_R <= X;
   end process;

   addsub: GenericFloatingPointAdderSubtractor
		generic map(name => name & "-addsub", tag_width => tag_length,
				exponent_width => 11,
				fraction_width => 52,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true,
				use_as_subtractor => false)
		port map(INA => addsub_L, INB => addsub_R,
				OUTADD => OUTADD,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => addsub_tag_out,
				env_rdy => addsubi_req, accept_rdy => addsubo_req,
				addi_rdy => addsubi_ack, addo_rdy => addsubo_ack);

   mul: GenericFloatingPointMultiplier
		generic map(name => name & "-mul", tag_width => tag_length,
				exponent_width => 11,
				fraction_width => 52,
                   		round_style => round_nearest,
                   		addguard => 3,
                   		check_error => true,
                   		denormalize => true)
		port map(INA => L, INB => R,
				OUTMUL => OUTMUL,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => mul_tag_out,
				env_rdy => muli_req, accept_rdy => mulo_req,
				muli_rdy => muli_ack, mulo_rdy => mulo_ack);

   data_to_omux <= OUTADD & addsub_tag_out & OUTMUL & mul_tag_out;
   reqi_omux(1) <= addsubo_ack;
   reqi_omux(0) <= mulo_ack;
   addsubo_req <= acki_omux(1);
   mulo_req <= acki_omux(0);


   omux:  OutputPortLevel generic map(name => name & "-omux", num_reqs => 2,
					data_width => data_from_omux'length,
					no_arbitration => false)
			port map(req => reqi_omux,
				ack => acki_omux,
				data => data_to_omux,
				oreq => fin_ack,
				oack => fin_req,
				odata => data_from_omux,
				clk => clk,
				reset => reset);

   ret_val_x_x <= data_from_omux(63+tag_length downto tag_length);
   tag_out <= data_from_omux(tag_length-1 downto 0);
			
end Struct;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity ram_1024x32_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    enable : in  std_logic_vector(0 downto 0);
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(9 downto 0);
    din : in  std_logic_vector(31 downto 0);
    dout : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity ram_1024x32_Operator;
architecture ram_1024x32_Operator_arch of ram_1024x32_Operator is -- 
	signal datain, dataout: std_logic_vector(31 downto 0);
	signal writebar: std_logic;
	signal addrin: std_logic_vector(9 downto 0);
	signal enable_base, enable_bb: std_logic;
	signal start_req, start_ack: std_logic;
	signal ureg_write_req, ureg_write_ack: std_logic;
begin --  
   p2l: Sample_Pulse_To_Level_Translate_Entity
                generic map(name => "ram_1024x32_Operator-p2l")
                port map (rL => sample_req, rR => start_req,
                                aL => sample_ack, aR => start_ack,
                                        clk => clk, reset => reset);

  -- 0 is write-port
  datain <= din;
  addrin <= addr;
  enable_bb <= enable_base and enable(0);
  writebar <= read_write_bar(0);

  bbsp: base_bank
		generic map ("ram_1024x32_base_bank",
					g_addr_width => 10, g_data_width => 32)
		port map (
			clk => clk, reset => reset,
			datain => datain,
			dataout => dataout,
         		addrin => addrin,
         		enable => enable_bb,
         		writebar  => writebar 
		);


   sfsm: SingleCycleStartFinFsm 
			port map (clk => clk, reset => reset,
					-- input
					start_req => start_req, 
					-- output
					start_ack => start_ack,
					-- input
					fin_req => ureg_write_ack, 
					-- output
					fin_ack => ureg_write_req,
					-- same as start-ack
					enable => enable_base);

   ureg: UnloadRegister 
		generic map (name => "ram1024x32:ureg",
				data_width => 32,
				  bypass_flag => true, nonblocking_read_flag => false)
		port map (write_data => dataout,
				write_req => ureg_write_req,
					write_ack => ureg_write_ack,
					    read_data => dout,
						unload_req => update_req,
						   unload_ack => update_ack,
							clk => clk,
							  reset => reset);


end ram_1024x32_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.mem_component_pack.all;

entity dpram_1w_1r_1024x32_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    read_enable : in  std_logic_vector(0 downto 0);
    write_enable : in  std_logic_vector(0 downto 0);
    read_addr : in  std_logic_vector(9 downto 0);
    write_addr : in  std_logic_vector(9 downto 0);
    write_data : in  std_logic_vector(31 downto 0);
    read_data : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity dpram_1w_1r_1024x32_Operator;
architecture dpram_1w_1r_1024x32_Operator_arch of dpram_1w_1r_1024x32_Operator is -- 
	signal datain_0, datain_1, dataout_0, dataout_1, dataout_1_reg, data_to_ulreg: std_logic_vector(31 downto 0);
	signal enable_0, enable_1, enable_1_reg, writebar_0, writebar_1: std_logic;
	signal addrin_0, addrin_1: std_logic_vector(9 downto 0);
	signal enable_base: std_logic;
	signal start_req, start_ack: std_logic;
	signal ureg_write_req, ureg_write_ack: std_logic;
begin 

   p2l: Sample_Pulse_To_Level_Translate_Entity
                generic map(name => "dpram_1w_1r_1024x32_Operator-p2l")
                port map (rL => sample_req, rR => start_req,
                                aL => sample_ack, aR => start_ack,
                                        clk => clk, reset => reset);

  -- 0 is write-port
  datain_0 <= write_data;
  addrin_0 <= write_addr;
  enable_0 <= enable_base and write_enable(0);
  writebar_0 <= '0';

  datain_1 <= (others => '0');
  addrin_1  <= read_addr;
  enable_1 <= enable_base and read_enable(0);
  writebar_1 <= '1';

  -- stabilize the outputs of the dpram.
  process(clk, reset)
  begin
	if(clk'event and clk = '1') then 
		if(reset = '1') then
			enable_1_reg <= '0';
		else
			enable_1_reg <= enable_1;
			if(enable_1_reg = '1') then
				dataout_1_reg <= dataout_1;
			end if;	
		end if;
	end if;
  end process;
  data_to_ulreg <= dataout_1 when (enable_1_reg = '1') else dataout_1_reg;

  bbdp: base_bank_dual_port 
		generic map ("dpram_1w_1r_1024x32_base_bank_dual_port",
					g_addr_width => 10, g_data_width => 32)
		port map (
			clk => clk, reset => reset,
			datain_0 => datain_0,
			dataout_0 => dataout_0,
         		addrin_0 => addrin_0,
         		enable_0 => enable_0,
         		writebar_0  => writebar_0 ,
	 		datain_1  => datain_1 ,
         		dataout_1 => dataout_1,
         		addrin_1 => addrin_1,
         		enable_1 => enable_1,
         		writebar_1  => writebar_1 
		);


   sfsm: SingleCycleStartFinFsm 
			port map (clk => clk, reset => reset,
					start_req => start_req, start_ack => start_ack,
						fin_req => ureg_write_ack, fin_ack => ureg_write_req,
							enable => enable_base);

   ureg: UnloadRegister 
		generic map (name => "dpram_1w_1r_1024x32_base_bank_dual_port:ureg",
				data_width => 32,
				  bypass_flag => true, nonblocking_read_flag => false)
		port map (write_data => data_to_ulreg,
				write_req => ureg_write_req,
					write_ack => ureg_write_ack,
					    read_data => read_data,
						unload_req => update_req,
						   unload_ack => update_ack,
							clk => clk,
							  reset => reset);

end dpram_1w_1r_1024x32_Operator_arch;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;


entity countDownTimer is -- 
    generic (tag_length : integer);
    port ( -- 
      time_count : in  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity countDownTimer;

architecture Behave of countDownTimer is
	type TimerState is (idle, busy, done);
	signal tstate : TimerState;
	signal count_sig : unsigned(31 downto 0);
	signal tag_reg: std_logic_vector(tag_length-1 downto 0);
begin

	process(clk,reset,tstate,count_sig,start_req,fin_req,tag_in)
		variable next_state: TimerState;
		variable latch_var, decr_count, latch_otag: boolean;
	begin
		next_state := tstate;

		start_ack <= '0';
		fin_ack <= '0';

		latch_var := false;
		decr_count := false;
		latch_otag := false;

		case tstate is 
			when idle =>
				start_ack <= '1';
				if(start_req = '1') then
					next_state := busy;
					latch_var  := true;
				end if;
			when busy =>
				decr_count := true;
				if(count_sig = 0) then
					next_state := done;
					latch_otag := true;
				end if;
			when done =>
				fin_ack <= '1';
				if(fin_req = '1') then
					next_state := idle;
				end if;
			when others =>
		end case;
		if(clk'event  and clk = '1') then
			if(reset = '1') then
				tstate <= idle;
			else
				tstate <= next_state;	
			end if;

			if(latch_var) then
				count_sig <= unsigned(time_count);
				tag_reg <= tag_in;
			elsif(decr_count) then
				count_sig <= count_sig - 1;
			end if;

			if(latch_otag) then
				tag_out <= tag_reg;	
			end if;
		end if;
	end process;

end Behave;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;


entity getClockTime is -- 
    generic (tag_length : integer);
    port ( -- 
      clock_time : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity getClockTime;

architecture Behave of getClockTime is

	type TimerState is (idle, done);
	signal tstate : TimerState;
	signal count_sig : unsigned(31 downto 0);

begin

	process(clk,reset,tstate,count_sig,start_req,fin_req,tag_in)
		variable next_state: TimerState;
		variable latch_var, decr_count, latch_otag: boolean;
	begin
		next_state := tstate;

		start_ack <= '0';
		fin_ack <= '0';

		latch_var := false;
		decr_count := false;

		case tstate is 
			when idle =>
				start_ack <= '1';
				if(start_req = '1') then
					next_state := done;
					latch_var  := true;
				end if;
			when done =>
				fin_ack <= '1';
				if(fin_req = '1') then
					next_state := idle;
				end if;
		end case;
		if(clk'event  and clk = '1') then
			if(reset = '1') then
				tstate <= idle;
				count_sig <= (others => '0');
			else
				tstate <= next_state;	
				count_sig <= count_sig + 1;
			end if;

			if(latch_var) then
				tag_out <= tag_in;
				clock_time <= std_logic_vector(count_sig);	
			end if;
		end if;
	end process;

end Behave;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;

entity uaddsub32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      carry_in: in std_logic_vector(0 downto 0);
      carry_out: out std_logic_vector(0 downto 0);
      subtract_flag: in std_logic_vector(0 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end entity uaddsub32_Operator;

architecture Struct of uaddsub32_Operator is
   signal pipeline_stall: std_logic;
   signal out_rdy_sig: std_logic;
   signal start_req, start_ack, fin_req, fin_ack: std_logic;
   signal tag_in, tag_out: std_logic_vector(0 downto 0);

   signal addsub_out, ret_val_x_x_reg : std_logic_vector(31 downto 0);
   signal update_ack_sig: boolean;
begin
   tag_in(0) <= '0';
   update_ack <= update_ack_sig;

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map(name => "uaddsub32-Operator-p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "uaddsub32-Operator-l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);
				

   pipeline_stall <= fin_ack and (not fin_req);
   start_ack <= not pipeline_stall;

   addsub_inst: UnsignedAdderSubtractor_n_n_n
		generic map( name => "uaddsub32-adder",
				tag_width => 1,
				operand_width => 32,
				chunk_width => 8)
		port map(slv_L => L,  slv_R => R, 
				slv_RESULT => addsub_out,
				slv_carry_in => carry_in(0),
				slv_carry_out => carry_out(0),
				subtract_op => subtract_flag(0),
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				stall => pipeline_stall,
				in_rdy => start_req, out_rdy => fin_ack);
   rrr: BypassRegister 
		generic map (data_width => 32, bypass => true)
		port map (clk => clk, reset => reset, enable => update_ack_sig, din => addsub_out, q => ret_val_x_x);
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;

entity uaddsub32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      carry_in: in std_logic_vector(0 downto 0);
      carry_out: out std_logic_vector(0 downto 0);
      subtract_flag: in std_logic_vector(0 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity uaddsub32;

architecture Struct of uaddsub32 is
   signal pipeline_stall: std_logic;
   signal out_rdy_sig: std_logic;
begin
   pipeline_stall <= out_rdy_sig and (not fin_req);
   start_ack <= not pipeline_stall;
   fin_ack <= out_rdy_sig;

   shift_inst: UnsignedAdderSubtractor_n_n_n
		generic map( name => "uaddsub32-adder",
				tag_width => tag_length,
				operand_width => 32,
				chunk_width => 8)
		port map(slv_L => L,  slv_R => R, 
				slv_RESULT => ret_val_x_x,
				slv_carry_in => carry_in(0),
				slv_carry_out => carry_out(0),
				subtract_op => subtract_flag(0),
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				stall => pipeline_stall,
				in_rdy => start_req, out_rdy => out_rdy_sig);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;


entity umul32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end entity umul32_Operator;

architecture Struct of umul32_Operator is
   signal in_data: std_logic_vector(63 downto 0);
   signal start_req, start_ack, fin_req, fin_ack: std_logic;
   signal tag_in, tag_out: std_logic_vector(0 downto 0);
   signal mul_out, ret_val_x_x_reg : std_logic_vector(63 downto 0);
   signal update_ack_sig: boolean;
begin
   tag_in(0) <= '0';
   update_ack <= update_ack_sig;

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map(name => "umul32_Operator_p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "umul32_Operator_l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);
				
   in_data <= L & R; -- concatenate..

   mul_inst: GenericApIntArithOperator
		generic map(op_id => "ApIntMul",
				name => "umul32-Operator-mul",
				tag_width => 1,
				in_operand_width => 32,
				num_non_constant_inputs => 2,
				first_operand_is_constant => false,
				second_operand_is_constant => false,
				constant_value => "0",
                   		out_result_width => 64)
		port map(in_data => in_data, 
				out_data => mul_out,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				op_i_rdy => start_ack, op_o_rdy => fin_ack);

			
   rrr: BypassRegister 
		generic map (data_width => 64, bypass => true)
		port map (clk => clk, reset =>reset, enable => update_ack_sig, din => mul_out, q => ret_val_x_x);
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;


entity umul32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity umul32;

architecture Struct of umul32 is
   signal in_data: std_logic_vector(63 downto 0);
begin
   in_data <= L & R; -- concatenate..

   mul_inst: GenericApIntArithOperator
		generic map(op_id => "ApIntMul",
				name => "umul32-mul",
				tag_width => tag_length,
				in_operand_width => 32,
				num_non_constant_inputs => 2,
				first_operand_is_constant => false,
				second_operand_is_constant => false,
				constant_value => "0",
                   		out_result_width => 64)
		port map(in_data => in_data, 
				out_data => ret_val_x_x,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				env_rdy => start_req, accept_rdy => fin_req,
				op_i_rdy => start_ack, op_o_rdy => fin_ack);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;


entity ushift32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      shift_right_flag: in std_logic_vector(0 downto 0);
      signed_flag: in std_logic_vector(0 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end entity ushift32_Operator;

architecture Struct of ushift32_Operator is
   signal pipeline_stall: std_logic;
   signal out_rdy_sig: std_logic;

   signal start_req, start_ack, fin_req, fin_ack: std_logic;
   signal tag_in, tag_out: std_logic_vector(0 downto 0);
   signal shift_out, ret_val_x_x_reg : std_logic_vector(31 downto 0);
   signal update_ack_sig: boolean;
begin

   tag_in(0) <= '0';
   update_ack <= update_ack_sig;

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map (name => "ushift32_Operator_p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map (name => "ushift32_Operator_l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);
				
   pipeline_stall <= fin_ack and (not fin_req);
   start_ack <= not pipeline_stall;

   shift_inst: UnsignedShifter_n_n_n
		generic map( name => "ushift32-shifter",
				tag_width => 1,
				operand_width => 32,
				shift_amount_width => 32)
		port map(slv_L => L,  slv_R => R, 
				slv_RESULT => shift_out,
				clk => clk, reset => reset,
				shift_right_flag => shift_right_flag(0),
				signed_flag => signed_flag(0),		
				tag_in => tag_in , tag_out => tag_out,
				stall => pipeline_stall,
				in_rdy => start_req, out_rdy => fin_ack);

   rrr: BypassRegister 
		generic map (data_width => 32, bypass => true)
		port map (clk => clk, reset =>reset, enable => update_ack_sig, din => shift_out, q => ret_val_x_x);

end Struct;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;


entity ushift32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      shift_right_flag: in std_logic_vector(0 downto 0);
      signed_flag: in std_logic_vector(0 downto 0);
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity ushift32;

architecture Struct of ushift32 is
   signal pipeline_stall: std_logic;
   signal out_rdy_sig: std_logic;
begin
   pipeline_stall <= out_rdy_sig and (not fin_req);
   start_ack <= not pipeline_stall;
   fin_ack <= out_rdy_sig;

   shift_inst: UnsignedShifter_n_n_n
		generic map( name => "ushift32-shifter",
				tag_width => tag_length,
				operand_width => 32,
				shift_amount_width => 32)
		port map(slv_L => L,  slv_R => R, 
				slv_RESULT => ret_val_x_x,
				clk => clk, reset => reset,
				shift_right_flag => shift_right_flag(0),
				signed_flag => signed_flag(0),		
				tag_in => tag_in , tag_out => tag_out,
				stall => pipeline_stall,
				in_rdy => start_req, out_rdy => out_rdy_sig);
			
end Struct;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- generic ap-int (signed/unsigned operator)
-- Madhav Desai.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;


-- 
-- mul/lshl/lshr/ashr.
-- 
entity GenericApIntArithOperator is
  generic (
	    name: string;
	    op_id: string;
	    tag_width : integer := 8;
	    in_operand_width: integer;
	    num_non_constant_inputs: integer;
            first_operand_is_constant: boolean;
            second_operand_is_constant: boolean;
	    constant_value: std_logic_vector;
	    out_result_width: integer
           );
  port(
    in_data: in std_logic_vector((num_non_constant_inputs*in_operand_width)-1 downto 0);
    out_data: out std_logic_vector(out_result_width-1 downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    env_rdy, accept_rdy: in std_logic;
    op_i_rdy, op_o_rdy: out std_logic);
end entity;

architecture rtl of GenericApIntArithOperator is

  signal pipeline_stall : std_logic;
  signal op_o_rdy_sig: std_logic;
  signal outR: std_logic_vector(out_result_width-1 downto 0);

begin

  assert (not (first_operand_is_constant and second_operand_is_constant))
	report "In " & " operator " & name & ", both operands are constants." severity failure;

  out_data <= outR;
  pipeline_stall <= op_o_rdy_sig and (not accept_rdy);
  op_o_rdy <= op_o_rdy_sig;
  op_i_rdy <= (not pipeline_stall);


  -- binary operator.
  arithOp: if ( (op_id = "ApIntMul") or
		(op_id = "ApIntSHL") or
		(op_id = "ApIntLSHR") or
		(op_id = "ApIntLASHR") or
		(op_id = "ApIntROL") or
		(op_id = "ApIntROR"))  generate
       gBlk: block
	signal inA, inB: std_logic_vector(in_operand_width-1 downto 0);
       begin
	     firstConstant: if (first_operand_is_constant) generate
	    	inA <= constant_value;
	     end generate firstConstant;

	     notfirstConstant: if (not first_operand_is_constant) generate
	    	inA <= in_data((2*in_operand_width)-1 downto in_operand_width);
	     end generate notfirstConstant;
	
	     secondConstant: if (second_operand_is_constant) generate
	    	inB <= constant_value;
	     end generate secondConstant;

	     notsecondConstant: if (not second_operand_is_constant) generate
	    	inB <= in_data(in_operand_width-1 downto 0);
             end generate notsecondConstant;

	     oprtr: GenericBinaryApIntArithOperatorPipelined
			generic map(name => name & ":binary" ,
					op_id => op_id,
					tag_width => tag_width,
					in_operand_width => in_operand_width,
					out_result_width => out_result_width)
			port map (inA => inA, inB => inB, outR => outR,
					pipeline_stall => pipeline_stall,
					tag_in => tag_in, tag_out => tag_out,
					env_rdy => env_rdy,
					op_o_rdy => op_o_rdy_sig,
					clk => clk, reset => reset);
       end block gBlk;
  end generate arithOp;

  notArithOp:if ( (op_id /= "ApIntMul") and
		(op_id /= "ApIntSHL") and
		(op_id /= "ApIntLSHR") and
		(op_id /= "ApIntLASHR"))  generate

 	assert false report op_id & " is not a pipelined binary arith operation" severity failure;

  end generate notArithOp;
end rtl;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- generic ap-int (signed/unsigned operator)
-- modified by Madhav Desai.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Subprograms.all;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;

entity GenericBinaryApIntArithOperatorPipelined is
  generic (
	    name : string;
	    op_id: string;
	    tag_width : integer := 8;
	    in_operand_width: integer;
	    out_result_width: integer
           );
  port(
    inA, inB: in std_logic_vector(in_operand_width-1 downto 0);
    outR: out std_logic_vector(out_result_width-1 downto 0);
    clk,reset: in std_logic;
    tag_in: in std_logic_vector(tag_width-1 downto 0);
    tag_out: out std_logic_vector(tag_width-1 downto 0);
    pipeline_stall: in std_logic;
    env_rdy: in std_logic;
    op_o_rdy: out std_logic);
end entity;

architecture rtl of GenericBinaryApIntArithOperatorPipelined is
begin


  -- binary operator.

  mulOp: if (op_id = "ApIntMul") generate
	op: UnsignedMultiplier_n_n_2n
		generic map (name => name & "-mul", 
				tag_width => tag_width,
				    operand_width => in_operand_width,
					chunk_width => 32)
		port map (
    				slv_L => inA,
				slv_R => inB,
    				slv_RESULT  => outR,
				clk => clk, 
				reset => reset,
    				in_rdy   => env_rdy,
    				out_rdy  => op_o_rdy,
    				stall    => pipeline_stall,
    				tag_in   => tag_in,
    				tag_out  => tag_out
			 );
  end generate mulOp;

  shiftOp: if ((op_id = "ApIntSHL") or (op_id = "ApIntLSHR") or (op_id = "ApIntASHR")) generate
    bb: block
       signal shift_right_flag: std_logic;
       signal signed_flag: std_logic;
    begin
	signed_flag <= '1' when (op_id = "ApIntASHR") else '0';
	shift_right_flag <= '1' when ((op_id = "ApIntLSHR") or (op_id = "ApIntASHR"))  else '0';

	op: UnsignedShifter_n_n_n
		generic map (
				name => name & "-shift",
				tag_width => tag_width,
				operand_width => in_operand_width,
				shift_amount_width => out_result_width
			    )
		port map (
				clk => clk, 
				reset => reset,
				slv_L => inA,
				slv_R => inB,
				slv_RESULT => outR,
				signed_flag => signed_flag,
				shift_right_flag => shift_right_flag,
				stall => pipeline_stall,
				tag_in => tag_in,
				tag_out => tag_out,
				in_rdy => env_rdy,
				out_rdy => op_o_rdy
			 );
    end block;
  end generate shiftOp;

  -- only mul and shifts here for now.
  assert ((op_id = "ApIntSHL") or (op_id = "ApIntLSHR") or (op_id = "ApIntASHR") or (op_id = "ApIntMul"))
	report "Currently unsupported operator " & op_id severity failure;

end rtl;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Types.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;
use ahir.BaseComponents.all;
use ahir.ApIntComponents.all;

entity PipelinedApIntOperator is
  generic (
      name : string;
      operator_id : string;
      no_arbitration: boolean := true;
      in_data_width: integer;
      out_data_width: integer;
      num_reqs : integer := 3; -- how many requesters?
      use_input_buffering: boolean := true;
      detailed_buffering_per_input: IntegerArray;
      detailed_buffering_per_output: IntegerArray;
      full_rate: boolean
    );
  port (
    -- req/ack follow level protocol
    reqL                     : in BooleanArray(num_reqs-1 downto 0);
    ackR                     : out BooleanArray(num_reqs-1 downto 0);
    ackL                     : out BooleanArray(num_reqs-1 downto 0);
    reqR                     : in  BooleanArray(num_reqs-1 downto 0);
    -- input data consists of concatenated pairs of ips
    dataL                    : in std_logic_vector((2*in_data_width*num_reqs)-1 downto 0);
    -- output data consists of concatenated pairs of ops.
    dataR                    : out std_logic_vector((out_data_width*num_reqs)-1 downto 0);
    -- with dataR
    clk, reset              : in std_logic);
end entity;

architecture Vanilla of PipelinedApIntOperator is

  constant num_operands : integer := 2;
  constant operand_width : integer := in_data_width;
  constant iwidth : integer := 2*operand_width;
  constant owidth : integer := out_data_width;
  
  constant tag_length: integer := Maximum(1,Ceil_Log2(reqL'length));
  signal itag,otag : std_logic_vector(tag_length-1 downto 0);
  signal ireq,iack, oreq, oack: std_logic;

  constant debug_flag : boolean := global_debug_flag;

  signal idata: std_logic_vector(iwidth-1 downto 0);
  signal odata: std_logic_vector(owidth-1 downto 0);
begin  -- Behave

  assert ackL'length = reqL'length report "mismatched req/ack vectors" severity error;
  assert ((operand_width = 32) or (operand_width = 64)) report "32/64 bit operand-support only!" severity error;
  assert ((operator_id = "ApFloatMul") or (operator_id = "ApFloatAdd") or (operator_id = "ApFloatSub"))
    report "operator_id must be either add or mul or sub" severity error;  

  -- DebugGen: if debug_flag generate 
    -- assert( (not ((reset = '0') and (clk'event and clk = '1') and no_arbitration)) or Is_At_Most_One_Hot(reqL))
    -- report "in no-arbitration case, at most one request should be hot on clock edge (in SplitOperatorShared)" severity error;
  -- end generate DebugGen;
  NoInBuffers : if not use_input_buffering generate 
    imux: InputMuxBase
      generic map(name => name & "-imux",
		  iwidth => iwidth*num_reqs,
                  owidth => iwidth, 
                  twidth => tag_length,
                  nreqs => num_reqs,
                  no_arbitration => no_arbitration,
                  registered_output => false)
      port map(
          reqL       => reqL,
        ackL       => ackL,
        reqR       => ireq,
        ackR       => iack,
        dataL      => dataL,
        dataR      => idata,
        tagR       => itag,
        clk        => clk,
        reset      => reset);
   end generate NoInBuffers;

  InBuffers: if use_input_buffering generate
    imuxWithInputBuf: InputMuxWithBuffering
      generic map(name => name & "-imux" , 
		iwidth => iwidth*num_reqs,
                owidth => iwidth, 
                twidth => tag_length,
                nreqs => num_reqs,
		buffering => detailed_buffering_per_input,
                no_arbitration => no_arbitration,
		full_rate => full_rate,
                registered_output => false)
      port map(
        reqL       => reqL,
        ackL       => ackL,
        reqR       => ireq,
        ackR       => iack,
        dataL      => dataL,
        dataR      => idata,
        tagR       => itag,
        clk        => clk,
        reset      => reset);
  end generate InBuffers;

   pipeOp: GenericApIntArithOperator
		generic map(name => name & "-int-operator", op_id => operator_id,
				tag_width => tag_length,
				 in_operand_width => in_data_width,
					num_non_constant_inputs => 0,	
					   first_operand_is_constant => false,
					    second_operand_is_constant => false,
						constant_value => "",
						out_result_width => out_data_width)
		port map ( in_data => idata,
    				out_data => odata,
    				clk => clk,
				reset => reset,
    				tag_in => itag,
    				tag_out => otag,
    				env_rdy => ireq,
		        	accept_rdy => oack, 
    				op_i_rdy => iack,
				op_o_rdy => oreq);


  odemux: OutputDeMuxBaseWithBuffering
    generic map (
        name => name & "-odemux",
  	iwidth => owidth,
  	owidth =>  owidth*num_reqs,
	twidth =>  tag_length,
	nreqs  => num_reqs,
	detailed_buffering_per_output => detailed_buffering_per_output,
	full_rate => full_rate)
    port map (
      reqL   => oreq,
      ackL   => oack,
      dataL => odata,
      tagL  => otag,
      reqR  => reqR,
      ackR  => ackR,
      dataR => dataR,
      clk   => clk,
      reset => reset);
  
end Vanilla;

------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- a basic unsigned adder..  if addition is specified, just
-- adds using a simple carry lookahead scheme.  if subtraction
-- is specified, takes the twos complement of the second operand
-- and adds the two numbers.  No overflow/negative checks
-- are performed.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;

entity AddSubCellX  is
	generic (operand_width: integer);
	port (A,B: in unsigned(operand_width-1 downto 0);
		Sum: out unsigned(operand_width-1 downto 0);
		BP,BG: out std_logic;
		stall: in std_logic;
		clk, reset: in std_logic);
end entity AddSubCellX;

architecture Behave of AddSubCellX is
begin
	process(clk, reset, A, B, stall )
		variable sumv: unsigned(operand_width-1 downto 0);
		variable prop, gen: std_logic;
	begin
		prop := '1';
		gen  := '0';

		sumv := A+B;

		for I in 0 to operand_width-1 loop
			prop := (prop and (A(I) or B(I)));
			gen  := (A(I) and B(I)) or (gen and (A(I) or B(I)));
		end loop;


		if(clk'event and clk = '1') then
		   if(stall = '0') then
			Sum <= sumv;
			BP <= prop;
			BG <= gen;
		   end if;
		end if;
	end process;
end Behave;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.SubPrograms.all;

entity UnsignedAdderSubtractor_n_n_n is
  
  generic (
    name : string;
    tag_width          : integer;
    operand_width      : integer;
    chunk_width        : integer
	);

  port (
    slv_L            : in  std_logic_vector(operand_width-1 downto 0);
    slv_R            : in  std_logic_vector(operand_width-1 downto 0);
    slv_RESULT       : out std_logic_vector(operand_width-1 downto 0);
    slv_carry_out    : out std_logic;
    slv_carry_in     : in std_logic;  
    subtract_op      : in std_logic;
    clk, reset       : in  std_logic;
    in_rdy           : in  std_logic;
    out_rdy          : out std_logic;
    stall            : in std_logic;
    tag_in           : in std_logic_vector(tag_width-1 downto 0);
    tag_out          : out std_logic_vector(tag_width-1 downto 0));

end entity;


architecture Pipelined of UnsignedAdderSubtractor_n_n_n is
 
  constant num_chunks: integer := Ceil(operand_width, chunk_width);
  constant padded_operand_width: integer := num_chunks  * chunk_width;
  signal Lpadded, Rpadded, Resultpadded : unsigned(padded_operand_width-1 downto 0);

  constant pipe_depth : integer := 3;
  signal stage_active : std_logic_vector(0 to pipe_depth);


  type CWORD is array (natural range <>) of unsigned(chunk_width-1 downto 0);
  type TWORD is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);  
  signal stage_tags: TWORD(0 to pipe_depth);


  signal addsubcell_Sum, addsubcell_Sum_Delayed, 
			addsubcell_A, addsubcell_B, final_sums: CWord(0 to num_chunks-1);
  signal addsubcell_BP, addsubcell_BG : std_logic_vector(0 to num_chunks-1);

  signal block_carries: std_logic_vector(0 to num_chunks);
  signal subtract_op_1, subtract_op_2: std_logic;

  component AddSubCellX  is
	generic ( operand_width: integer);
	port (A,B: in unsigned(operand_width-1 downto 0);
		Sum: out unsigned(operand_width-1 downto 0);
		BP,BG: out std_logic;
		stall: in std_logic;
		clk, reset: in std_logic);
  end component AddSubCellX;
   
  signal L             : unsigned(operand_width-1 downto 0);
  signal R             : unsigned(operand_width-1 downto 0);
  signal RESULT        : unsigned(operand_width-1 downto 0);
  signal lsChunk_carry_in : std_logic;
  
begin  -- Pipelined

  -- slv <-> unsigned
  L <= To_Unsigned(slv_L);
  R <= To_Unsigned(slv_R);
  slv_RESULT <= To_SLV(RESULT);


  stage_active(0) <= in_rdy;
  out_rdy <= stage_active(pipe_depth);
  stage_tags(0) <= tag_in;
  tag_out <= stage_tags(3);

  RESULT <= ResultPadded(operand_width-1 downto 0);


  -- note: if subtract_op = '1', then complement R (see below) and add 1.
  -- pad. also if subtract_op = '1' then complement R and add 1 addsubcell_Cin).
  process(L,R,subtract_op)
	variable ltmp, rtmp: unsigned(padded_operand_width-1 downto 0);
	variable sign_bit : std_logic;
  begin
        
	ltmp := (others => L(operand_width-1)); ltmp(operand_width-1 downto 0) := L;
	rtmp := (others => R(operand_width-1)); rtmp(operand_width-1 downto 0) := R;
	Lpadded <= ltmp;

	if(subtract_op = '0') then
		Rpadded <= rtmp;
	else
		Rpadded <= not rtmp;
	end if;
  end process;

  -- carry into least significant block.
  lsChunk_carry_in <=  '1' when ((slv_carry_in = '1') xor (subtract_op = '1')) else '0';
  
  Stage1:  for I in  0 to num_chunks-1 generate

	addsubcell_A(I) <= Lpadded(((I+1)*chunk_width)-1 downto (I*chunk_width));
	addsubcell_B(I) <= Rpadded(((I+1)*chunk_width)-1 downto (I*chunk_width));

	asCellX: AddSubCellX generic map(operand_width => chunk_width)
		port  map( A => addsubcell_A(I),
			   B => addsubcell_B(I),	
			   Sum => addsubcell_Sum(I),
			   BP => addsubcell_BP(I),
			   BG => addsubcell_BG(I),
			   stall => stall,
			   clk => clk,
			   reset => reset);
  end generate Stage1;

  process(clk)
  begin
	if(clk'event and clk = '1') then
		if(stall = '0') then
			stage_tags(1) <= stage_tags(0);
			subtract_op_1 <= subtract_op;
		end if;
		if(reset = '1') then
			stage_active(1) <= '0';
		elsif stall = '0' then
			stage_active(1) <= stage_active(0);
		end if;
	end if;
  end process;

  -- stage two: calculate the block carries.
  process(clk, reset, stall, stage_active, lsChunk_carry_in, addsubcell_Sum, addsubcell_BP, addsubcell_BG)	
	variable cin: std_logic_vector(0 to num_chunks);
  begin
	cin(0) := lsChunk_carry_in;
	for I in 1 to num_chunks loop
		cin(I) := (cin(I-1) and addsubcell_BP(I-1))  or addsubcell_BG(I-1);
	end loop;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			stage_active(2) <= '0';
		elsif(stall = '0') then
			block_carries <= cin;
			stage_tags(2) <= stage_tags(1);
			addsubcell_Sum_Delayed <= addsubcell_Sum;
			subtract_op_2 <= subtract_op_1;
			stage_active(2) <= stage_active(1);
		end if;
	end if;
  end process;


  -- stage three: final sums
  process(clk)
	variable correction, tmp: unsigned(chunk_width-1 downto 0);
	variable is_negative: boolean;
  begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			stage_active(3) <= '0';
		elsif(stall = '0') then
			for I in 0 to num_chunks-1 loop
				correction := (others => '0');
				if(block_carries(I) = '1') then
					correction(0) := '1';
				end if;
				final_sums(I) <= addsubcell_Sum_Delayed(I) + correction;
			end loop;

			stage_tags(3) <= stage_tags(2);
			stage_active(3) <= stage_active(2);
		end if;
	end if;
  end process;


  -- collect final-sums into RESULT
  process(final_sums)
  begin
	for I in 0 to num_chunks-1 loop
		ResultPadded(((I+1)*chunk_width)-1 downto (I*chunk_width)) <= final_sums(I);
	end loop;
  end process;



end Pipelined;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- a basic unsigned multiplier.
--    basic architecture
--    pipelined array multiplier
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity DelayCellX is
   generic (operand_width: integer; delay: natural);
   port (Din: in unsigned(operand_width-1 downto 0);
	 Dout: out unsigned(operand_width-1 downto 0);
	 clk: in std_logic;
	 stall: in std_logic);
end entity DelayCellX;

architecture Behave of DelayCellX is
	type DArray is array (natural range <>) of unsigned(operand_width-1 downto 0);
	signal data_array: DArray(0 to delay);
begin

	data_array(0) <= Din;
	NonZeroDelay: if delay > 0 generate
	   SRgen: for I in 1 to delay generate
		process(clk)
		begin
			if(clk'event and clk = '1') then
				if(stall = '0') then
					data_array(I) <= data_array(I-1);
				end if;
			end if;
			
		end process;
	    end generate SRgen;
	end generate NonZeroDelay;
	
	Dout <= data_array(delay);
end Behave;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SumCellX is
 	generic (operand_width: integer; ignore_diag: boolean; ignore_right: boolean);
	port (SU,SDiagIn: in unsigned(operand_width-1 downto 0);
              SR: in unsigned(1 downto 0);
	      SDiagOut: out unsigned(operand_width-1 downto 0);
	      SL: out unsigned(1 downto 0);
	      stall: in std_logic;
	      clk: in std_logic);
end entity SumCellX;

architecture Behave of SumCellX is
begin

	process(clk)
		variable x, y, z, sum: unsigned(operand_width+1 downto 0);
		variable t: unsigned(1 downto 0);
	begin

		if(clk'event and clk = '1') then
			if(stall = '0') then
				x := "00" & SU;
				y := (1 => SR(1), 0 => SR(0), others => '0');
				z := "00" & SDiagIn;
		
				if(not (ignore_diag  or ignore_right)) then
					sum := x + y + z;
				elsif (ignore_diag and ignore_right) then
					sum := x;
				elsif (ignore_diag and (not ignore_right)) then
					sum := (x + y);
				else
					sum := (x + z);
				end if;
	
				t := sum(operand_width+1 downto operand_width);

				SDiagOut <= sum(operand_width-1 downto 0);
				SL <= t;
			end if;
		end if;
	end process;
end Behave;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MultiplierCellX is
  generic (operand_width: integer);
  port (MT, MR, ST, DiagIn: in unsigned(operand_width-1 downto 0);
        ML, MD, SD, DiagOut: out unsigned(operand_width-1 downto 0);
        stall: in std_logic;
	clk: in std_logic);
end entity MultiplierCellX;

architecture Simple of MultiplierCellX is
	constant zero_const : unsigned(operand_width-2 downto 0) := (others => '0');
begin

	-- sent through without any delay.
	ML <= MR;

	process(clk)
		variable tmp,wext: unsigned((2*operand_width)-1 downto 0);
		variable u, v, w: unsigned(operand_width downto 0);
	begin
		if(clk'event and clk = '1') then
			if(stall = '0') then
				tmp := MT*MR;
		
				-- pad one bit to incoming summands.
				u :=  "0" & DiagIn;
                                v :=  "0" & ST;
		
				-- this is a operand_width+1 size addition
				w := (u + v);

				-- pad to 2*operand_width
				wext := zero_const & w;
		
				-- a full 2*operand_width addition.
				tmp := tmp + wext;

				-- send down the vertical operand
				-- with a cycle delay.
				MD <= MT;

				-- top half of result goes down to 
				-- next row (to be summed)
				SD <= tmp((2*operand_width)-1 downto operand_width);

				-- bottom half of the result goes out
				-- on the diagonal..
				DiagOut <= tmp(operand_width-1 downto 0);
			end if;
		end if;
	end process;
end Simple;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.Utilities.all;
use ahir.SubPrograms.all;

entity UnsignedMultiplier_n_n_2n is
  
  generic (
    name: string;
    tag_width     : integer;
    operand_width : integer;
    chunk_width   : integer := 16);

  port (
    slv_L, slv_R       : in  std_logic_vector(operand_width-1 downto 0);
    slv_RESULT     : out std_logic_vector((2*operand_width)-1 downto 0);
    clk, reset : in  std_logic;
    in_rdy     : in  std_logic;
    out_rdy    : out std_logic;
    stall      : in std_logic;
    tag_in     : in std_logic_vector(tag_width-1 downto 0);
    tag_out    : out std_logic_vector(tag_width-1 downto 0));
end entity;

architecture Pipelined of UnsignedMultiplier_n_n_2n is

  constant pipe_depth : integer := operand_width/chunk_width;

  type RWORD is array (natural range <>) of unsigned((2*operand_width)-1 downto 0);
  type TWORD is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);  


  signal intermediate_results : RWORD(0 to pipe_depth);
  signal intermediate_tags : TWORD(0 to pipe_depth);  
  signal stage_active : std_logic_vector(0 to pipe_depth);
  
  signal L,R: unsigned (operand_width-1 downto 0);
  signal RESULT: unsigned((2*operand_width)-1 downto 0);

begin  -- Pipelined

  -- unsigned <-> slv
  L <= To_Unsigned(slv_L);
  R <= To_Unsigned(slv_R);
  slv_RESULT <= To_SLV(RESULT);
  
  -- for now, just multiply..
  intermediate_results(0) <= L*R;


  -- I/O
  intermediate_tags(0) <= tag_in;
  stage_active(0) <= in_rdy;
  out_rdy <= stage_active(pipe_depth);
  tag_out <= intermediate_tags(pipe_depth);
  RESULT <= intermediate_results(pipe_depth);
  
  -- for now, just add stages after the multiply
  -- the synthesis tool should retime.  Later
  -- we'll get around to doing the array multiplier
  -- right.
  Pipeline: for STAGE in 1 to pipe_depth generate

    process(clk)
    begin
      if(clk'event and clk = '1') then
        if(reset = '1') then
          stage_active(STAGE) <= '0';
        elsif(stall = '0') then
          stage_active(STAGE) <= stage_active(STAGE-1);
        end if;

        if(stall = '0') then
          intermediate_results(STAGE) <= intermediate_results(STAGE-1);
          intermediate_tags(STAGE) <= intermediate_tags(STAGE-1);
        end if;
        
      end if;
    end process;
    
  end generate Pipeline;
end Pipelined;


 
architecture ArrayMul of UnsignedMultiplier_n_n_2n is

	constant NumChunks : integer := Ceil(operand_width, chunk_width);

	constant padded_operand_width: integer  := NumChunks*chunk_width;
	signal Lpadded, Rpadded: unsigned(padded_operand_width-1 downto 0);
	signal RESULTpadded: unsigned((2*padded_operand_width)-1 downto 0);

	type TwoDTagArray is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);
	signal tag_array: TwoDTagArray(0 to 2*NumChunks);

	type TwoDChunkArray is array (natural range <>, natural range <>) of unsigned(chunk_width-1 downto 0);
	signal MT, ML, ST, DiagIn, SD, MR, MD, DiagOut: TwoDChunkArray(0 to NumChunks-1, 0 to NumChunks-1);



	signal rdy_array: std_logic_vector(0 to 2*NumChunks);

        -- the multiplier cells are arranged in a NumChunk X NumChunk array.
        -- CellX (I,J) receives R(I) (MT),  L(J) (MR) and a partial sum from above (ST).
	-- CellX (I,J) receives an incoming diagonal sum from CellX (I-1,J+1) and
        -- passes on its sum to the diagonal block CellX (I+1,J-1).
	--
	component DelayCellX 
   		generic (operand_width: integer; delay: natural);
   		port (Din: in unsigned(operand_width-1 downto 0);
	 		Dout: out unsigned(operand_width-1 downto 0);
	 		clk: in std_logic;
	 		stall: in std_logic);
	end component DelayCellX;

	component MultiplierCellX is
  		generic (operand_width: integer);
  		port (MT, MR, ST, DiagIn: in unsigned(operand_width-1 downto 0);
        		ML, MD, SD, DiagOut: out unsigned(operand_width-1 downto 0);
        		stall: in std_logic;
			clk: in std_logic);
	end component MultiplierCellX;

	component SumCellX is
 		generic (operand_width: integer; ignore_diag: boolean; ignore_right: boolean);
		port (SU,SDiagIn: in unsigned(operand_width-1 downto 0);
              		SR: in unsigned(1 downto 0);
	      		SDiagOut: out unsigned(operand_width-1 downto 0);
	      		SL: out unsigned(1 downto 0);
	      		stall: in std_logic;
	      		clk: in std_logic);
	end component SumCellX;

	type OneDChunkArray is array (natural range <>) of unsigned(chunk_width-1 downto 0);
	signal SU,SDiagIn,SDiagOut: OneDChunkArray(0 to NumChunks-1);

	type OneD2BitArray is array (natural range <>) of unsigned(1 downto 0);
        signal SR,SL: OneD2BitArray(0 to NumChunks-1);

	signal result_array : OneDChunkArray(0 to (2*NumChunks)-1);
  
	signal L,R: unsigned (operand_width-1 downto 0);
  	signal RESULT: unsigned((2*operand_width)-1 downto 0);
begin
  	-- unsigned <-> slv
  	L <= To_Unsigned(slv_L);
  	R <= To_Unsigned(slv_R);
  	slv_RESULT <= To_SLV(RESULT);

	process(L)
		variable lpad : unsigned(padded_operand_width-1 downto 0);
	begin
		lpad := (others => '0');
		lpad(operand_width-1 downto 0) := L;
		Lpadded <= lpad;
	end process;

	process(R)
		variable rpad : unsigned(padded_operand_width-1 downto 0);
	begin
		rpad := (others => '0');
		rpad(operand_width-1 downto 0) := R;
		Rpadded <= rpad;
	end process;

	RESULT <= RESULTpadded((2*operand_width)-1 downto 0);

	tag_array(0) <= tag_in;
	rdy_array(0) <= in_rdy;
	
	Tags: for ROW in 1 to (2*NumChunks) generate
		process(clk)
		begin
			if(clk'event and clk = '1') then
				if(reset = '1') then
					rdy_array(ROW) <= '0';
					tag_array(ROW) <= (others => '0');
				elsif(stall = '0') then
					tag_array(ROW) <= tag_array(ROW-1);
					rdy_array(ROW) <= rdy_array(ROW-1);
				end if;
			end if;
		end process;
	end generate Tags;
	tag_out <= tag_array(2*NumChunks);
	out_rdy <= rdy_array(2*NumChunks);

	Rows: for ROW in 0 to NumChunks-1 generate
		Cols: for COL in 0 to NumChunks-1 generate

			-- incoming  L values get into MT(0,-).
			ROWBC: if ROW = 0 generate
                                MT(ROW,COL) <= Lpadded(((COL+1)*chunk_width)-1 downto (COL*chunk_width));

				-- incoming signals to top row are 0.
				DiagIn(ROW,COL) <= (others => '0');
				ST(ROW,COL) <= (others => '0');

			end generate ROWBC;

		        COLBC: if COL=NumChunks-1 and ROW>0 generate
				-- left border column has incoming diagonals 0
				DiagIn(ROW,COL) <= (others => '0');
			end generate COLBC;

			-- from the right, R values enter with each row 
			-- getting an appropriate delay.
			COLBC2: if COL = 0 generate
				delInst: DelayCellX generic map(operand_width => chunk_width,
								delay => ROW)
					port map(Din => Rpadded(((ROW+1)*chunk_width)-1 downto (ROW*chunk_width)),
						 Dout => MR(ROW,COL),
						 clk => clk,
						 stall => stall);
			end generate COLBC2;

			-- passing from right to left.
			Cols1: if COL > 0 generate
				MR(ROW,COL) <= ML(ROW,COL-1);
			end generate Cols1;

			ConnectArray: if ROW>0 generate

				-- from top to bottom
				MT(ROW,COL) <= MD(ROW-1,COL);
				ST(ROW,COL) <= SD(ROW-1,COL);
				
				-- diagonally.
				Cols2: if COL < NumChunks-1 generate
					DiagIn(ROW,COL) <= DiagOut(ROW-1,COL+1);
				end generate Cols2;
			end generate ConnectArray;

			mulCellX: MultiplierCellX generic map(operand_width => chunk_width)
				port map(MT => MT(ROW,COL),
					 ML => ML(ROW,COL),
					 ST => ST(ROW,COL),
					 DiagIn => DiagIn(ROW,COL),
					 SD => SD(ROW,COL),
					 MR => MR(ROW,COL),
					 MD => MD(ROW,COL),
					 stall => stall,
					 DiagOut => DiagOut(ROW,COL),
					 clk => clk);
		end generate Cols;
	end generate Rows;


	--  instantiate an array of sum cells to take
	--  care of the SD correction.
	sumArray: for Cols in 0 to NumChunks-1 generate
	
		scell: SumCellX generic map (operand_width => chunk_width,
						ignore_diag => (Cols = NumChunks-1),
						ignore_right => (Cols = 0))
			port map(SU => SU(Cols),
				 SDiagIn => SDiagIn(Cols),
				 SR => SR(Cols),
				 SDiagOut => SDiagOut(Cols),
				 SL => SL(Cols),
				 stall => stall,
				 clk => clk);

		BR: if(Cols = 0) generate
			-- 0s from the right at the right boundary
			SR(Cols) <= (others => '0');
		end generate BR;
				
		BL: if(Cols = NumChunks-1) generate
			-- 0s from the diagonal at the left boundary.
			SDiagIn(Cols) <= (others => '0');
		end generate BL;

		--   inputs to the cells are delayed to match the sum
		--   propagation.

		--  sum coming down..
		dSU: DelayCellX generic map(operand_width => chunk_width, delay => Cols)
			port map(Din => SD(NumChunks-1,Cols),
				 Dout => SU(Cols),
				 clk => clk,
				 stall => stall);
		
		Cntr1: if(Cols > 0) generate
			SR(Cols) <= SL(Cols-1);
		end generate Cntr1;
		
		Cntr2: if (Cols < NumChunks-1) generate
			-- diagonal coming in..  the leftmost cell has no incoming diagonal.
			dSDiagIn: DelayCellX generic map(operand_width => chunk_width, delay => Cols)
				port map(Din => DiagOut(NumChunks-1,Cols+1),
				 Dout => SDiagIn(Cols),
				 clk => clk,
				 stall => stall);
		end generate Cntr2;
		
	end generate sumArray;


	--       instantiate delay elements to match delays
        --       inserted due to sum-cell array.


	-- the right column and 2*N-1 delays inserted.
	RightColumn:  for Rows in 0 to NumChunks-1 generate
		dRc: DelayCellX generic map(operand_width => chunk_width, delay => ((2*NumChunks)-1)-Rows)
			port map(Din => DiagOut(Rows,0),
				 Dout => result_array(Rows),
				 stall => stall,
				 clk => clk);
	end generate RightColumn;

	-- the bottom row as N-C delays inserted as C goes from 0 to N-2
	BottomRow: for Cols in 0 to NumChunks-2 generate
		dBr: DelayCellX generic map(operand_width => chunk_width, delay => NumChunks-(Cols+1))
			port map(Din => SDiagOut(Cols),
				 Dout => result_array(Cols+NumChunks),
				 stall => stall,
				 clk => clk);
		
	end generate BottomRow;

	-- leftmost element has no delays inserted.
	result_array((2*NumChunks)-1) <= SDiagOut(NumChunks-1);


	-- result: pack the diagonals into the result vector.
	process(result_array)
	begin
		for I in 0 to (2*NumChunks)-1 loop
			RESULTpadded(((I+1)*chunk_width)-1 downto (I*chunk_width))
				<= result_array(I);
		end loop;
	end process;

end ArrayMul;
------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- a basic unsigned shifter.
--
-- for the moment, this just does a shift and adds delay stages at
-- the end; presumably, the synthesis tool will retime things
-- appropriately..
--
-- TODO: pipeline this explicitly!
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.GlobalConstants.all;
use ahir.Utilities.all;
use ahir.SubPrograms.all;

entity UnsignedShifter_n_n_n is
  generic (
    name: string;
    tag_width          : integer;
    operand_width      : integer;
    shift_amount_width : integer);

  port (
    slv_L       : in  std_logic_vector(operand_width-1 downto 0);
    slv_R       : in  std_logic_vector(shift_amount_width-1 downto 0);
    slv_RESULT  : out std_logic_vector(operand_width-1 downto 0);
    clk, reset  : in  std_logic;
    in_rdy      : in  std_logic;
    out_rdy     : out std_logic;
    shift_right_flag : in std_logic;
    signed_flag : in std_logic;
    stall       : in std_logic;
    tag_in      : in std_logic_vector(tag_width-1 downto 0);
    tag_out     : out std_logic_vector(tag_width-1 downto 0));

end entity;


architecture Pipelined of UnsignedShifter_n_n_n is

  -- depth of multiplexor..
  constant phases_per_stage: integer := 8;

  constant num_sig_bits: integer := Maximum(1,Minimum(shift_amount_width, Ceil_Log2(operand_width)));
  constant pipe_depth : integer := Ceil(num_sig_bits,phases_per_stage);

  type RWORD is array (natural range <>) of std_logic_vector(operand_width-1 downto 0);
  type TWORD is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);  

  type SWORD is array (natural range <>) of unsigned(num_sig_bits-1 downto 0);  

  signal intermediate_results : RWORD(0 to pipe_depth);
  signal intermediate_tags : TWORD(0 to pipe_depth);  
  signal intermediate_shift_amount : SWORD(0 to pipe_depth);  
  signal stage_active : std_logic_vector(0 to pipe_depth);

  
  constant debug_flag: boolean := global_debug_flag;

  function shift_right_signed ( X: std_logic_vector; Y: integer )
		return std_logic_vector is
	variable ret_val: std_logic_vector(1 to X'length);
  begin
	ret_val := To_SLV( shift_right(To_Signed(X),Y));
	return(ret_val);
  end shift_right_signed;

  function shift_right_unsigned ( X: std_logic_vector; Y: integer )
		return std_logic_vector is
	variable ret_val: std_logic_vector(1 to X'length);
  begin
	ret_val := To_SLV(shift_right(To_Unsigned(X),Y));
	return(ret_val);
  end shift_right_unsigned;

  constant ZZZ: std_logic_vector(operand_width-1 downto 0) := (others => '0');

begin  -- Pipelined


   
  TrivOp: if operand_width = 1 generate
	intermediate_results(0) <= (others => '0') when (slv_R /= ZZZ) else slv_L;
  end generate TrivOp;
  

  NonTrivOp: if operand_width > 1 generate

        genStages: for STAGE in 1 to pipe_depth generate
  		process(clk, reset, signed_flag, intermediate_results, intermediate_shift_amount, shift_right_flag)
			variable shifted_L: std_logic_vector(operand_width-1 downto 0);
			variable shift_amount: unsigned(num_sig_bits-1 downto 0);
  		begin
			shifted_L := intermediate_results(STAGE-1);
			shift_amount := intermediate_shift_amount(STAGE-1);

			for I in ((STAGE-1)*phases_per_stage) to 
					Minimum(num_sig_bits-1,(STAGE*phases_per_stage)-1) loop  
				if(shift_amount(I) = '1') then
					if(shift_right_flag = '1') then
						if(signed_flag = '1') then
							shifted_L := shift_right_signed(shifted_L, 2**I);
						else 
							shifted_L := shift_right_unsigned(shifted_L, 2**I);
						end if;
					else
						shifted_L :=  To_SLV(shift_left(To_Unsigned(shifted_L),2**I));
					end if;
				end if;
			end loop;

			if(clk'event and clk='1') then

                                if(reset = '1') then
					stage_active(STAGE) <=  '0';
				elsif stall = '0' then
					stage_active(STAGE) <= stage_active(STAGE-1);
  					intermediate_results(STAGE) <= shifted_L;
  					intermediate_tags(STAGE) <= intermediate_tags(STAGE-1);
					intermediate_shift_amount(STAGE) <= 
							intermediate_shift_amount(STAGE-1);
				end if;
			end if;
  		end process;
	end generate genStages;

  end generate NonTrivOp;


  -- I/O
  intermediate_results(0) <=  slv_L;
  intermediate_tags(0) <= tag_in;
  intermediate_shift_amount(0) <= To_Unsigned(slv_R(num_sig_bits-1 downto 0));
  stage_active(0) <= in_rdy;
  out_rdy <= stage_active(pipe_depth);
  tag_out <= intermediate_tags(pipe_depth);
  slv_RESULT <= intermediate_results(pipe_depth);
  
end Pipelined;
