
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.types.all;
use ahir.components.all;

entity test_floats_cp is
  port(
    LambdaIn : in BooleanArray(323 downto 1);
    LambdaOut : out BooleanArray(323 downto 1);
    clk : in std_logic;
    reset : in std_logic);
end test_floats_cp;

architecture default_arch of test_floats_cp is
  signal place_0_preds : BooleanArray(0 downto 0);
  signal place_0_succs : BooleanArray(0 downto 0);
  signal place_0_token : boolean;
  signal place_5_preds : BooleanArray(0 downto 0);
  signal place_5_succs : BooleanArray(0 downto 0);
  signal place_5_token : boolean;
  signal place_12_preds : BooleanArray(0 downto 0);
  signal place_12_succs : BooleanArray(0 downto 0);
  signal place_12_token : boolean;
  signal place_13_preds : BooleanArray(0 downto 0);
  signal place_13_succs : BooleanArray(0 downto 0);
  signal place_13_token : boolean;
  signal place_14_preds : BooleanArray(0 downto 0);
  signal place_14_succs : BooleanArray(0 downto 0);
  signal place_14_token : boolean;
  signal place_19_preds : BooleanArray(0 downto 0);
  signal place_19_succs : BooleanArray(0 downto 0);
  signal place_19_token : boolean;
  signal place_20_preds : BooleanArray(0 downto 0);
  signal place_20_succs : BooleanArray(0 downto 0);
  signal place_20_token : boolean;
  signal place_21_preds : BooleanArray(0 downto 0);
  signal place_21_succs : BooleanArray(0 downto 0);
  signal place_21_token : boolean;
  signal place_26_preds : BooleanArray(0 downto 0);
  signal place_26_succs : BooleanArray(0 downto 0);
  signal place_26_token : boolean;
  signal place_27_preds : BooleanArray(0 downto 0);
  signal place_27_succs : BooleanArray(0 downto 0);
  signal place_27_token : boolean;
  signal place_28_preds : BooleanArray(0 downto 0);
  signal place_28_succs : BooleanArray(0 downto 0);
  signal place_28_token : boolean;
  signal place_34_preds : BooleanArray(0 downto 0);
  signal place_34_succs : BooleanArray(0 downto 0);
  signal place_34_token : boolean;
  signal place_35_preds : BooleanArray(0 downto 0);
  signal place_35_succs : BooleanArray(0 downto 0);
  signal place_35_token : boolean;
  signal place_36_preds : BooleanArray(0 downto 0);
  signal place_36_succs : BooleanArray(0 downto 0);
  signal place_36_token : boolean;
  signal place_41_preds : BooleanArray(0 downto 0);
  signal place_41_succs : BooleanArray(0 downto 0);
  signal place_41_token : boolean;
  signal place_42_preds : BooleanArray(0 downto 0);
  signal place_42_succs : BooleanArray(0 downto 0);
  signal place_42_token : boolean;
  signal place_43_preds : BooleanArray(0 downto 0);
  signal place_43_succs : BooleanArray(0 downto 0);
  signal place_43_token : boolean;
  signal place_49_preds : BooleanArray(0 downto 0);
  signal place_49_succs : BooleanArray(0 downto 0);
  signal place_49_token : boolean;
  signal place_50_preds : BooleanArray(0 downto 0);
  signal place_50_succs : BooleanArray(0 downto 0);
  signal place_50_token : boolean;
  signal place_51_preds : BooleanArray(0 downto 0);
  signal place_51_succs : BooleanArray(0 downto 0);
  signal place_51_token : boolean;
  signal place_52_preds : BooleanArray(0 downto 0);
  signal place_52_succs : BooleanArray(0 downto 0);
  signal place_52_token : boolean;
  signal place_56_preds : BooleanArray(0 downto 0);
  signal place_56_succs : BooleanArray(0 downto 0);
  signal place_56_token : boolean;
  signal place_64_preds : BooleanArray(0 downto 0);
  signal place_64_succs : BooleanArray(0 downto 0);
  signal place_64_token : boolean;
  signal place_65_preds : BooleanArray(0 downto 0);
  signal place_65_succs : BooleanArray(0 downto 0);
  signal place_65_token : boolean;
  signal place_66_preds : BooleanArray(0 downto 0);
  signal place_66_succs : BooleanArray(0 downto 0);
  signal place_66_token : boolean;
  signal place_71_preds : BooleanArray(0 downto 0);
  signal place_71_succs : BooleanArray(0 downto 0);
  signal place_71_token : boolean;
  signal place_72_preds : BooleanArray(0 downto 0);
  signal place_72_succs : BooleanArray(0 downto 0);
  signal place_72_token : boolean;
  signal place_73_preds : BooleanArray(0 downto 0);
  signal place_73_succs : BooleanArray(0 downto 0);
  signal place_73_token : boolean;
  signal place_78_preds : BooleanArray(0 downto 0);
  signal place_78_succs : BooleanArray(0 downto 0);
  signal place_78_token : boolean;
  signal place_79_preds : BooleanArray(0 downto 0);
  signal place_79_succs : BooleanArray(0 downto 0);
  signal place_79_token : boolean;
  signal place_80_preds : BooleanArray(0 downto 0);
  signal place_80_succs : BooleanArray(0 downto 0);
  signal place_80_token : boolean;
  signal place_86_preds : BooleanArray(0 downto 0);
  signal place_86_succs : BooleanArray(0 downto 0);
  signal place_86_token : boolean;
  signal place_87_preds : BooleanArray(0 downto 0);
  signal place_87_succs : BooleanArray(0 downto 0);
  signal place_87_token : boolean;
  signal place_88_preds : BooleanArray(0 downto 0);
  signal place_88_succs : BooleanArray(0 downto 0);
  signal place_88_token : boolean;
  signal place_93_preds : BooleanArray(0 downto 0);
  signal place_93_succs : BooleanArray(0 downto 0);
  signal place_93_token : boolean;
  signal place_94_preds : BooleanArray(0 downto 0);
  signal place_94_succs : BooleanArray(0 downto 0);
  signal place_94_token : boolean;
  signal place_95_preds : BooleanArray(0 downto 0);
  signal place_95_succs : BooleanArray(0 downto 0);
  signal place_95_token : boolean;
  signal place_101_preds : BooleanArray(0 downto 0);
  signal place_101_succs : BooleanArray(0 downto 0);
  signal place_101_token : boolean;
  signal place_102_preds : BooleanArray(0 downto 0);
  signal place_102_succs : BooleanArray(0 downto 0);
  signal place_102_token : boolean;
  signal place_103_preds : BooleanArray(0 downto 0);
  signal place_103_succs : BooleanArray(0 downto 0);
  signal place_103_token : boolean;
  signal place_104_preds : BooleanArray(0 downto 0);
  signal place_104_succs : BooleanArray(0 downto 0);
  signal place_104_token : boolean;
  signal place_108_preds : BooleanArray(0 downto 0);
  signal place_108_succs : BooleanArray(0 downto 0);
  signal place_108_token : boolean;
  signal place_116_preds : BooleanArray(0 downto 0);
  signal place_116_succs : BooleanArray(0 downto 0);
  signal place_116_token : boolean;
  signal place_117_preds : BooleanArray(0 downto 0);
  signal place_117_succs : BooleanArray(0 downto 0);
  signal place_117_token : boolean;
  signal place_118_preds : BooleanArray(0 downto 0);
  signal place_118_succs : BooleanArray(0 downto 0);
  signal place_118_token : boolean;
  signal place_125_preds : BooleanArray(0 downto 0);
  signal place_125_succs : BooleanArray(0 downto 0);
  signal place_125_token : boolean;
  signal place_126_preds : BooleanArray(0 downto 0);
  signal place_126_succs : BooleanArray(0 downto 0);
  signal place_126_token : boolean;
  signal place_127_preds : BooleanArray(0 downto 0);
  signal place_127_succs : BooleanArray(0 downto 0);
  signal place_127_token : boolean;
  signal place_132_preds : BooleanArray(0 downto 0);
  signal place_132_succs : BooleanArray(0 downto 0);
  signal place_132_token : boolean;
  signal place_133_preds : BooleanArray(0 downto 0);
  signal place_133_succs : BooleanArray(0 downto 0);
  signal place_133_token : boolean;
  signal place_134_preds : BooleanArray(0 downto 0);
  signal place_134_succs : BooleanArray(0 downto 0);
  signal place_134_token : boolean;
  signal place_139_preds : BooleanArray(0 downto 0);
  signal place_139_succs : BooleanArray(0 downto 0);
  signal place_139_token : boolean;
  signal place_140_preds : BooleanArray(0 downto 0);
  signal place_140_succs : BooleanArray(0 downto 0);
  signal place_140_token : boolean;
  signal place_141_preds : BooleanArray(0 downto 0);
  signal place_141_succs : BooleanArray(0 downto 0);
  signal place_141_token : boolean;
  signal place_147_preds : BooleanArray(0 downto 0);
  signal place_147_succs : BooleanArray(0 downto 0);
  signal place_147_token : boolean;
  signal place_148_preds : BooleanArray(0 downto 0);
  signal place_148_succs : BooleanArray(0 downto 0);
  signal place_148_token : boolean;
  signal place_149_preds : BooleanArray(0 downto 0);
  signal place_149_succs : BooleanArray(0 downto 0);
  signal place_149_token : boolean;
  signal place_154_preds : BooleanArray(0 downto 0);
  signal place_154_succs : BooleanArray(0 downto 0);
  signal place_154_token : boolean;
  signal place_155_preds : BooleanArray(0 downto 0);
  signal place_155_succs : BooleanArray(0 downto 0);
  signal place_155_token : boolean;
  signal place_156_preds : BooleanArray(0 downto 0);
  signal place_156_succs : BooleanArray(0 downto 0);
  signal place_156_token : boolean;
  signal place_162_preds : BooleanArray(0 downto 0);
  signal place_162_succs : BooleanArray(0 downto 0);
  signal place_162_token : boolean;
  signal place_163_preds : BooleanArray(0 downto 0);
  signal place_163_succs : BooleanArray(0 downto 0);
  signal place_163_token : boolean;
  signal place_164_preds : BooleanArray(0 downto 0);
  signal place_164_succs : BooleanArray(0 downto 0);
  signal place_164_token : boolean;
  signal place_165_preds : BooleanArray(0 downto 0);
  signal place_165_succs : BooleanArray(0 downto 0);
  signal place_165_token : boolean;
  signal place_174_preds : BooleanArray(0 downto 0);
  signal place_174_succs : BooleanArray(0 downto 0);
  signal place_174_token : boolean;
  signal place_175_preds : BooleanArray(0 downto 0);
  signal place_175_succs : BooleanArray(0 downto 0);
  signal place_175_token : boolean;
  signal place_176_preds : BooleanArray(0 downto 0);
  signal place_176_succs : BooleanArray(0 downto 0);
  signal place_176_token : boolean;
  signal place_181_preds : BooleanArray(0 downto 0);
  signal place_181_succs : BooleanArray(0 downto 0);
  signal place_181_token : boolean;
  signal place_182_preds : BooleanArray(0 downto 0);
  signal place_182_succs : BooleanArray(0 downto 0);
  signal place_182_token : boolean;
  signal place_183_preds : BooleanArray(0 downto 0);
  signal place_183_succs : BooleanArray(0 downto 0);
  signal place_183_token : boolean;
  signal place_188_preds : BooleanArray(0 downto 0);
  signal place_188_succs : BooleanArray(0 downto 0);
  signal place_188_token : boolean;
  signal place_189_preds : BooleanArray(0 downto 0);
  signal place_189_succs : BooleanArray(0 downto 0);
  signal place_189_token : boolean;
  signal place_190_preds : BooleanArray(0 downto 0);
  signal place_190_succs : BooleanArray(0 downto 0);
  signal place_190_token : boolean;
  signal place_196_preds : BooleanArray(0 downto 0);
  signal place_196_succs : BooleanArray(0 downto 0);
  signal place_196_token : boolean;
  signal place_197_preds : BooleanArray(0 downto 0);
  signal place_197_succs : BooleanArray(0 downto 0);
  signal place_197_token : boolean;
  signal place_198_preds : BooleanArray(0 downto 0);
  signal place_198_succs : BooleanArray(0 downto 0);
  signal place_198_token : boolean;
  signal place_203_preds : BooleanArray(0 downto 0);
  signal place_203_succs : BooleanArray(0 downto 0);
  signal place_203_token : boolean;
  signal place_204_preds : BooleanArray(0 downto 0);
  signal place_204_succs : BooleanArray(0 downto 0);
  signal place_204_token : boolean;
  signal place_205_preds : BooleanArray(0 downto 0);
  signal place_205_succs : BooleanArray(0 downto 0);
  signal place_205_token : boolean;
  signal place_211_preds : BooleanArray(0 downto 0);
  signal place_211_succs : BooleanArray(0 downto 0);
  signal place_211_token : boolean;
  signal place_212_preds : BooleanArray(0 downto 0);
  signal place_212_succs : BooleanArray(0 downto 0);
  signal place_212_token : boolean;
  signal place_213_preds : BooleanArray(0 downto 0);
  signal place_213_succs : BooleanArray(0 downto 0);
  signal place_213_token : boolean;
  signal place_214_preds : BooleanArray(0 downto 0);
  signal place_214_succs : BooleanArray(0 downto 0);
  signal place_214_token : boolean;
  signal place_218_preds : BooleanArray(0 downto 0);
  signal place_218_succs : BooleanArray(0 downto 0);
  signal place_218_token : boolean;
  signal place_226_preds : BooleanArray(0 downto 0);
  signal place_226_succs : BooleanArray(0 downto 0);
  signal place_226_token : boolean;
  signal place_227_preds : BooleanArray(0 downto 0);
  signal place_227_succs : BooleanArray(0 downto 0);
  signal place_227_token : boolean;
  signal place_228_preds : BooleanArray(0 downto 0);
  signal place_228_succs : BooleanArray(0 downto 0);
  signal place_228_token : boolean;
  signal place_233_preds : BooleanArray(0 downto 0);
  signal place_233_succs : BooleanArray(0 downto 0);
  signal place_233_token : boolean;
  signal place_234_preds : BooleanArray(0 downto 0);
  signal place_234_succs : BooleanArray(0 downto 0);
  signal place_234_token : boolean;
  signal place_235_preds : BooleanArray(0 downto 0);
  signal place_235_succs : BooleanArray(0 downto 0);
  signal place_235_token : boolean;
  signal place_240_preds : BooleanArray(0 downto 0);
  signal place_240_succs : BooleanArray(0 downto 0);
  signal place_240_token : boolean;
  signal place_241_preds : BooleanArray(0 downto 0);
  signal place_241_succs : BooleanArray(0 downto 0);
  signal place_241_token : boolean;
  signal place_242_preds : BooleanArray(0 downto 0);
  signal place_242_succs : BooleanArray(0 downto 0);
  signal place_242_token : boolean;
  signal place_248_preds : BooleanArray(0 downto 0);
  signal place_248_succs : BooleanArray(0 downto 0);
  signal place_248_token : boolean;
  signal place_249_preds : BooleanArray(0 downto 0);
  signal place_249_succs : BooleanArray(0 downto 0);
  signal place_249_token : boolean;
  signal place_250_preds : BooleanArray(0 downto 0);
  signal place_250_succs : BooleanArray(0 downto 0);
  signal place_250_token : boolean;
  signal place_255_preds : BooleanArray(0 downto 0);
  signal place_255_succs : BooleanArray(0 downto 0);
  signal place_255_token : boolean;
  signal place_256_preds : BooleanArray(0 downto 0);
  signal place_256_succs : BooleanArray(0 downto 0);
  signal place_256_token : boolean;
  signal place_257_preds : BooleanArray(0 downto 0);
  signal place_257_succs : BooleanArray(0 downto 0);
  signal place_257_token : boolean;
  signal place_263_preds : BooleanArray(0 downto 0);
  signal place_263_succs : BooleanArray(0 downto 0);
  signal place_263_token : boolean;
  signal place_264_preds : BooleanArray(0 downto 0);
  signal place_264_succs : BooleanArray(0 downto 0);
  signal place_264_token : boolean;
  signal place_265_preds : BooleanArray(0 downto 0);
  signal place_265_succs : BooleanArray(0 downto 0);
  signal place_265_token : boolean;
  signal place_266_preds : BooleanArray(0 downto 0);
  signal place_266_succs : BooleanArray(0 downto 0);
  signal place_266_token : boolean;
  signal place_270_preds : BooleanArray(0 downto 0);
  signal place_270_succs : BooleanArray(0 downto 0);
  signal place_270_token : boolean;
  signal place_278_preds : BooleanArray(0 downto 0);
  signal place_278_succs : BooleanArray(0 downto 0);
  signal place_278_token : boolean;
  signal place_279_preds : BooleanArray(0 downto 0);
  signal place_279_succs : BooleanArray(0 downto 0);
  signal place_279_token : boolean;
  signal place_280_preds : BooleanArray(0 downto 0);
  signal place_280_succs : BooleanArray(0 downto 0);
  signal place_280_token : boolean;
  signal place_287_preds : BooleanArray(0 downto 0);
  signal place_287_succs : BooleanArray(0 downto 0);
  signal place_287_token : boolean;
  signal place_288_preds : BooleanArray(0 downto 0);
  signal place_288_succs : BooleanArray(0 downto 0);
  signal place_288_token : boolean;
  signal place_289_preds : BooleanArray(0 downto 0);
  signal place_289_succs : BooleanArray(0 downto 0);
  signal place_289_token : boolean;
  signal place_294_preds : BooleanArray(0 downto 0);
  signal place_294_succs : BooleanArray(0 downto 0);
  signal place_294_token : boolean;
  signal place_295_preds : BooleanArray(0 downto 0);
  signal place_295_succs : BooleanArray(0 downto 0);
  signal place_295_token : boolean;
  signal place_296_preds : BooleanArray(0 downto 0);
  signal place_296_succs : BooleanArray(0 downto 0);
  signal place_296_token : boolean;
  signal place_301_preds : BooleanArray(0 downto 0);
  signal place_301_succs : BooleanArray(0 downto 0);
  signal place_301_token : boolean;
  signal place_302_preds : BooleanArray(0 downto 0);
  signal place_302_succs : BooleanArray(0 downto 0);
  signal place_302_token : boolean;
  signal place_303_preds : BooleanArray(0 downto 0);
  signal place_303_succs : BooleanArray(0 downto 0);
  signal place_303_token : boolean;
  signal place_309_preds : BooleanArray(0 downto 0);
  signal place_309_succs : BooleanArray(0 downto 0);
  signal place_309_token : boolean;
  signal place_310_preds : BooleanArray(0 downto 0);
  signal place_310_succs : BooleanArray(0 downto 0);
  signal place_310_token : boolean;
  signal place_311_preds : BooleanArray(0 downto 0);
  signal place_311_succs : BooleanArray(0 downto 0);
  signal place_311_token : boolean;
  signal place_316_preds : BooleanArray(0 downto 0);
  signal place_316_succs : BooleanArray(0 downto 0);
  signal place_316_token : boolean;
  signal place_317_preds : BooleanArray(0 downto 0);
  signal place_317_succs : BooleanArray(0 downto 0);
  signal place_317_token : boolean;
  signal place_318_preds : BooleanArray(0 downto 0);
  signal place_318_succs : BooleanArray(0 downto 0);
  signal place_318_token : boolean;
  signal place_324_preds : BooleanArray(0 downto 0);
  signal place_324_succs : BooleanArray(0 downto 0);
  signal place_324_token : boolean;
  signal place_325_preds : BooleanArray(0 downto 0);
  signal place_325_succs : BooleanArray(0 downto 0);
  signal place_325_token : boolean;
  signal place_326_preds : BooleanArray(0 downto 0);
  signal place_326_succs : BooleanArray(0 downto 0);
  signal place_326_token : boolean;
  signal place_327_preds : BooleanArray(0 downto 0);
  signal place_327_succs : BooleanArray(0 downto 0);
  signal place_327_token : boolean;
  signal place_336_preds : BooleanArray(0 downto 0);
  signal place_336_succs : BooleanArray(0 downto 0);
  signal place_336_token : boolean;
  signal place_337_preds : BooleanArray(0 downto 0);
  signal place_337_succs : BooleanArray(0 downto 0);
  signal place_337_token : boolean;
  signal place_338_preds : BooleanArray(0 downto 0);
  signal place_338_succs : BooleanArray(0 downto 0);
  signal place_338_token : boolean;
  signal place_343_preds : BooleanArray(0 downto 0);
  signal place_343_succs : BooleanArray(0 downto 0);
  signal place_343_token : boolean;
  signal place_344_preds : BooleanArray(0 downto 0);
  signal place_344_succs : BooleanArray(0 downto 0);
  signal place_344_token : boolean;
  signal place_345_preds : BooleanArray(0 downto 0);
  signal place_345_succs : BooleanArray(0 downto 0);
  signal place_345_token : boolean;
  signal place_350_preds : BooleanArray(0 downto 0);
  signal place_350_succs : BooleanArray(0 downto 0);
  signal place_350_token : boolean;
  signal place_351_preds : BooleanArray(0 downto 0);
  signal place_351_succs : BooleanArray(0 downto 0);
  signal place_351_token : boolean;
  signal place_352_preds : BooleanArray(0 downto 0);
  signal place_352_succs : BooleanArray(0 downto 0);
  signal place_352_token : boolean;
  signal place_358_preds : BooleanArray(0 downto 0);
  signal place_358_succs : BooleanArray(0 downto 0);
  signal place_358_token : boolean;
  signal place_359_preds : BooleanArray(0 downto 0);
  signal place_359_succs : BooleanArray(0 downto 0);
  signal place_359_token : boolean;
  signal place_360_preds : BooleanArray(0 downto 0);
  signal place_360_succs : BooleanArray(0 downto 0);
  signal place_360_token : boolean;
  signal place_365_preds : BooleanArray(0 downto 0);
  signal place_365_succs : BooleanArray(0 downto 0);
  signal place_365_token : boolean;
  signal place_366_preds : BooleanArray(0 downto 0);
  signal place_366_succs : BooleanArray(0 downto 0);
  signal place_366_token : boolean;
  signal place_367_preds : BooleanArray(0 downto 0);
  signal place_367_succs : BooleanArray(0 downto 0);
  signal place_367_token : boolean;
  signal place_373_preds : BooleanArray(0 downto 0);
  signal place_373_succs : BooleanArray(0 downto 0);
  signal place_373_token : boolean;
  signal place_374_preds : BooleanArray(0 downto 0);
  signal place_374_succs : BooleanArray(0 downto 0);
  signal place_374_token : boolean;
  signal place_375_preds : BooleanArray(0 downto 0);
  signal place_375_succs : BooleanArray(0 downto 0);
  signal place_375_token : boolean;
  signal place_376_preds : BooleanArray(0 downto 0);
  signal place_376_succs : BooleanArray(0 downto 0);
  signal place_376_token : boolean;
  signal place_380_preds : BooleanArray(0 downto 0);
  signal place_380_succs : BooleanArray(0 downto 0);
  signal place_380_token : boolean;
  signal place_388_preds : BooleanArray(0 downto 0);
  signal place_388_succs : BooleanArray(0 downto 0);
  signal place_388_token : boolean;
  signal place_389_preds : BooleanArray(0 downto 0);
  signal place_389_succs : BooleanArray(0 downto 0);
  signal place_389_token : boolean;
  signal place_390_preds : BooleanArray(0 downto 0);
  signal place_390_succs : BooleanArray(0 downto 0);
  signal place_390_token : boolean;
  signal place_395_preds : BooleanArray(0 downto 0);
  signal place_395_succs : BooleanArray(0 downto 0);
  signal place_395_token : boolean;
  signal place_396_preds : BooleanArray(0 downto 0);
  signal place_396_succs : BooleanArray(0 downto 0);
  signal place_396_token : boolean;
  signal place_397_preds : BooleanArray(0 downto 0);
  signal place_397_succs : BooleanArray(0 downto 0);
  signal place_397_token : boolean;
  signal place_402_preds : BooleanArray(0 downto 0);
  signal place_402_succs : BooleanArray(0 downto 0);
  signal place_402_token : boolean;
  signal place_403_preds : BooleanArray(0 downto 0);
  signal place_403_succs : BooleanArray(0 downto 0);
  signal place_403_token : boolean;
  signal place_404_preds : BooleanArray(0 downto 0);
  signal place_404_succs : BooleanArray(0 downto 0);
  signal place_404_token : boolean;
  signal place_410_preds : BooleanArray(0 downto 0);
  signal place_410_succs : BooleanArray(0 downto 0);
  signal place_410_token : boolean;
  signal place_411_preds : BooleanArray(0 downto 0);
  signal place_411_succs : BooleanArray(0 downto 0);
  signal place_411_token : boolean;
  signal place_412_preds : BooleanArray(0 downto 0);
  signal place_412_succs : BooleanArray(0 downto 0);
  signal place_412_token : boolean;
  signal place_417_preds : BooleanArray(0 downto 0);
  signal place_417_succs : BooleanArray(0 downto 0);
  signal place_417_token : boolean;
  signal place_418_preds : BooleanArray(0 downto 0);
  signal place_418_succs : BooleanArray(0 downto 0);
  signal place_418_token : boolean;
  signal place_419_preds : BooleanArray(0 downto 0);
  signal place_419_succs : BooleanArray(0 downto 0);
  signal place_419_token : boolean;
  signal place_425_preds : BooleanArray(0 downto 0);
  signal place_425_succs : BooleanArray(0 downto 0);
  signal place_425_token : boolean;
  signal place_426_preds : BooleanArray(0 downto 0);
  signal place_426_succs : BooleanArray(0 downto 0);
  signal place_426_token : boolean;
  signal place_427_preds : BooleanArray(0 downto 0);
  signal place_427_succs : BooleanArray(0 downto 0);
  signal place_427_token : boolean;
  signal place_428_preds : BooleanArray(0 downto 0);
  signal place_428_succs : BooleanArray(0 downto 0);
  signal place_428_token : boolean;
  signal place_432_preds : BooleanArray(0 downto 0);
  signal place_432_succs : BooleanArray(0 downto 0);
  signal place_432_token : boolean;
  signal place_440_preds : BooleanArray(0 downto 0);
  signal place_440_succs : BooleanArray(0 downto 0);
  signal place_440_token : boolean;
  signal place_441_preds : BooleanArray(0 downto 0);
  signal place_441_succs : BooleanArray(0 downto 0);
  signal place_441_token : boolean;
  signal place_442_preds : BooleanArray(0 downto 0);
  signal place_442_succs : BooleanArray(0 downto 0);
  signal place_442_token : boolean;
  signal place_449_preds : BooleanArray(0 downto 0);
  signal place_449_succs : BooleanArray(0 downto 0);
  signal place_449_token : boolean;
  signal place_450_preds : BooleanArray(0 downto 0);
  signal place_450_succs : BooleanArray(0 downto 0);
  signal place_450_token : boolean;
  signal place_451_preds : BooleanArray(0 downto 0);
  signal place_451_succs : BooleanArray(0 downto 0);
  signal place_451_token : boolean;
  signal place_456_preds : BooleanArray(0 downto 0);
  signal place_456_succs : BooleanArray(0 downto 0);
  signal place_456_token : boolean;
  signal place_457_preds : BooleanArray(0 downto 0);
  signal place_457_succs : BooleanArray(0 downto 0);
  signal place_457_token : boolean;
  signal place_458_preds : BooleanArray(0 downto 0);
  signal place_458_succs : BooleanArray(0 downto 0);
  signal place_458_token : boolean;
  signal place_463_preds : BooleanArray(0 downto 0);
  signal place_463_succs : BooleanArray(0 downto 0);
  signal place_463_token : boolean;
  signal place_464_preds : BooleanArray(0 downto 0);
  signal place_464_succs : BooleanArray(0 downto 0);
  signal place_464_token : boolean;
  signal place_465_preds : BooleanArray(0 downto 0);
  signal place_465_succs : BooleanArray(0 downto 0);
  signal place_465_token : boolean;
  signal place_471_preds : BooleanArray(0 downto 0);
  signal place_471_succs : BooleanArray(0 downto 0);
  signal place_471_token : boolean;
  signal place_472_preds : BooleanArray(0 downto 0);
  signal place_472_succs : BooleanArray(0 downto 0);
  signal place_472_token : boolean;
  signal place_473_preds : BooleanArray(0 downto 0);
  signal place_473_succs : BooleanArray(0 downto 0);
  signal place_473_token : boolean;
  signal place_478_preds : BooleanArray(0 downto 0);
  signal place_478_succs : BooleanArray(0 downto 0);
  signal place_478_token : boolean;
  signal place_479_preds : BooleanArray(0 downto 0);
  signal place_479_succs : BooleanArray(0 downto 0);
  signal place_479_token : boolean;
  signal place_480_preds : BooleanArray(0 downto 0);
  signal place_480_succs : BooleanArray(0 downto 0);
  signal place_480_token : boolean;
  signal place_486_preds : BooleanArray(0 downto 0);
  signal place_486_succs : BooleanArray(0 downto 0);
  signal place_486_token : boolean;
  signal place_487_preds : BooleanArray(0 downto 0);
  signal place_487_succs : BooleanArray(0 downto 0);
  signal place_487_token : boolean;
  signal place_488_preds : BooleanArray(0 downto 0);
  signal place_488_succs : BooleanArray(0 downto 0);
  signal place_488_token : boolean;
  signal place_489_preds : BooleanArray(0 downto 0);
  signal place_489_succs : BooleanArray(0 downto 0);
  signal place_489_token : boolean;
  signal place_497_preds : BooleanArray(0 downto 0);
  signal place_497_succs : BooleanArray(0 downto 0);
  signal place_497_token : boolean;
  signal place_498_preds : BooleanArray(0 downto 0);
  signal place_498_succs : BooleanArray(0 downto 0);
  signal place_498_token : boolean;
  signal place_499_preds : BooleanArray(0 downto 0);
  signal place_499_succs : BooleanArray(0 downto 0);
  signal place_499_token : boolean;
  signal place_505_preds : BooleanArray(0 downto 0);
  signal place_505_succs : BooleanArray(0 downto 0);
  signal place_505_token : boolean;
  signal place_506_preds : BooleanArray(0 downto 0);
  signal place_506_succs : BooleanArray(0 downto 0);
  signal place_506_token : boolean;
  signal place_507_preds : BooleanArray(0 downto 0);
  signal place_507_succs : BooleanArray(0 downto 0);
  signal place_507_token : boolean;
  signal place_512_preds : BooleanArray(0 downto 0);
  signal place_512_succs : BooleanArray(0 downto 0);
  signal place_512_token : boolean;
  signal place_513_preds : BooleanArray(0 downto 0);
  signal place_513_succs : BooleanArray(0 downto 0);
  signal place_513_token : boolean;
  signal place_514_preds : BooleanArray(0 downto 0);
  signal place_514_succs : BooleanArray(0 downto 0);
  signal place_514_token : boolean;
  signal place_519_preds : BooleanArray(0 downto 0);
  signal place_519_succs : BooleanArray(0 downto 0);
  signal place_519_token : boolean;
  signal place_520_preds : BooleanArray(0 downto 0);
  signal place_520_succs : BooleanArray(0 downto 0);
  signal place_520_token : boolean;
  signal place_521_preds : BooleanArray(0 downto 0);
  signal place_521_succs : BooleanArray(0 downto 0);
  signal place_521_token : boolean;
  signal place_526_preds : BooleanArray(0 downto 0);
  signal place_526_succs : BooleanArray(0 downto 0);
  signal place_526_token : boolean;
  signal place_527_preds : BooleanArray(0 downto 0);
  signal place_527_succs : BooleanArray(0 downto 0);
  signal place_527_token : boolean;
  signal place_528_preds : BooleanArray(0 downto 0);
  signal place_528_succs : BooleanArray(0 downto 0);
  signal place_528_token : boolean;
  signal place_534_preds : BooleanArray(0 downto 0);
  signal place_534_succs : BooleanArray(0 downto 0);
  signal place_534_token : boolean;
  signal place_535_preds : BooleanArray(0 downto 0);
  signal place_535_succs : BooleanArray(0 downto 0);
  signal place_535_token : boolean;
  signal place_536_preds : BooleanArray(0 downto 0);
  signal place_536_succs : BooleanArray(0 downto 0);
  signal place_536_token : boolean;
  signal place_541_preds : BooleanArray(0 downto 0);
  signal place_541_succs : BooleanArray(0 downto 0);
  signal place_541_token : boolean;
  signal place_542_preds : BooleanArray(0 downto 0);
  signal place_542_succs : BooleanArray(0 downto 0);
  signal place_542_token : boolean;
  signal place_543_preds : BooleanArray(0 downto 0);
  signal place_543_succs : BooleanArray(0 downto 0);
  signal place_543_token : boolean;
  signal place_549_preds : BooleanArray(0 downto 0);
  signal place_549_succs : BooleanArray(0 downto 0);
  signal place_549_token : boolean;
  signal place_550_preds : BooleanArray(0 downto 0);
  signal place_550_succs : BooleanArray(0 downto 0);
  signal place_550_token : boolean;
  signal place_551_preds : BooleanArray(0 downto 0);
  signal place_551_succs : BooleanArray(0 downto 0);
  signal place_551_token : boolean;
  signal place_552_preds : BooleanArray(0 downto 0);
  signal place_552_succs : BooleanArray(0 downto 0);
  signal place_552_token : boolean;
  signal place_560_preds : BooleanArray(0 downto 0);
  signal place_560_succs : BooleanArray(0 downto 0);
  signal place_560_token : boolean;
  signal place_561_preds : BooleanArray(0 downto 0);
  signal place_561_succs : BooleanArray(0 downto 0);
  signal place_561_token : boolean;
  signal place_562_preds : BooleanArray(0 downto 0);
  signal place_562_succs : BooleanArray(0 downto 0);
  signal place_562_token : boolean;
  signal place_568_preds : BooleanArray(0 downto 0);
  signal place_568_succs : BooleanArray(0 downto 0);
  signal place_568_token : boolean;
  signal place_569_preds : BooleanArray(0 downto 0);
  signal place_569_succs : BooleanArray(0 downto 0);
  signal place_569_token : boolean;
  signal place_570_preds : BooleanArray(0 downto 0);
  signal place_570_succs : BooleanArray(0 downto 0);
  signal place_570_token : boolean;
  signal place_575_preds : BooleanArray(0 downto 0);
  signal place_575_succs : BooleanArray(0 downto 0);
  signal place_575_token : boolean;
  signal place_576_preds : BooleanArray(0 downto 0);
  signal place_576_succs : BooleanArray(0 downto 0);
  signal place_576_token : boolean;
  signal place_577_preds : BooleanArray(0 downto 0);
  signal place_577_succs : BooleanArray(0 downto 0);
  signal place_577_token : boolean;
  signal place_582_preds : BooleanArray(0 downto 0);
  signal place_582_succs : BooleanArray(0 downto 0);
  signal place_582_token : boolean;
  signal place_583_preds : BooleanArray(0 downto 0);
  signal place_583_succs : BooleanArray(0 downto 0);
  signal place_583_token : boolean;
  signal place_584_preds : BooleanArray(0 downto 0);
  signal place_584_succs : BooleanArray(0 downto 0);
  signal place_584_token : boolean;
  signal place_589_preds : BooleanArray(0 downto 0);
  signal place_589_succs : BooleanArray(0 downto 0);
  signal place_589_token : boolean;
  signal place_590_preds : BooleanArray(0 downto 0);
  signal place_590_succs : BooleanArray(0 downto 0);
  signal place_590_token : boolean;
  signal place_591_preds : BooleanArray(0 downto 0);
  signal place_591_succs : BooleanArray(0 downto 0);
  signal place_591_token : boolean;
  signal place_597_preds : BooleanArray(0 downto 0);
  signal place_597_succs : BooleanArray(0 downto 0);
  signal place_597_token : boolean;
  signal place_598_preds : BooleanArray(0 downto 0);
  signal place_598_succs : BooleanArray(0 downto 0);
  signal place_598_token : boolean;
  signal place_599_preds : BooleanArray(0 downto 0);
  signal place_599_succs : BooleanArray(0 downto 0);
  signal place_599_token : boolean;
  signal place_604_preds : BooleanArray(0 downto 0);
  signal place_604_succs : BooleanArray(0 downto 0);
  signal place_604_token : boolean;
  signal place_605_preds : BooleanArray(0 downto 0);
  signal place_605_succs : BooleanArray(0 downto 0);
  signal place_605_token : boolean;
  signal place_606_preds : BooleanArray(0 downto 0);
  signal place_606_succs : BooleanArray(0 downto 0);
  signal place_606_token : boolean;
  signal place_612_preds : BooleanArray(0 downto 0);
  signal place_612_succs : BooleanArray(0 downto 0);
  signal place_612_token : boolean;
  signal place_613_preds : BooleanArray(0 downto 0);
  signal place_613_succs : BooleanArray(0 downto 0);
  signal place_613_token : boolean;
  signal place_614_preds : BooleanArray(0 downto 0);
  signal place_614_succs : BooleanArray(0 downto 0);
  signal place_614_token : boolean;
  signal place_615_preds : BooleanArray(0 downto 0);
  signal place_615_succs : BooleanArray(0 downto 0);
  signal place_615_token : boolean;
  signal place_623_preds : BooleanArray(0 downto 0);
  signal place_623_succs : BooleanArray(0 downto 0);
  signal place_623_token : boolean;
  signal place_624_preds : BooleanArray(0 downto 0);
  signal place_624_succs : BooleanArray(0 downto 0);
  signal place_624_token : boolean;
  signal place_625_preds : BooleanArray(0 downto 0);
  signal place_625_succs : BooleanArray(0 downto 0);
  signal place_625_token : boolean;
  signal place_631_preds : BooleanArray(0 downto 0);
  signal place_631_succs : BooleanArray(0 downto 0);
  signal place_631_token : boolean;
  signal place_632_preds : BooleanArray(0 downto 0);
  signal place_632_succs : BooleanArray(0 downto 0);
  signal place_632_token : boolean;
  signal place_633_preds : BooleanArray(0 downto 0);
  signal place_633_succs : BooleanArray(0 downto 0);
  signal place_633_token : boolean;
  signal place_638_preds : BooleanArray(0 downto 0);
  signal place_638_succs : BooleanArray(0 downto 0);
  signal place_638_token : boolean;
  signal place_639_preds : BooleanArray(0 downto 0);
  signal place_639_succs : BooleanArray(0 downto 0);
  signal place_639_token : boolean;
  signal place_640_preds : BooleanArray(0 downto 0);
  signal place_640_succs : BooleanArray(0 downto 0);
  signal place_640_token : boolean;
  signal place_645_preds : BooleanArray(0 downto 0);
  signal place_645_succs : BooleanArray(0 downto 0);
  signal place_645_token : boolean;
  signal place_646_preds : BooleanArray(0 downto 0);
  signal place_646_succs : BooleanArray(0 downto 0);
  signal place_646_token : boolean;
  signal place_647_preds : BooleanArray(0 downto 0);
  signal place_647_succs : BooleanArray(0 downto 0);
  signal place_647_token : boolean;
  signal place_652_preds : BooleanArray(0 downto 0);
  signal place_652_succs : BooleanArray(0 downto 0);
  signal place_652_token : boolean;
  signal place_653_preds : BooleanArray(0 downto 0);
  signal place_653_succs : BooleanArray(0 downto 0);
  signal place_653_token : boolean;
  signal place_654_preds : BooleanArray(0 downto 0);
  signal place_654_succs : BooleanArray(0 downto 0);
  signal place_654_token : boolean;
  signal place_660_preds : BooleanArray(0 downto 0);
  signal place_660_succs : BooleanArray(0 downto 0);
  signal place_660_token : boolean;
  signal place_661_preds : BooleanArray(0 downto 0);
  signal place_661_succs : BooleanArray(0 downto 0);
  signal place_661_token : boolean;
  signal place_662_preds : BooleanArray(0 downto 0);
  signal place_662_succs : BooleanArray(0 downto 0);
  signal place_662_token : boolean;
  signal place_667_preds : BooleanArray(0 downto 0);
  signal place_667_succs : BooleanArray(0 downto 0);
  signal place_667_token : boolean;
  signal place_668_preds : BooleanArray(0 downto 0);
  signal place_668_succs : BooleanArray(0 downto 0);
  signal place_668_token : boolean;
  signal place_669_preds : BooleanArray(0 downto 0);
  signal place_669_succs : BooleanArray(0 downto 0);
  signal place_669_token : boolean;
  signal place_675_preds : BooleanArray(0 downto 0);
  signal place_675_succs : BooleanArray(0 downto 0);
  signal place_675_token : boolean;
  signal place_676_preds : BooleanArray(0 downto 0);
  signal place_676_succs : BooleanArray(0 downto 0);
  signal place_676_token : boolean;
  signal place_677_preds : BooleanArray(0 downto 0);
  signal place_677_succs : BooleanArray(0 downto 0);
  signal place_677_token : boolean;
  signal place_678_preds : BooleanArray(0 downto 0);
  signal place_678_succs : BooleanArray(0 downto 0);
  signal place_678_token : boolean;
  signal place_687_preds : BooleanArray(0 downto 0);
  signal place_687_succs : BooleanArray(0 downto 0);
  signal place_687_token : boolean;
  signal place_688_preds : BooleanArray(0 downto 0);
  signal place_688_succs : BooleanArray(0 downto 0);
  signal place_688_token : boolean;
  signal place_689_preds : BooleanArray(0 downto 0);
  signal place_689_succs : BooleanArray(0 downto 0);
  signal place_689_token : boolean;
  signal place_694_preds : BooleanArray(0 downto 0);
  signal place_694_succs : BooleanArray(0 downto 0);
  signal place_694_token : boolean;
  signal place_695_preds : BooleanArray(0 downto 0);
  signal place_695_succs : BooleanArray(0 downto 0);
  signal place_695_token : boolean;
  signal place_696_preds : BooleanArray(0 downto 0);
  signal place_696_succs : BooleanArray(0 downto 0);
  signal place_696_token : boolean;
  signal place_701_preds : BooleanArray(0 downto 0);
  signal place_701_succs : BooleanArray(0 downto 0);
  signal place_701_token : boolean;
  signal place_702_preds : BooleanArray(0 downto 0);
  signal place_702_succs : BooleanArray(0 downto 0);
  signal place_702_token : boolean;
  signal place_703_preds : BooleanArray(0 downto 0);
  signal place_703_succs : BooleanArray(0 downto 0);
  signal place_703_token : boolean;
  signal place_709_preds : BooleanArray(0 downto 0);
  signal place_709_succs : BooleanArray(0 downto 0);
  signal place_709_token : boolean;
  signal place_710_preds : BooleanArray(0 downto 0);
  signal place_710_succs : BooleanArray(0 downto 0);
  signal place_710_token : boolean;
  signal place_711_preds : BooleanArray(0 downto 0);
  signal place_711_succs : BooleanArray(0 downto 0);
  signal place_711_token : boolean;
  signal place_716_preds : BooleanArray(0 downto 0);
  signal place_716_succs : BooleanArray(0 downto 0);
  signal place_716_token : boolean;
  signal place_717_preds : BooleanArray(0 downto 0);
  signal place_717_succs : BooleanArray(0 downto 0);
  signal place_717_token : boolean;
  signal place_718_preds : BooleanArray(0 downto 0);
  signal place_718_succs : BooleanArray(0 downto 0);
  signal place_718_token : boolean;
  signal place_724_preds : BooleanArray(0 downto 0);
  signal place_724_succs : BooleanArray(0 downto 0);
  signal place_724_token : boolean;
  signal place_725_preds : BooleanArray(0 downto 0);
  signal place_725_succs : BooleanArray(0 downto 0);
  signal place_725_token : boolean;
  signal place_726_preds : BooleanArray(0 downto 0);
  signal place_726_succs : BooleanArray(0 downto 0);
  signal place_726_token : boolean;
  signal place_727_preds : BooleanArray(0 downto 0);
  signal place_727_succs : BooleanArray(0 downto 0);
  signal place_727_token : boolean;
  signal place_731_preds : BooleanArray(0 downto 0);
  signal place_731_succs : BooleanArray(0 downto 0);
  signal place_731_token : boolean;
  signal place_738_preds : BooleanArray(0 downto 0);
  signal place_738_succs : BooleanArray(0 downto 0);
  signal place_738_token : boolean;
  signal place_739_preds : BooleanArray(0 downto 0);
  signal place_739_succs : BooleanArray(0 downto 0);
  signal place_739_token : boolean;
  signal place_740_preds : BooleanArray(0 downto 0);
  signal place_740_succs : BooleanArray(0 downto 0);
  signal place_740_token : boolean;
  signal place_745_preds : BooleanArray(0 downto 0);
  signal place_745_succs : BooleanArray(0 downto 0);
  signal place_745_token : boolean;
  signal place_746_preds : BooleanArray(0 downto 0);
  signal place_746_succs : BooleanArray(0 downto 0);
  signal place_746_token : boolean;
  signal place_747_preds : BooleanArray(0 downto 0);
  signal place_747_succs : BooleanArray(0 downto 0);
  signal place_747_token : boolean;
  signal place_752_preds : BooleanArray(0 downto 0);
  signal place_752_succs : BooleanArray(0 downto 0);
  signal place_752_token : boolean;
  signal place_753_preds : BooleanArray(0 downto 0);
  signal place_753_succs : BooleanArray(0 downto 0);
  signal place_753_token : boolean;
  signal place_754_preds : BooleanArray(0 downto 0);
  signal place_754_succs : BooleanArray(0 downto 0);
  signal place_754_token : boolean;
  signal place_760_preds : BooleanArray(0 downto 0);
  signal place_760_succs : BooleanArray(0 downto 0);
  signal place_760_token : boolean;
  signal place_761_preds : BooleanArray(0 downto 0);
  signal place_761_succs : BooleanArray(0 downto 0);
  signal place_761_token : boolean;
  signal place_762_preds : BooleanArray(0 downto 0);
  signal place_762_succs : BooleanArray(0 downto 0);
  signal place_762_token : boolean;
  signal place_767_preds : BooleanArray(0 downto 0);
  signal place_767_succs : BooleanArray(0 downto 0);
  signal place_767_token : boolean;
  signal place_768_preds : BooleanArray(0 downto 0);
  signal place_768_succs : BooleanArray(0 downto 0);
  signal place_768_token : boolean;
  signal place_769_preds : BooleanArray(0 downto 0);
  signal place_769_succs : BooleanArray(0 downto 0);
  signal place_769_token : boolean;
  signal place_775_preds : BooleanArray(0 downto 0);
  signal place_775_succs : BooleanArray(0 downto 0);
  signal place_775_token : boolean;
  signal place_776_preds : BooleanArray(0 downto 0);
  signal place_776_succs : BooleanArray(0 downto 0);
  signal place_776_token : boolean;
  signal place_777_preds : BooleanArray(0 downto 0);
  signal place_777_succs : BooleanArray(0 downto 0);
  signal place_777_token : boolean;
  signal place_778_preds : BooleanArray(0 downto 0);
  signal place_778_succs : BooleanArray(0 downto 0);
  signal place_778_token : boolean;
  signal place_782_preds : BooleanArray(0 downto 0);
  signal place_782_succs : BooleanArray(0 downto 0);
  signal place_782_token : boolean;
  signal place_789_preds : BooleanArray(0 downto 0);
  signal place_789_succs : BooleanArray(0 downto 0);
  signal place_789_token : boolean;
  signal place_790_preds : BooleanArray(0 downto 0);
  signal place_790_succs : BooleanArray(0 downto 0);
  signal place_790_token : boolean;
  signal place_791_preds : BooleanArray(0 downto 0);
  signal place_791_succs : BooleanArray(0 downto 0);
  signal place_791_token : boolean;
  signal place_797_preds : BooleanArray(0 downto 0);
  signal place_797_succs : BooleanArray(0 downto 0);
  signal place_797_token : boolean;
  signal place_798_preds : BooleanArray(0 downto 0);
  signal place_798_succs : BooleanArray(0 downto 0);
  signal place_798_token : boolean;
  signal place_799_preds : BooleanArray(0 downto 0);
  signal place_799_succs : BooleanArray(0 downto 0);
  signal place_799_token : boolean;
  signal place_804_preds : BooleanArray(0 downto 0);
  signal place_804_succs : BooleanArray(0 downto 0);
  signal place_804_token : boolean;
  signal place_805_preds : BooleanArray(0 downto 0);
  signal place_805_succs : BooleanArray(0 downto 0);
  signal place_805_token : boolean;
  signal place_806_preds : BooleanArray(0 downto 0);
  signal place_806_succs : BooleanArray(0 downto 0);
  signal place_806_token : boolean;
  signal place_811_preds : BooleanArray(0 downto 0);
  signal place_811_succs : BooleanArray(0 downto 0);
  signal place_811_token : boolean;
  signal place_812_preds : BooleanArray(0 downto 0);
  signal place_812_succs : BooleanArray(0 downto 0);
  signal place_812_token : boolean;
  signal place_813_preds : BooleanArray(0 downto 0);
  signal place_813_succs : BooleanArray(0 downto 0);
  signal place_813_token : boolean;
  signal place_818_preds : BooleanArray(0 downto 0);
  signal place_818_succs : BooleanArray(0 downto 0);
  signal place_818_token : boolean;
  signal place_819_preds : BooleanArray(0 downto 0);
  signal place_819_succs : BooleanArray(0 downto 0);
  signal place_819_token : boolean;
  signal place_820_preds : BooleanArray(0 downto 0);
  signal place_820_succs : BooleanArray(0 downto 0);
  signal place_820_token : boolean;
  signal place_826_preds : BooleanArray(0 downto 0);
  signal place_826_succs : BooleanArray(0 downto 0);
  signal place_826_token : boolean;
  signal place_827_preds : BooleanArray(0 downto 0);
  signal place_827_succs : BooleanArray(0 downto 0);
  signal place_827_token : boolean;
  signal place_828_preds : BooleanArray(0 downto 0);
  signal place_828_succs : BooleanArray(0 downto 0);
  signal place_828_token : boolean;
  signal place_833_preds : BooleanArray(0 downto 0);
  signal place_833_succs : BooleanArray(0 downto 0);
  signal place_833_token : boolean;
  signal place_834_preds : BooleanArray(0 downto 0);
  signal place_834_succs : BooleanArray(0 downto 0);
  signal place_834_token : boolean;
  signal place_835_preds : BooleanArray(0 downto 0);
  signal place_835_succs : BooleanArray(0 downto 0);
  signal place_835_token : boolean;
  signal place_841_preds : BooleanArray(0 downto 0);
  signal place_841_succs : BooleanArray(0 downto 0);
  signal place_841_token : boolean;
  signal place_842_preds : BooleanArray(0 downto 0);
  signal place_842_succs : BooleanArray(0 downto 0);
  signal place_842_token : boolean;
  signal place_843_preds : BooleanArray(0 downto 0);
  signal place_843_succs : BooleanArray(0 downto 0);
  signal place_843_token : boolean;
  signal place_844_preds : BooleanArray(0 downto 0);
  signal place_844_succs : BooleanArray(0 downto 0);
  signal place_844_token : boolean;
  signal place_853_preds : BooleanArray(0 downto 0);
  signal place_853_succs : BooleanArray(0 downto 0);
  signal place_853_token : boolean;
  signal place_854_preds : BooleanArray(0 downto 0);
  signal place_854_succs : BooleanArray(0 downto 0);
  signal place_854_token : boolean;
  signal place_855_preds : BooleanArray(0 downto 0);
  signal place_855_succs : BooleanArray(0 downto 0);
  signal place_855_token : boolean;
  signal place_860_preds : BooleanArray(0 downto 0);
  signal place_860_succs : BooleanArray(0 downto 0);
  signal place_860_token : boolean;
  signal place_861_preds : BooleanArray(0 downto 0);
  signal place_861_succs : BooleanArray(0 downto 0);
  signal place_861_token : boolean;
  signal place_862_preds : BooleanArray(0 downto 0);
  signal place_862_succs : BooleanArray(0 downto 0);
  signal place_862_token : boolean;
  signal place_867_preds : BooleanArray(0 downto 0);
  signal place_867_succs : BooleanArray(0 downto 0);
  signal place_867_token : boolean;
  signal place_868_preds : BooleanArray(0 downto 0);
  signal place_868_succs : BooleanArray(0 downto 0);
  signal place_868_token : boolean;
  signal place_869_preds : BooleanArray(0 downto 0);
  signal place_869_succs : BooleanArray(0 downto 0);
  signal place_869_token : boolean;
  signal place_875_preds : BooleanArray(0 downto 0);
  signal place_875_succs : BooleanArray(0 downto 0);
  signal place_875_token : boolean;
  signal place_876_preds : BooleanArray(0 downto 0);
  signal place_876_succs : BooleanArray(0 downto 0);
  signal place_876_token : boolean;
  signal place_877_preds : BooleanArray(0 downto 0);
  signal place_877_succs : BooleanArray(0 downto 0);
  signal place_877_token : boolean;
  signal place_882_preds : BooleanArray(0 downto 0);
  signal place_882_succs : BooleanArray(0 downto 0);
  signal place_882_token : boolean;
  signal place_883_preds : BooleanArray(0 downto 0);
  signal place_883_succs : BooleanArray(0 downto 0);
  signal place_883_token : boolean;
  signal place_884_preds : BooleanArray(0 downto 0);
  signal place_884_succs : BooleanArray(0 downto 0);
  signal place_884_token : boolean;
  signal place_890_preds : BooleanArray(0 downto 0);
  signal place_890_succs : BooleanArray(0 downto 0);
  signal place_890_token : boolean;
  signal place_891_preds : BooleanArray(0 downto 0);
  signal place_891_succs : BooleanArray(0 downto 0);
  signal place_891_token : boolean;
  signal place_892_preds : BooleanArray(0 downto 0);
  signal place_892_succs : BooleanArray(0 downto 0);
  signal place_892_token : boolean;
  signal place_893_preds : BooleanArray(0 downto 0);
  signal place_893_succs : BooleanArray(0 downto 0);
  signal place_893_token : boolean;
  signal place_897_preds : BooleanArray(0 downto 0);
  signal place_897_succs : BooleanArray(0 downto 0);
  signal place_897_token : boolean;
  signal place_904_preds : BooleanArray(0 downto 0);
  signal place_904_succs : BooleanArray(0 downto 0);
  signal place_904_token : boolean;
  signal place_905_preds : BooleanArray(0 downto 0);
  signal place_905_succs : BooleanArray(0 downto 0);
  signal place_905_token : boolean;
  signal place_906_preds : BooleanArray(0 downto 0);
  signal place_906_succs : BooleanArray(0 downto 0);
  signal place_906_token : boolean;
  signal place_911_preds : BooleanArray(0 downto 0);
  signal place_911_succs : BooleanArray(0 downto 0);
  signal place_911_token : boolean;
  signal place_912_preds : BooleanArray(0 downto 0);
  signal place_912_succs : BooleanArray(0 downto 0);
  signal place_912_token : boolean;
  signal place_913_preds : BooleanArray(0 downto 0);
  signal place_913_succs : BooleanArray(0 downto 0);
  signal place_913_token : boolean;
  signal place_918_preds : BooleanArray(0 downto 0);
  signal place_918_succs : BooleanArray(0 downto 0);
  signal place_918_token : boolean;
  signal place_919_preds : BooleanArray(0 downto 0);
  signal place_919_succs : BooleanArray(0 downto 0);
  signal place_919_token : boolean;
  signal place_920_preds : BooleanArray(0 downto 0);
  signal place_920_succs : BooleanArray(0 downto 0);
  signal place_920_token : boolean;
  signal place_926_preds : BooleanArray(0 downto 0);
  signal place_926_succs : BooleanArray(0 downto 0);
  signal place_926_token : boolean;
  signal place_927_preds : BooleanArray(0 downto 0);
  signal place_927_succs : BooleanArray(0 downto 0);
  signal place_927_token : boolean;
  signal place_928_preds : BooleanArray(0 downto 0);
  signal place_928_succs : BooleanArray(0 downto 0);
  signal place_928_token : boolean;
  signal place_933_preds : BooleanArray(0 downto 0);
  signal place_933_succs : BooleanArray(0 downto 0);
  signal place_933_token : boolean;
  signal place_934_preds : BooleanArray(0 downto 0);
  signal place_934_succs : BooleanArray(0 downto 0);
  signal place_934_token : boolean;
  signal place_935_preds : BooleanArray(0 downto 0);
  signal place_935_succs : BooleanArray(0 downto 0);
  signal place_935_token : boolean;
  signal place_941_preds : BooleanArray(0 downto 0);
  signal place_941_succs : BooleanArray(0 downto 0);
  signal place_941_token : boolean;
  signal place_942_preds : BooleanArray(0 downto 0);
  signal place_942_succs : BooleanArray(0 downto 0);
  signal place_942_token : boolean;
  signal place_943_preds : BooleanArray(0 downto 0);
  signal place_943_succs : BooleanArray(0 downto 0);
  signal place_943_token : boolean;
  signal place_944_preds : BooleanArray(0 downto 0);
  signal place_944_succs : BooleanArray(0 downto 0);
  signal place_944_token : boolean;
  signal place_948_preds : BooleanArray(0 downto 0);
  signal place_948_succs : BooleanArray(0 downto 0);
  signal place_948_token : boolean;
  signal place_955_preds : BooleanArray(0 downto 0);
  signal place_955_succs : BooleanArray(0 downto 0);
  signal place_955_token : boolean;
  signal place_956_preds : BooleanArray(0 downto 0);
  signal place_956_succs : BooleanArray(0 downto 0);
  signal place_956_token : boolean;
  signal place_957_preds : BooleanArray(0 downto 0);
  signal place_957_succs : BooleanArray(0 downto 0);
  signal place_957_token : boolean;
  signal place_963_preds : BooleanArray(0 downto 0);
  signal place_963_succs : BooleanArray(0 downto 0);
  signal place_963_token : boolean;
  signal place_964_preds : BooleanArray(0 downto 0);
  signal place_964_succs : BooleanArray(0 downto 0);
  signal place_964_token : boolean;
  signal place_965_preds : BooleanArray(0 downto 0);
  signal place_965_succs : BooleanArray(0 downto 0);
  signal place_965_token : boolean;
  signal place_970_preds : BooleanArray(0 downto 0);
  signal place_970_succs : BooleanArray(0 downto 0);
  signal place_970_token : boolean;
  signal place_971_preds : BooleanArray(0 downto 0);
  signal place_971_succs : BooleanArray(0 downto 0);
  signal place_971_token : boolean;
  signal place_972_preds : BooleanArray(0 downto 0);
  signal place_972_succs : BooleanArray(0 downto 0);
  signal place_972_token : boolean;
  signal place_977_preds : BooleanArray(0 downto 0);
  signal place_977_succs : BooleanArray(0 downto 0);
  signal place_977_token : boolean;
  signal place_978_preds : BooleanArray(0 downto 0);
  signal place_978_succs : BooleanArray(0 downto 0);
  signal place_978_token : boolean;
  signal place_979_preds : BooleanArray(0 downto 0);
  signal place_979_succs : BooleanArray(0 downto 0);
  signal place_979_token : boolean;
  signal place_984_preds : BooleanArray(0 downto 0);
  signal place_984_succs : BooleanArray(0 downto 0);
  signal place_984_token : boolean;
  signal place_985_preds : BooleanArray(0 downto 0);
  signal place_985_succs : BooleanArray(0 downto 0);
  signal place_985_token : boolean;
  signal place_986_preds : BooleanArray(0 downto 0);
  signal place_986_succs : BooleanArray(0 downto 0);
  signal place_986_token : boolean;
  signal place_992_preds : BooleanArray(0 downto 0);
  signal place_992_succs : BooleanArray(0 downto 0);
  signal place_992_token : boolean;
  signal place_993_preds : BooleanArray(0 downto 0);
  signal place_993_succs : BooleanArray(0 downto 0);
  signal place_993_token : boolean;
  signal place_994_preds : BooleanArray(0 downto 0);
  signal place_994_succs : BooleanArray(0 downto 0);
  signal place_994_token : boolean;
  signal place_999_preds : BooleanArray(0 downto 0);
  signal place_999_succs : BooleanArray(0 downto 0);
  signal place_999_token : boolean;
  signal place_1000_preds : BooleanArray(0 downto 0);
  signal place_1000_succs : BooleanArray(0 downto 0);
  signal place_1000_token : boolean;
  signal place_1001_preds : BooleanArray(0 downto 0);
  signal place_1001_succs : BooleanArray(0 downto 0);
  signal place_1001_token : boolean;
  signal place_1007_preds : BooleanArray(0 downto 0);
  signal place_1007_succs : BooleanArray(0 downto 0);
  signal place_1007_token : boolean;
  signal place_1008_preds : BooleanArray(0 downto 0);
  signal place_1008_succs : BooleanArray(0 downto 0);
  signal place_1008_token : boolean;
  signal place_1009_preds : BooleanArray(0 downto 0);
  signal place_1009_succs : BooleanArray(0 downto 0);
  signal place_1009_token : boolean;
  signal place_1010_preds : BooleanArray(0 downto 0);
  signal place_1010_succs : BooleanArray(0 downto 0);
  signal place_1010_token : boolean;
  signal place_1019_preds : BooleanArray(0 downto 0);
  signal place_1019_succs : BooleanArray(0 downto 0);
  signal place_1019_token : boolean;
  signal place_1020_preds : BooleanArray(0 downto 0);
  signal place_1020_succs : BooleanArray(0 downto 0);
  signal place_1020_token : boolean;
  signal place_1021_preds : BooleanArray(0 downto 0);
  signal place_1021_succs : BooleanArray(0 downto 0);
  signal place_1021_token : boolean;
  signal place_1026_preds : BooleanArray(0 downto 0);
  signal place_1026_succs : BooleanArray(0 downto 0);
  signal place_1026_token : boolean;
  signal place_1027_preds : BooleanArray(0 downto 0);
  signal place_1027_succs : BooleanArray(0 downto 0);
  signal place_1027_token : boolean;
  signal place_1028_preds : BooleanArray(0 downto 0);
  signal place_1028_succs : BooleanArray(0 downto 0);
  signal place_1028_token : boolean;
  signal place_1033_preds : BooleanArray(0 downto 0);
  signal place_1033_succs : BooleanArray(0 downto 0);
  signal place_1033_token : boolean;
  signal place_1034_preds : BooleanArray(0 downto 0);
  signal place_1034_succs : BooleanArray(0 downto 0);
  signal place_1034_token : boolean;
  signal place_1035_preds : BooleanArray(0 downto 0);
  signal place_1035_succs : BooleanArray(0 downto 0);
  signal place_1035_token : boolean;
  signal place_1041_preds : BooleanArray(0 downto 0);
  signal place_1041_succs : BooleanArray(0 downto 0);
  signal place_1041_token : boolean;
  signal place_1042_preds : BooleanArray(0 downto 0);
  signal place_1042_succs : BooleanArray(0 downto 0);
  signal place_1042_token : boolean;
  signal place_1043_preds : BooleanArray(0 downto 0);
  signal place_1043_succs : BooleanArray(0 downto 0);
  signal place_1043_token : boolean;
  signal place_1048_preds : BooleanArray(0 downto 0);
  signal place_1048_succs : BooleanArray(0 downto 0);
  signal place_1048_token : boolean;
  signal place_1049_preds : BooleanArray(0 downto 0);
  signal place_1049_succs : BooleanArray(0 downto 0);
  signal place_1049_token : boolean;
  signal place_1050_preds : BooleanArray(0 downto 0);
  signal place_1050_succs : BooleanArray(0 downto 0);
  signal place_1050_token : boolean;
  signal place_1056_preds : BooleanArray(0 downto 0);
  signal place_1056_succs : BooleanArray(0 downto 0);
  signal place_1056_token : boolean;
  signal place_1057_preds : BooleanArray(0 downto 0);
  signal place_1057_succs : BooleanArray(0 downto 0);
  signal place_1057_token : boolean;
  signal place_1058_preds : BooleanArray(0 downto 0);
  signal place_1058_succs : BooleanArray(0 downto 0);
  signal place_1058_token : boolean;
  signal place_1059_preds : BooleanArray(0 downto 0);
  signal place_1059_succs : BooleanArray(0 downto 0);
  signal place_1059_token : boolean;
  signal place_1063_preds : BooleanArray(0 downto 0);
  signal place_1063_succs : BooleanArray(0 downto 0);
  signal place_1063_token : boolean;
  signal place_1070_preds : BooleanArray(0 downto 0);
  signal place_1070_succs : BooleanArray(0 downto 0);
  signal place_1070_token : boolean;
  signal place_1071_preds : BooleanArray(0 downto 0);
  signal place_1071_succs : BooleanArray(0 downto 0);
  signal place_1071_token : boolean;
  signal place_1072_preds : BooleanArray(0 downto 0);
  signal place_1072_succs : BooleanArray(0 downto 0);
  signal place_1072_token : boolean;
  signal place_1077_preds : BooleanArray(0 downto 0);
  signal place_1077_succs : BooleanArray(0 downto 0);
  signal place_1077_token : boolean;
  signal place_1078_preds : BooleanArray(0 downto 0);
  signal place_1078_succs : BooleanArray(0 downto 0);
  signal place_1078_token : boolean;
  signal place_1079_preds : BooleanArray(0 downto 0);
  signal place_1079_succs : BooleanArray(0 downto 0);
  signal place_1079_token : boolean;
  signal place_1084_preds : BooleanArray(0 downto 0);
  signal place_1084_succs : BooleanArray(0 downto 0);
  signal place_1084_token : boolean;
  signal place_1085_preds : BooleanArray(0 downto 0);
  signal place_1085_succs : BooleanArray(0 downto 0);
  signal place_1085_token : boolean;
  signal place_1086_preds : BooleanArray(0 downto 0);
  signal place_1086_succs : BooleanArray(0 downto 0);
  signal place_1086_token : boolean;
  signal place_1092_preds : BooleanArray(0 downto 0);
  signal place_1092_succs : BooleanArray(0 downto 0);
  signal place_1092_token : boolean;
  signal place_1093_preds : BooleanArray(0 downto 0);
  signal place_1093_succs : BooleanArray(0 downto 0);
  signal place_1093_token : boolean;
  signal place_1094_preds : BooleanArray(0 downto 0);
  signal place_1094_succs : BooleanArray(0 downto 0);
  signal place_1094_token : boolean;
  signal place_1099_preds : BooleanArray(0 downto 0);
  signal place_1099_succs : BooleanArray(0 downto 0);
  signal place_1099_token : boolean;
  signal place_1100_preds : BooleanArray(0 downto 0);
  signal place_1100_succs : BooleanArray(0 downto 0);
  signal place_1100_token : boolean;
  signal place_1101_preds : BooleanArray(0 downto 0);
  signal place_1101_succs : BooleanArray(0 downto 0);
  signal place_1101_token : boolean;
  signal place_1107_preds : BooleanArray(0 downto 0);
  signal place_1107_succs : BooleanArray(0 downto 0);
  signal place_1107_token : boolean;
  signal place_1108_preds : BooleanArray(0 downto 0);
  signal place_1108_succs : BooleanArray(0 downto 0);
  signal place_1108_token : boolean;
  signal place_1109_preds : BooleanArray(0 downto 0);
  signal place_1109_succs : BooleanArray(0 downto 0);
  signal place_1109_token : boolean;
  signal place_1110_preds : BooleanArray(0 downto 0);
  signal place_1110_succs : BooleanArray(0 downto 0);
  signal place_1110_token : boolean;
  signal place_1114_preds : BooleanArray(0 downto 0);
  signal place_1114_succs : BooleanArray(0 downto 0);
  signal place_1114_token : boolean;
  signal place_1121_preds : BooleanArray(0 downto 0);
  signal place_1121_succs : BooleanArray(0 downto 0);
  signal place_1121_token : boolean;
  signal place_1122_preds : BooleanArray(0 downto 0);
  signal place_1122_succs : BooleanArray(0 downto 0);
  signal place_1122_token : boolean;
  signal place_1123_preds : BooleanArray(0 downto 0);
  signal place_1123_succs : BooleanArray(0 downto 0);
  signal place_1123_token : boolean;
  signal place_1129_preds : BooleanArray(0 downto 0);
  signal place_1129_succs : BooleanArray(0 downto 0);
  signal place_1129_token : boolean;
  signal place_1130_preds : BooleanArray(0 downto 0);
  signal place_1130_succs : BooleanArray(0 downto 0);
  signal place_1130_token : boolean;
  signal place_1131_preds : BooleanArray(0 downto 0);
  signal place_1131_succs : BooleanArray(0 downto 0);
  signal place_1131_token : boolean;
  signal place_1136_preds : BooleanArray(0 downto 0);
  signal place_1136_succs : BooleanArray(0 downto 0);
  signal place_1136_token : boolean;
  signal place_1137_preds : BooleanArray(0 downto 0);
  signal place_1137_succs : BooleanArray(0 downto 0);
  signal place_1137_token : boolean;
  signal place_1138_preds : BooleanArray(0 downto 0);
  signal place_1138_succs : BooleanArray(0 downto 0);
  signal place_1138_token : boolean;
  signal place_1143_preds : BooleanArray(0 downto 0);
  signal place_1143_succs : BooleanArray(0 downto 0);
  signal place_1143_token : boolean;
  signal place_1144_preds : BooleanArray(0 downto 0);
  signal place_1144_succs : BooleanArray(0 downto 0);
  signal place_1144_token : boolean;
  signal place_1145_preds : BooleanArray(0 downto 0);
  signal place_1145_succs : BooleanArray(0 downto 0);
  signal place_1145_token : boolean;
  signal place_1150_preds : BooleanArray(0 downto 0);
  signal place_1150_succs : BooleanArray(0 downto 0);
  signal place_1150_token : boolean;
  signal place_1151_preds : BooleanArray(0 downto 0);
  signal place_1151_succs : BooleanArray(0 downto 0);
  signal place_1151_token : boolean;
  signal place_1152_preds : BooleanArray(0 downto 0);
  signal place_1152_succs : BooleanArray(0 downto 0);
  signal place_1152_token : boolean;
  signal place_1158_preds : BooleanArray(0 downto 0);
  signal place_1158_succs : BooleanArray(0 downto 0);
  signal place_1158_token : boolean;
  signal place_1159_preds : BooleanArray(0 downto 0);
  signal place_1159_succs : BooleanArray(0 downto 0);
  signal place_1159_token : boolean;
  signal place_1160_preds : BooleanArray(0 downto 0);
  signal place_1160_succs : BooleanArray(0 downto 0);
  signal place_1160_token : boolean;
  signal place_1165_preds : BooleanArray(0 downto 0);
  signal place_1165_succs : BooleanArray(0 downto 0);
  signal place_1165_token : boolean;
  signal place_1166_preds : BooleanArray(0 downto 0);
  signal place_1166_succs : BooleanArray(0 downto 0);
  signal place_1166_token : boolean;
  signal place_1167_preds : BooleanArray(0 downto 0);
  signal place_1167_succs : BooleanArray(0 downto 0);
  signal place_1167_token : boolean;
  signal place_1173_preds : BooleanArray(0 downto 0);
  signal place_1173_succs : BooleanArray(0 downto 0);
  signal place_1173_token : boolean;
  signal place_1174_preds : BooleanArray(0 downto 0);
  signal place_1174_succs : BooleanArray(0 downto 0);
  signal place_1174_token : boolean;
  signal place_1175_preds : BooleanArray(0 downto 0);
  signal place_1175_succs : BooleanArray(0 downto 0);
  signal place_1175_token : boolean;
  signal place_1176_preds : BooleanArray(0 downto 0);
  signal place_1176_succs : BooleanArray(0 downto 0);
  signal place_1176_token : boolean;
  signal place_1184_preds : BooleanArray(0 downto 0);
  signal place_1184_succs : BooleanArray(0 downto 0);
  signal place_1184_token : boolean;
  signal place_1185_preds : BooleanArray(0 downto 0);
  signal place_1185_succs : BooleanArray(0 downto 0);
  signal place_1185_token : boolean;
  signal place_1186_preds : BooleanArray(0 downto 0);
  signal place_1186_succs : BooleanArray(0 downto 0);
  signal place_1186_token : boolean;
  signal place_1192_preds : BooleanArray(0 downto 0);
  signal place_1192_succs : BooleanArray(0 downto 0);
  signal place_1192_token : boolean;
  signal place_1193_preds : BooleanArray(0 downto 0);
  signal place_1193_succs : BooleanArray(0 downto 0);
  signal place_1193_token : boolean;
  signal place_1194_preds : BooleanArray(0 downto 0);
  signal place_1194_succs : BooleanArray(0 downto 0);
  signal place_1194_token : boolean;
  signal place_1200_preds : BooleanArray(0 downto 0);
  signal place_1200_succs : BooleanArray(0 downto 0);
  signal place_1200_token : boolean;
  signal place_1201_preds : BooleanArray(0 downto 0);
  signal place_1201_succs : BooleanArray(0 downto 0);
  signal place_1201_token : boolean;
  signal place_1202_preds : BooleanArray(0 downto 0);
  signal place_1202_succs : BooleanArray(0 downto 0);
  signal place_1202_token : boolean;
  signal place_1203_preds : BooleanArray(0 downto 0);
  signal place_1203_succs : BooleanArray(0 downto 0);
  signal place_1203_token : boolean;
  signal place_1206_preds : BooleanArray(0 downto 0);
  signal place_1206_succs : BooleanArray(0 downto 0);
  signal place_1206_token : boolean;
  signal place_1207_preds : BooleanArray(0 downto 0);
  signal place_1207_succs : BooleanArray(0 downto 0);
  signal place_1207_token : boolean;
  signal place_1208_preds : BooleanArray(0 downto 0);
  signal place_1208_succs : BooleanArray(0 downto 0);
  signal place_1208_token : boolean;
  signal place_1209_preds : BooleanArray(0 downto 0);
  signal place_1209_succs : BooleanArray(0 downto 0);
  signal place_1209_token : boolean;
  signal place_1210_preds : BooleanArray(0 downto 0);
  signal place_1210_succs : BooleanArray(0 downto 0);
  signal place_1210_token : boolean;
  signal place_1211_preds : BooleanArray(0 downto 0);
  signal place_1211_succs : BooleanArray(0 downto 0);
  signal place_1211_token : boolean;
  signal place_1212_preds : BooleanArray(0 downto 0);
  signal place_1212_succs : BooleanArray(0 downto 0);
  signal place_1212_token : boolean;
  signal place_1213_preds : BooleanArray(0 downto 0);
  signal place_1213_succs : BooleanArray(0 downto 0);
  signal place_1213_token : boolean;
  signal place_1214_preds : BooleanArray(0 downto 0);
  signal place_1214_succs : BooleanArray(0 downto 0);
  signal place_1214_token : boolean;
  signal place_1215_preds : BooleanArray(0 downto 0);
  signal place_1215_succs : BooleanArray(0 downto 0);
  signal place_1215_token : boolean;
  signal place_1216_preds : BooleanArray(0 downto 0);
  signal place_1216_succs : BooleanArray(0 downto 0);
  signal place_1216_token : boolean;
  signal place_1217_preds : BooleanArray(0 downto 0);
  signal place_1217_succs : BooleanArray(0 downto 0);
  signal place_1217_token : boolean;
  signal place_1218_preds : BooleanArray(0 downto 0);
  signal place_1218_succs : BooleanArray(0 downto 0);
  signal place_1218_token : boolean;
  signal place_1219_preds : BooleanArray(0 downto 0);
  signal place_1219_succs : BooleanArray(0 downto 0);
  signal place_1219_token : boolean;
  signal place_1220_preds : BooleanArray(0 downto 0);
  signal place_1220_succs : BooleanArray(0 downto 0);
  signal place_1220_token : boolean;
  signal place_1221_preds : BooleanArray(0 downto 0);
  signal place_1221_succs : BooleanArray(0 downto 0);
  signal place_1221_token : boolean;
  signal place_1222_preds : BooleanArray(0 downto 0);
  signal place_1222_succs : BooleanArray(0 downto 0);
  signal place_1222_token : boolean;
  signal place_1223_preds : BooleanArray(0 downto 0);
  signal place_1223_succs : BooleanArray(0 downto 0);
  signal place_1223_token : boolean;
  signal place_1224_preds : BooleanArray(0 downto 0);
  signal place_1224_succs : BooleanArray(0 downto 0);
  signal place_1224_token : boolean;
  signal place_1225_preds : BooleanArray(0 downto 0);
  signal place_1225_succs : BooleanArray(0 downto 0);
  signal place_1225_token : boolean;
  signal place_1226_preds : BooleanArray(0 downto 0);
  signal place_1226_succs : BooleanArray(0 downto 0);
  signal place_1226_token : boolean;
  signal place_1227_preds : BooleanArray(0 downto 0);
  signal place_1227_succs : BooleanArray(0 downto 0);
  signal place_1227_token : boolean;
  signal place_1228_preds : BooleanArray(0 downto 0);
  signal place_1228_succs : BooleanArray(0 downto 0);
  signal place_1228_token : boolean;
  signal place_1229_preds : BooleanArray(0 downto 0);
  signal place_1229_succs : BooleanArray(0 downto 0);
  signal place_1229_token : boolean;
  signal place_1230_preds : BooleanArray(0 downto 0);
  signal place_1230_succs : BooleanArray(0 downto 0);
  signal place_1230_token : boolean;
  signal place_1231_preds : BooleanArray(0 downto 0);
  signal place_1231_succs : BooleanArray(0 downto 0);
  signal place_1231_token : boolean;
  signal place_1232_preds : BooleanArray(0 downto 0);
  signal place_1232_succs : BooleanArray(0 downto 0);
  signal place_1232_token : boolean;
  signal place_1233_preds : BooleanArray(0 downto 0);
  signal place_1233_succs : BooleanArray(0 downto 0);
  signal place_1233_token : boolean;
  signal place_1234_preds : BooleanArray(0 downto 0);
  signal place_1234_succs : BooleanArray(0 downto 0);
  signal place_1234_token : boolean;
  signal place_1235_preds : BooleanArray(0 downto 0);
  signal place_1235_succs : BooleanArray(0 downto 0);
  signal place_1235_token : boolean;
  signal place_1236_preds : BooleanArray(0 downto 0);
  signal place_1236_succs : BooleanArray(0 downto 0);
  signal place_1236_token : boolean;
  signal place_1237_preds : BooleanArray(0 downto 0);
  signal place_1237_succs : BooleanArray(0 downto 0);
  signal place_1237_token : boolean;
  signal place_1238_preds : BooleanArray(0 downto 0);
  signal place_1238_succs : BooleanArray(0 downto 0);
  signal place_1238_token : boolean;
  signal place_1239_preds : BooleanArray(0 downto 0);
  signal place_1239_succs : BooleanArray(0 downto 0);
  signal place_1239_token : boolean;
  signal place_1240_preds : BooleanArray(0 downto 0);
  signal place_1240_succs : BooleanArray(0 downto 0);
  signal place_1240_token : boolean;
  signal place_1241_preds : BooleanArray(0 downto 0);
  signal place_1241_succs : BooleanArray(0 downto 0);
  signal place_1241_token : boolean;
  signal place_1242_preds : BooleanArray(0 downto 0);
  signal place_1242_succs : BooleanArray(0 downto 0);
  signal place_1242_token : boolean;
  signal place_1243_preds : BooleanArray(0 downto 0);
  signal place_1243_succs : BooleanArray(0 downto 0);
  signal place_1243_token : boolean;
  signal place_1244_preds : BooleanArray(0 downto 0);
  signal place_1244_succs : BooleanArray(0 downto 0);
  signal place_1244_token : boolean;
  signal place_1245_preds : BooleanArray(0 downto 0);
  signal place_1245_succs : BooleanArray(0 downto 0);
  signal place_1245_token : boolean;
  signal place_1246_preds : BooleanArray(0 downto 0);
  signal place_1246_succs : BooleanArray(0 downto 0);
  signal place_1246_token : boolean;
  signal place_1247_preds : BooleanArray(0 downto 0);
  signal place_1247_succs : BooleanArray(0 downto 0);
  signal place_1247_token : boolean;
  signal place_1248_preds : BooleanArray(0 downto 0);
  signal place_1248_succs : BooleanArray(0 downto 0);
  signal place_1248_token : boolean;
  signal place_1249_preds : BooleanArray(0 downto 0);
  signal place_1249_succs : BooleanArray(0 downto 0);
  signal place_1249_token : boolean;
  signal place_1250_preds : BooleanArray(0 downto 0);
  signal place_1250_succs : BooleanArray(0 downto 0);
  signal place_1250_token : boolean;
  signal place_1251_preds : BooleanArray(0 downto 0);
  signal place_1251_succs : BooleanArray(0 downto 0);
  signal place_1251_token : boolean;
  signal place_1252_preds : BooleanArray(0 downto 0);
  signal place_1252_succs : BooleanArray(0 downto 0);
  signal place_1252_token : boolean;
  signal place_1253_preds : BooleanArray(0 downto 0);
  signal place_1253_succs : BooleanArray(0 downto 0);
  signal place_1253_token : boolean;
  signal place_1254_preds : BooleanArray(0 downto 0);
  signal place_1254_succs : BooleanArray(0 downto 0);
  signal place_1254_token : boolean;
  signal place_1255_preds : BooleanArray(0 downto 0);
  signal place_1255_succs : BooleanArray(0 downto 0);
  signal place_1255_token : boolean;
  signal place_1256_preds : BooleanArray(0 downto 0);
  signal place_1256_succs : BooleanArray(0 downto 0);
  signal place_1256_token : boolean;
  signal place_1257_preds : BooleanArray(0 downto 0);
  signal place_1257_succs : BooleanArray(0 downto 0);
  signal place_1257_token : boolean;
  signal place_1258_preds : BooleanArray(0 downto 0);
  signal place_1258_succs : BooleanArray(0 downto 0);
  signal place_1258_token : boolean;
  signal place_1259_preds : BooleanArray(0 downto 0);
  signal place_1259_succs : BooleanArray(0 downto 0);
  signal place_1259_token : boolean;
  signal place_1260_preds : BooleanArray(0 downto 0);
  signal place_1260_succs : BooleanArray(0 downto 0);
  signal place_1260_token : boolean;
  signal place_1261_preds : BooleanArray(0 downto 0);
  signal place_1261_succs : BooleanArray(0 downto 0);
  signal place_1261_token : boolean;
  signal place_1262_preds : BooleanArray(0 downto 0);
  signal place_1262_succs : BooleanArray(0 downto 0);
  signal place_1262_token : boolean;
  signal place_1263_preds : BooleanArray(0 downto 0);
  signal place_1263_succs : BooleanArray(0 downto 0);
  signal place_1263_token : boolean;
  signal place_1264_preds : BooleanArray(0 downto 0);
  signal place_1264_succs : BooleanArray(0 downto 0);
  signal place_1264_token : boolean;
  signal place_1265_preds : BooleanArray(0 downto 0);
  signal place_1265_succs : BooleanArray(0 downto 0);
  signal place_1265_token : boolean;
  signal place_1266_preds : BooleanArray(0 downto 0);
  signal place_1266_succs : BooleanArray(0 downto 0);
  signal place_1266_token : boolean;
  signal place_1267_preds : BooleanArray(0 downto 0);
  signal place_1267_succs : BooleanArray(0 downto 0);
  signal place_1267_token : boolean;
  signal place_1268_preds : BooleanArray(0 downto 0);
  signal place_1268_succs : BooleanArray(0 downto 0);
  signal place_1268_token : boolean;
  signal place_1269_preds : BooleanArray(0 downto 0);
  signal place_1269_succs : BooleanArray(0 downto 0);
  signal place_1269_token : boolean;
  signal place_1270_preds : BooleanArray(0 downto 0);
  signal place_1270_succs : BooleanArray(0 downto 0);
  signal place_1270_token : boolean;
  signal place_1271_preds : BooleanArray(0 downto 0);
  signal place_1271_succs : BooleanArray(0 downto 0);
  signal place_1271_token : boolean;
  signal place_1272_preds : BooleanArray(0 downto 0);
  signal place_1272_succs : BooleanArray(0 downto 0);
  signal place_1272_token : boolean;
  signal place_1273_preds : BooleanArray(0 downto 0);
  signal place_1273_succs : BooleanArray(0 downto 0);
  signal place_1273_token : boolean;
  signal place_1274_preds : BooleanArray(0 downto 0);
  signal place_1274_succs : BooleanArray(0 downto 0);
  signal place_1274_token : boolean;
  signal place_1275_preds : BooleanArray(0 downto 0);
  signal place_1275_succs : BooleanArray(0 downto 0);
  signal place_1275_token : boolean;
  signal place_1276_preds : BooleanArray(0 downto 0);
  signal place_1276_succs : BooleanArray(0 downto 0);
  signal place_1276_token : boolean;
  signal place_1277_preds : BooleanArray(0 downto 0);
  signal place_1277_succs : BooleanArray(0 downto 0);
  signal place_1277_token : boolean;
  signal place_1278_preds : BooleanArray(0 downto 0);
  signal place_1278_succs : BooleanArray(0 downto 0);
  signal place_1278_token : boolean;
  signal place_1279_preds : BooleanArray(0 downto 0);
  signal place_1279_succs : BooleanArray(0 downto 0);
  signal place_1279_token : boolean;
  signal place_1280_preds : BooleanArray(0 downto 0);
  signal place_1280_succs : BooleanArray(0 downto 0);
  signal place_1280_token : boolean;
  signal place_1281_preds : BooleanArray(0 downto 0);
  signal place_1281_succs : BooleanArray(0 downto 0);
  signal place_1281_token : boolean;
  signal place_1282_preds : BooleanArray(0 downto 0);
  signal place_1282_succs : BooleanArray(0 downto 0);
  signal place_1282_token : boolean;
  signal place_1283_preds : BooleanArray(0 downto 0);
  signal place_1283_succs : BooleanArray(0 downto 0);
  signal place_1283_token : boolean;
  signal place_1284_preds : BooleanArray(0 downto 0);
  signal place_1284_succs : BooleanArray(0 downto 0);
  signal place_1284_token : boolean;
  signal place_1285_preds : BooleanArray(0 downto 0);
  signal place_1285_succs : BooleanArray(0 downto 0);
  signal place_1285_token : boolean;
  signal place_1286_preds : BooleanArray(0 downto 0);
  signal place_1286_succs : BooleanArray(0 downto 0);
  signal place_1286_token : boolean;
  signal place_1287_preds : BooleanArray(0 downto 0);
  signal place_1287_succs : BooleanArray(0 downto 0);
  signal place_1287_token : boolean;
  signal place_1288_preds : BooleanArray(0 downto 0);
  signal place_1288_succs : BooleanArray(0 downto 0);
  signal place_1288_token : boolean;
  signal place_1289_preds : BooleanArray(0 downto 0);
  signal place_1289_succs : BooleanArray(0 downto 0);
  signal place_1289_token : boolean;
  signal place_1290_preds : BooleanArray(0 downto 0);
  signal place_1290_succs : BooleanArray(0 downto 0);
  signal place_1290_token : boolean;
  signal place_1291_preds : BooleanArray(0 downto 0);
  signal place_1291_succs : BooleanArray(0 downto 0);
  signal place_1291_token : boolean;
  signal place_1292_preds : BooleanArray(0 downto 0);
  signal place_1292_succs : BooleanArray(0 downto 0);
  signal place_1292_token : boolean;
  signal place_1293_preds : BooleanArray(0 downto 0);
  signal place_1293_succs : BooleanArray(0 downto 0);
  signal place_1293_token : boolean;
  signal place_1294_preds : BooleanArray(0 downto 0);
  signal place_1294_succs : BooleanArray(0 downto 0);
  signal place_1294_token : boolean;
  signal place_1295_preds : BooleanArray(0 downto 0);
  signal place_1295_succs : BooleanArray(0 downto 0);
  signal place_1295_token : boolean;
  signal place_1296_preds : BooleanArray(0 downto 0);
  signal place_1296_succs : BooleanArray(0 downto 0);
  signal place_1296_token : boolean;
  signal place_1297_preds : BooleanArray(0 downto 0);
  signal place_1297_succs : BooleanArray(0 downto 0);
  signal place_1297_token : boolean;
  signal place_1298_preds : BooleanArray(0 downto 0);
  signal place_1298_succs : BooleanArray(0 downto 0);
  signal place_1298_token : boolean;
  signal place_1299_preds : BooleanArray(0 downto 0);
  signal place_1299_succs : BooleanArray(0 downto 0);
  signal place_1299_token : boolean;
  signal place_1300_preds : BooleanArray(0 downto 0);
  signal place_1300_succs : BooleanArray(0 downto 0);
  signal place_1300_token : boolean;
  signal place_1301_preds : BooleanArray(0 downto 0);
  signal place_1301_succs : BooleanArray(0 downto 0);
  signal place_1301_token : boolean;
  signal place_1302_preds : BooleanArray(0 downto 0);
  signal place_1302_succs : BooleanArray(0 downto 0);
  signal place_1302_token : boolean;
  signal place_1303_preds : BooleanArray(0 downto 0);
  signal place_1303_succs : BooleanArray(0 downto 0);
  signal place_1303_token : boolean;
  signal place_1304_preds : BooleanArray(0 downto 0);
  signal place_1304_succs : BooleanArray(0 downto 0);
  signal place_1304_token : boolean;
  signal place_1305_preds : BooleanArray(0 downto 0);
  signal place_1305_succs : BooleanArray(0 downto 0);
  signal place_1305_token : boolean;
  signal place_1306_preds : BooleanArray(0 downto 0);
  signal place_1306_succs : BooleanArray(0 downto 0);
  signal place_1306_token : boolean;
  signal place_1307_preds : BooleanArray(0 downto 0);
  signal place_1307_succs : BooleanArray(0 downto 0);
  signal place_1307_token : boolean;
  signal place_1308_preds : BooleanArray(0 downto 0);
  signal place_1308_succs : BooleanArray(0 downto 0);
  signal place_1308_token : boolean;
  signal place_1309_preds : BooleanArray(0 downto 0);
  signal place_1309_succs : BooleanArray(0 downto 0);
  signal place_1309_token : boolean;
  signal place_1310_preds : BooleanArray(0 downto 0);
  signal place_1310_succs : BooleanArray(0 downto 0);
  signal place_1310_token : boolean;
  signal place_1311_preds : BooleanArray(0 downto 0);
  signal place_1311_succs : BooleanArray(0 downto 0);
  signal place_1311_token : boolean;
  signal place_1312_preds : BooleanArray(0 downto 0);
  signal place_1312_succs : BooleanArray(0 downto 0);
  signal place_1312_token : boolean;
  signal place_1313_preds : BooleanArray(0 downto 0);
  signal place_1313_succs : BooleanArray(0 downto 0);
  signal place_1313_token : boolean;
  signal place_1314_preds : BooleanArray(0 downto 0);
  signal place_1314_succs : BooleanArray(0 downto 0);
  signal place_1314_token : boolean;
  signal place_1315_preds : BooleanArray(0 downto 0);
  signal place_1315_succs : BooleanArray(0 downto 0);
  signal place_1315_token : boolean;
  signal place_1316_preds : BooleanArray(0 downto 0);
  signal place_1316_succs : BooleanArray(0 downto 0);
  signal place_1316_token : boolean;
  signal place_1317_preds : BooleanArray(0 downto 0);
  signal place_1317_succs : BooleanArray(0 downto 0);
  signal place_1317_token : boolean;
  signal place_1318_preds : BooleanArray(0 downto 0);
  signal place_1318_succs : BooleanArray(0 downto 0);
  signal place_1318_token : boolean;
  signal place_1319_preds : BooleanArray(0 downto 0);
  signal place_1319_succs : BooleanArray(0 downto 0);
  signal place_1319_token : boolean;
  signal place_1320_preds : BooleanArray(0 downto 0);
  signal place_1320_succs : BooleanArray(0 downto 0);
  signal place_1320_token : boolean;
  signal place_1321_preds : BooleanArray(0 downto 0);
  signal place_1321_succs : BooleanArray(0 downto 0);
  signal place_1321_token : boolean;
  signal place_1322_preds : BooleanArray(0 downto 0);
  signal place_1322_succs : BooleanArray(0 downto 0);
  signal place_1322_token : boolean;
  signal place_1323_preds : BooleanArray(0 downto 0);
  signal place_1323_succs : BooleanArray(0 downto 0);
  signal place_1323_token : boolean;
  signal place_1324_preds : BooleanArray(0 downto 0);
  signal place_1324_succs : BooleanArray(0 downto 0);
  signal place_1324_token : boolean;
  signal place_1325_preds : BooleanArray(0 downto 0);
  signal place_1325_succs : BooleanArray(0 downto 0);
  signal place_1325_token : boolean;
  signal place_1326_preds : BooleanArray(0 downto 0);
  signal place_1326_succs : BooleanArray(0 downto 0);
  signal place_1326_token : boolean;
  signal place_1327_preds : BooleanArray(0 downto 0);
  signal place_1327_succs : BooleanArray(0 downto 0);
  signal place_1327_token : boolean;
  signal place_1328_preds : BooleanArray(0 downto 0);
  signal place_1328_succs : BooleanArray(0 downto 0);
  signal place_1328_token : boolean;
  signal place_1329_preds : BooleanArray(0 downto 0);
  signal place_1329_succs : BooleanArray(0 downto 0);
  signal place_1329_token : boolean;
  signal place_1330_preds : BooleanArray(0 downto 0);
  signal place_1330_succs : BooleanArray(0 downto 0);
  signal place_1330_token : boolean;
  signal place_1331_preds : BooleanArray(0 downto 0);
  signal place_1331_succs : BooleanArray(0 downto 0);
  signal place_1331_token : boolean;
  signal place_1332_preds : BooleanArray(0 downto 0);
  signal place_1332_succs : BooleanArray(0 downto 0);
  signal place_1332_token : boolean;
  signal place_1333_preds : BooleanArray(0 downto 0);
  signal place_1333_succs : BooleanArray(0 downto 0);
  signal place_1333_token : boolean;
  signal place_1334_preds : BooleanArray(0 downto 0);
  signal place_1334_succs : BooleanArray(0 downto 0);
  signal place_1334_token : boolean;
  signal place_1335_preds : BooleanArray(0 downto 0);
  signal place_1335_succs : BooleanArray(0 downto 0);
  signal place_1335_token : boolean;
  signal place_1336_preds : BooleanArray(0 downto 0);
  signal place_1336_succs : BooleanArray(0 downto 0);
  signal place_1336_token : boolean;
  signal place_1337_preds : BooleanArray(0 downto 0);
  signal place_1337_succs : BooleanArray(0 downto 0);
  signal place_1337_token : boolean;
  signal place_1338_preds : BooleanArray(0 downto 0);
  signal place_1338_succs : BooleanArray(0 downto 0);
  signal place_1338_token : boolean;
  signal place_1339_preds : BooleanArray(0 downto 0);
  signal place_1339_succs : BooleanArray(0 downto 0);
  signal place_1339_token : boolean;
  signal place_1340_preds : BooleanArray(0 downto 0);
  signal place_1340_succs : BooleanArray(0 downto 0);
  signal place_1340_token : boolean;
  signal place_1341_preds : BooleanArray(0 downto 0);
  signal place_1341_succs : BooleanArray(0 downto 0);
  signal place_1341_token : boolean;
  signal place_1342_preds : BooleanArray(0 downto 0);
  signal place_1342_succs : BooleanArray(0 downto 0);
  signal place_1342_token : boolean;
  signal place_1343_preds : BooleanArray(0 downto 0);
  signal place_1343_succs : BooleanArray(0 downto 0);
  signal place_1343_token : boolean;
  signal place_1344_preds : BooleanArray(0 downto 0);
  signal place_1344_succs : BooleanArray(0 downto 0);
  signal place_1344_token : boolean;
  signal place_1345_preds : BooleanArray(0 downto 0);
  signal place_1345_succs : BooleanArray(0 downto 0);
  signal place_1345_token : boolean;
  signal place_1346_preds : BooleanArray(0 downto 0);
  signal place_1346_succs : BooleanArray(0 downto 0);
  signal place_1346_token : boolean;
  signal place_1347_preds : BooleanArray(0 downto 0);
  signal place_1347_succs : BooleanArray(0 downto 0);
  signal place_1347_token : boolean;
  signal place_1348_preds : BooleanArray(0 downto 0);
  signal place_1348_succs : BooleanArray(0 downto 0);
  signal place_1348_token : boolean;
  signal place_1349_preds : BooleanArray(0 downto 0);
  signal place_1349_succs : BooleanArray(0 downto 0);
  signal place_1349_token : boolean;
  signal place_1350_preds : BooleanArray(0 downto 0);
  signal place_1350_succs : BooleanArray(0 downto 0);
  signal place_1350_token : boolean;
  signal place_1351_preds : BooleanArray(0 downto 0);
  signal place_1351_succs : BooleanArray(0 downto 0);
  signal place_1351_token : boolean;
  signal place_1352_preds : BooleanArray(0 downto 0);
  signal place_1352_succs : BooleanArray(0 downto 0);
  signal place_1352_token : boolean;
  signal place_1353_preds : BooleanArray(0 downto 0);
  signal place_1353_succs : BooleanArray(0 downto 0);
  signal place_1353_token : boolean;
  signal place_1354_preds : BooleanArray(0 downto 0);
  signal place_1354_succs : BooleanArray(0 downto 0);
  signal place_1354_token : boolean;
  signal place_1355_preds : BooleanArray(0 downto 0);
  signal place_1355_succs : BooleanArray(0 downto 0);
  signal place_1355_token : boolean;
  signal place_1356_preds : BooleanArray(0 downto 0);
  signal place_1356_succs : BooleanArray(0 downto 0);
  signal place_1356_token : boolean;
  signal place_1357_preds : BooleanArray(0 downto 0);
  signal place_1357_succs : BooleanArray(0 downto 0);
  signal place_1357_token : boolean;
  signal place_1358_preds : BooleanArray(0 downto 0);
  signal place_1358_succs : BooleanArray(0 downto 0);
  signal place_1358_token : boolean;
  signal place_1359_preds : BooleanArray(0 downto 0);
  signal place_1359_succs : BooleanArray(0 downto 0);
  signal place_1359_token : boolean;
  signal place_1360_preds : BooleanArray(0 downto 0);
  signal place_1360_succs : BooleanArray(0 downto 0);
  signal place_1360_token : boolean;
  signal place_1361_preds : BooleanArray(0 downto 0);
  signal place_1361_succs : BooleanArray(0 downto 0);
  signal place_1361_token : boolean;
  signal place_1362_preds : BooleanArray(0 downto 0);
  signal place_1362_succs : BooleanArray(0 downto 0);
  signal place_1362_token : boolean;
  signal place_1363_preds : BooleanArray(0 downto 0);
  signal place_1363_succs : BooleanArray(0 downto 0);
  signal place_1363_token : boolean;
  signal place_1364_preds : BooleanArray(0 downto 0);
  signal place_1364_succs : BooleanArray(0 downto 0);
  signal place_1364_token : boolean;
  signal place_1365_preds : BooleanArray(0 downto 0);
  signal place_1365_succs : BooleanArray(0 downto 0);
  signal place_1365_token : boolean;
  signal place_1366_preds : BooleanArray(0 downto 0);
  signal place_1366_succs : BooleanArray(0 downto 0);
  signal place_1366_token : boolean;
  signal place_1367_preds : BooleanArray(0 downto 0);
  signal place_1367_succs : BooleanArray(0 downto 0);
  signal place_1367_token : boolean;
  signal place_1368_preds : BooleanArray(0 downto 0);
  signal place_1368_succs : BooleanArray(0 downto 0);
  signal place_1368_token : boolean;
  signal place_1369_preds : BooleanArray(0 downto 0);
  signal place_1369_succs : BooleanArray(0 downto 0);
  signal place_1369_token : boolean;
  signal place_1370_preds : BooleanArray(0 downto 0);
  signal place_1370_succs : BooleanArray(0 downto 0);
  signal place_1370_token : boolean;
  signal place_1371_preds : BooleanArray(0 downto 0);
  signal place_1371_succs : BooleanArray(0 downto 0);
  signal place_1371_token : boolean;
  signal place_1372_preds : BooleanArray(0 downto 0);
  signal place_1372_succs : BooleanArray(0 downto 0);
  signal place_1372_token : boolean;
  signal place_1373_preds : BooleanArray(0 downto 0);
  signal place_1373_succs : BooleanArray(0 downto 0);
  signal place_1373_token : boolean;
  signal place_1374_preds : BooleanArray(0 downto 0);
  signal place_1374_succs : BooleanArray(0 downto 0);
  signal place_1374_token : boolean;
  signal place_1375_preds : BooleanArray(0 downto 0);
  signal place_1375_succs : BooleanArray(0 downto 0);
  signal place_1375_token : boolean;
  signal place_1376_preds : BooleanArray(0 downto 0);
  signal place_1376_succs : BooleanArray(0 downto 0);
  signal place_1376_token : boolean;
  signal place_1377_preds : BooleanArray(0 downto 0);
  signal place_1377_succs : BooleanArray(0 downto 0);
  signal place_1377_token : boolean;
  signal place_1378_preds : BooleanArray(0 downto 0);
  signal place_1378_succs : BooleanArray(0 downto 0);
  signal place_1378_token : boolean;
  signal place_1379_preds : BooleanArray(0 downto 0);
  signal place_1379_succs : BooleanArray(0 downto 0);
  signal place_1379_token : boolean;
  signal place_1380_preds : BooleanArray(0 downto 0);
  signal place_1380_succs : BooleanArray(0 downto 0);
  signal place_1380_token : boolean;
  signal place_1381_preds : BooleanArray(0 downto 0);
  signal place_1381_succs : BooleanArray(0 downto 0);
  signal place_1381_token : boolean;
  signal place_1382_preds : BooleanArray(0 downto 0);
  signal place_1382_succs : BooleanArray(0 downto 0);
  signal place_1382_token : boolean;
  signal place_1383_preds : BooleanArray(0 downto 0);
  signal place_1383_succs : BooleanArray(0 downto 0);
  signal place_1383_token : boolean;
  signal place_1384_preds : BooleanArray(0 downto 0);
  signal place_1384_succs : BooleanArray(0 downto 0);
  signal place_1384_token : boolean;
  signal place_1385_preds : BooleanArray(0 downto 0);
  signal place_1385_succs : BooleanArray(0 downto 0);
  signal place_1385_token : boolean;
  signal place_1386_preds : BooleanArray(0 downto 0);
  signal place_1386_succs : BooleanArray(0 downto 0);
  signal place_1386_token : boolean;
  signal place_1387_preds : BooleanArray(0 downto 0);
  signal place_1387_succs : BooleanArray(0 downto 0);
  signal place_1387_token : boolean;
  signal place_1388_preds : BooleanArray(0 downto 0);
  signal place_1388_succs : BooleanArray(0 downto 0);
  signal place_1388_token : boolean;
  signal place_1389_preds : BooleanArray(0 downto 0);
  signal place_1389_succs : BooleanArray(0 downto 0);
  signal place_1389_token : boolean;
  signal place_1390_preds : BooleanArray(0 downto 0);
  signal place_1390_succs : BooleanArray(0 downto 0);
  signal place_1390_token : boolean;
  signal place_1391_preds : BooleanArray(0 downto 0);
  signal place_1391_succs : BooleanArray(0 downto 0);
  signal place_1391_token : boolean;
  signal place_1392_preds : BooleanArray(0 downto 0);
  signal place_1392_succs : BooleanArray(0 downto 0);
  signal place_1392_token : boolean;
  signal place_1393_preds : BooleanArray(0 downto 0);
  signal place_1393_succs : BooleanArray(0 downto 0);
  signal place_1393_token : boolean;
  signal place_1394_preds : BooleanArray(0 downto 0);
  signal place_1394_succs : BooleanArray(0 downto 0);
  signal place_1394_token : boolean;
  signal place_1395_preds : BooleanArray(0 downto 0);
  signal place_1395_succs : BooleanArray(0 downto 0);
  signal place_1395_token : boolean;
  signal place_1396_preds : BooleanArray(0 downto 0);
  signal place_1396_succs : BooleanArray(0 downto 0);
  signal place_1396_token : boolean;
  signal place_1397_preds : BooleanArray(0 downto 0);
  signal place_1397_succs : BooleanArray(0 downto 0);
  signal place_1397_token : boolean;
  signal place_1398_preds : BooleanArray(0 downto 0);
  signal place_1398_succs : BooleanArray(0 downto 0);
  signal place_1398_token : boolean;
  signal place_1399_preds : BooleanArray(0 downto 0);
  signal place_1399_succs : BooleanArray(0 downto 0);
  signal place_1399_token : boolean;
  signal place_1400_preds : BooleanArray(0 downto 0);
  signal place_1400_succs : BooleanArray(0 downto 0);
  signal place_1400_token : boolean;
  signal place_1401_preds : BooleanArray(0 downto 0);
  signal place_1401_succs : BooleanArray(0 downto 0);
  signal place_1401_token : boolean;
  signal place_1402_preds : BooleanArray(0 downto 0);
  signal place_1402_succs : BooleanArray(0 downto 0);
  signal place_1402_token : boolean;
  signal place_1403_preds : BooleanArray(0 downto 0);
  signal place_1403_succs : BooleanArray(0 downto 0);
  signal place_1403_token : boolean;
  signal place_1404_preds : BooleanArray(0 downto 0);
  signal place_1404_succs : BooleanArray(0 downto 0);
  signal place_1404_token : boolean;
  signal place_1405_preds : BooleanArray(0 downto 0);
  signal place_1405_succs : BooleanArray(0 downto 0);
  signal place_1405_token : boolean;
  signal place_1406_preds : BooleanArray(0 downto 0);
  signal place_1406_succs : BooleanArray(0 downto 0);
  signal place_1406_token : boolean;
  signal place_1407_preds : BooleanArray(0 downto 0);
  signal place_1407_succs : BooleanArray(0 downto 0);
  signal place_1407_token : boolean;
  signal place_1408_preds : BooleanArray(0 downto 0);
  signal place_1408_succs : BooleanArray(0 downto 0);
  signal place_1408_token : boolean;
  signal place_1409_preds : BooleanArray(0 downto 0);
  signal place_1409_succs : BooleanArray(0 downto 0);
  signal place_1409_token : boolean;
  signal place_1410_preds : BooleanArray(0 downto 0);
  signal place_1410_succs : BooleanArray(0 downto 0);
  signal place_1410_token : boolean;
  signal place_1411_preds : BooleanArray(0 downto 0);
  signal place_1411_succs : BooleanArray(0 downto 0);
  signal place_1411_token : boolean;
  signal place_1412_preds : BooleanArray(0 downto 0);
  signal place_1412_succs : BooleanArray(0 downto 0);
  signal place_1412_token : boolean;
  signal place_1413_preds : BooleanArray(0 downto 0);
  signal place_1413_succs : BooleanArray(0 downto 0);
  signal place_1413_token : boolean;
  signal place_1414_preds : BooleanArray(0 downto 0);
  signal place_1414_succs : BooleanArray(0 downto 0);
  signal place_1414_token : boolean;
  signal place_1415_preds : BooleanArray(0 downto 0);
  signal place_1415_succs : BooleanArray(0 downto 0);
  signal place_1415_token : boolean;
  signal place_1416_preds : BooleanArray(0 downto 0);
  signal place_1416_succs : BooleanArray(0 downto 0);
  signal place_1416_token : boolean;
  signal place_1417_preds : BooleanArray(0 downto 0);
  signal place_1417_succs : BooleanArray(0 downto 0);
  signal place_1417_token : boolean;
  signal place_1418_preds : BooleanArray(0 downto 0);
  signal place_1418_succs : BooleanArray(0 downto 0);
  signal place_1418_token : boolean;
  signal place_1419_preds : BooleanArray(0 downto 0);
  signal place_1419_succs : BooleanArray(0 downto 0);
  signal place_1419_token : boolean;
  signal place_1420_preds : BooleanArray(0 downto 0);
  signal place_1420_succs : BooleanArray(0 downto 0);
  signal place_1420_token : boolean;
  signal place_1421_preds : BooleanArray(0 downto 0);
  signal place_1421_succs : BooleanArray(0 downto 0);
  signal place_1421_token : boolean;
  signal place_1422_preds : BooleanArray(0 downto 0);
  signal place_1422_succs : BooleanArray(0 downto 0);
  signal place_1422_token : boolean;
  signal place_1423_preds : BooleanArray(0 downto 0);
  signal place_1423_succs : BooleanArray(0 downto 0);
  signal place_1423_token : boolean;
  signal place_1424_preds : BooleanArray(0 downto 0);
  signal place_1424_succs : BooleanArray(0 downto 0);
  signal place_1424_token : boolean;
  signal place_1425_preds : BooleanArray(0 downto 0);
  signal place_1425_succs : BooleanArray(0 downto 0);
  signal place_1425_token : boolean;
  signal place_1426_preds : BooleanArray(0 downto 0);
  signal place_1426_succs : BooleanArray(0 downto 0);
  signal place_1426_token : boolean;
  signal place_1427_preds : BooleanArray(0 downto 0);
  signal place_1427_succs : BooleanArray(0 downto 0);
  signal place_1427_token : boolean;
  signal place_1428_preds : BooleanArray(0 downto 0);
  signal place_1428_succs : BooleanArray(0 downto 0);
  signal place_1428_token : boolean;
  signal place_1429_preds : BooleanArray(0 downto 0);
  signal place_1429_succs : BooleanArray(0 downto 0);
  signal place_1429_token : boolean;
  signal place_1430_preds : BooleanArray(0 downto 0);
  signal place_1430_succs : BooleanArray(0 downto 0);
  signal place_1430_token : boolean;
  signal place_1431_preds : BooleanArray(0 downto 0);
  signal place_1431_succs : BooleanArray(0 downto 0);
  signal place_1431_token : boolean;
  signal place_1432_preds : BooleanArray(0 downto 0);
  signal place_1432_succs : BooleanArray(0 downto 0);
  signal place_1432_token : boolean;
  signal place_1433_preds : BooleanArray(0 downto 0);
  signal place_1433_succs : BooleanArray(0 downto 0);
  signal place_1433_token : boolean;
  signal place_1434_preds : BooleanArray(0 downto 0);
  signal place_1434_succs : BooleanArray(0 downto 0);
  signal place_1434_token : boolean;
  signal place_1435_preds : BooleanArray(0 downto 0);
  signal place_1435_succs : BooleanArray(0 downto 0);
  signal place_1435_token : boolean;
  signal place_1436_preds : BooleanArray(0 downto 0);
  signal place_1436_succs : BooleanArray(0 downto 0);
  signal place_1436_token : boolean;
  signal place_1437_preds : BooleanArray(0 downto 0);
  signal place_1437_succs : BooleanArray(0 downto 0);
  signal place_1437_token : boolean;
  signal place_1438_preds : BooleanArray(0 downto 0);
  signal place_1438_succs : BooleanArray(0 downto 0);
  signal place_1438_token : boolean;
  signal place_1439_preds : BooleanArray(0 downto 0);
  signal place_1439_succs : BooleanArray(0 downto 0);
  signal place_1439_token : boolean;
  signal place_1440_preds : BooleanArray(0 downto 0);
  signal place_1440_succs : BooleanArray(0 downto 0);
  signal place_1440_token : boolean;
  signal place_1441_preds : BooleanArray(0 downto 0);
  signal place_1441_succs : BooleanArray(0 downto 0);
  signal place_1441_token : boolean;
  signal place_1442_preds : BooleanArray(0 downto 0);
  signal place_1442_succs : BooleanArray(0 downto 0);
  signal place_1442_token : boolean;
  signal place_1443_preds : BooleanArray(0 downto 0);
  signal place_1443_succs : BooleanArray(0 downto 0);
  signal place_1443_token : boolean;
  signal place_1444_preds : BooleanArray(0 downto 0);
  signal place_1444_succs : BooleanArray(0 downto 0);
  signal place_1444_token : boolean;
  signal place_1445_preds : BooleanArray(0 downto 0);
  signal place_1445_succs : BooleanArray(0 downto 0);
  signal place_1445_token : boolean;
  signal place_1446_preds : BooleanArray(0 downto 0);
  signal place_1446_succs : BooleanArray(0 downto 0);
  signal place_1446_token : boolean;
  signal place_1447_preds : BooleanArray(0 downto 0);
  signal place_1447_succs : BooleanArray(0 downto 0);
  signal place_1447_token : boolean;
  signal place_1448_preds : BooleanArray(0 downto 0);
  signal place_1448_succs : BooleanArray(0 downto 0);
  signal place_1448_token : boolean;
  signal place_1449_preds : BooleanArray(0 downto 0);
  signal place_1449_succs : BooleanArray(0 downto 0);
  signal place_1449_token : boolean;
  signal place_1450_preds : BooleanArray(0 downto 0);
  signal place_1450_succs : BooleanArray(0 downto 0);
  signal place_1450_token : boolean;
  signal place_1451_preds : BooleanArray(0 downto 0);
  signal place_1451_succs : BooleanArray(0 downto 0);
  signal place_1451_token : boolean;
  signal place_1452_preds : BooleanArray(0 downto 0);
  signal place_1452_succs : BooleanArray(0 downto 0);
  signal place_1452_token : boolean;
  signal place_1453_preds : BooleanArray(0 downto 0);
  signal place_1453_succs : BooleanArray(0 downto 0);
  signal place_1453_token : boolean;
  signal place_1454_preds : BooleanArray(0 downto 0);
  signal place_1454_succs : BooleanArray(0 downto 0);
  signal place_1454_token : boolean;
  signal place_1455_preds : BooleanArray(0 downto 0);
  signal place_1455_succs : BooleanArray(0 downto 0);
  signal place_1455_token : boolean;
  signal place_1456_preds : BooleanArray(0 downto 0);
  signal place_1456_succs : BooleanArray(0 downto 0);
  signal place_1456_token : boolean;
  signal place_1457_preds : BooleanArray(0 downto 0);
  signal place_1457_succs : BooleanArray(0 downto 0);
  signal place_1457_token : boolean;
  signal place_1458_preds : BooleanArray(0 downto 0);
  signal place_1458_succs : BooleanArray(0 downto 0);
  signal place_1458_token : boolean;
  signal place_1459_preds : BooleanArray(0 downto 0);
  signal place_1459_succs : BooleanArray(0 downto 0);
  signal place_1459_token : boolean;
  signal place_1460_preds : BooleanArray(0 downto 0);
  signal place_1460_succs : BooleanArray(0 downto 0);
  signal place_1460_token : boolean;
  signal place_1461_preds : BooleanArray(0 downto 0);
  signal place_1461_succs : BooleanArray(0 downto 0);
  signal place_1461_token : boolean;
  signal place_1462_preds : BooleanArray(0 downto 0);
  signal place_1462_succs : BooleanArray(0 downto 0);
  signal place_1462_token : boolean;
  signal place_1463_preds : BooleanArray(0 downto 0);
  signal place_1463_succs : BooleanArray(0 downto 0);
  signal place_1463_token : boolean;
  signal place_1464_preds : BooleanArray(0 downto 0);
  signal place_1464_succs : BooleanArray(0 downto 0);
  signal place_1464_token : boolean;
  signal place_1465_preds : BooleanArray(0 downto 0);
  signal place_1465_succs : BooleanArray(0 downto 0);
  signal place_1465_token : boolean;
  signal place_1466_preds : BooleanArray(0 downto 0);
  signal place_1466_succs : BooleanArray(0 downto 0);
  signal place_1466_token : boolean;
  signal place_1467_preds : BooleanArray(0 downto 0);
  signal place_1467_succs : BooleanArray(0 downto 0);
  signal place_1467_token : boolean;
  signal place_1468_preds : BooleanArray(0 downto 0);
  signal place_1468_succs : BooleanArray(0 downto 0);
  signal place_1468_token : boolean;
  signal place_1469_preds : BooleanArray(0 downto 0);
  signal place_1469_succs : BooleanArray(0 downto 0);
  signal place_1469_token : boolean;
  signal place_1470_preds : BooleanArray(0 downto 0);
  signal place_1470_succs : BooleanArray(0 downto 0);
  signal place_1470_token : boolean;
  signal place_1471_preds : BooleanArray(0 downto 0);
  signal place_1471_succs : BooleanArray(0 downto 0);
  signal place_1471_token : boolean;
  signal place_1472_preds : BooleanArray(0 downto 0);
  signal place_1472_succs : BooleanArray(0 downto 0);
  signal place_1472_token : boolean;
  signal place_1473_preds : BooleanArray(0 downto 0);
  signal place_1473_succs : BooleanArray(0 downto 0);
  signal place_1473_token : boolean;
  signal place_1474_preds : BooleanArray(0 downto 0);
  signal place_1474_succs : BooleanArray(0 downto 0);
  signal place_1474_token : boolean;
  signal place_1475_preds : BooleanArray(0 downto 0);
  signal place_1475_succs : BooleanArray(0 downto 0);
  signal place_1475_token : boolean;
  signal place_1476_preds : BooleanArray(0 downto 0);
  signal place_1476_succs : BooleanArray(0 downto 0);
  signal place_1476_token : boolean;
  signal place_1477_preds : BooleanArray(0 downto 0);
  signal place_1477_succs : BooleanArray(0 downto 0);
  signal place_1477_token : boolean;
  signal place_1478_preds : BooleanArray(0 downto 0);
  signal place_1478_succs : BooleanArray(0 downto 0);
  signal place_1478_token : boolean;
  signal place_1479_preds : BooleanArray(0 downto 0);
  signal place_1479_succs : BooleanArray(0 downto 0);
  signal place_1479_token : boolean;
  signal place_1480_preds : BooleanArray(0 downto 0);
  signal place_1480_succs : BooleanArray(0 downto 0);
  signal place_1480_token : boolean;
  signal place_1481_preds : BooleanArray(0 downto 0);
  signal place_1481_succs : BooleanArray(0 downto 0);
  signal place_1481_token : boolean;
  signal place_1482_preds : BooleanArray(0 downto 0);
  signal place_1482_succs : BooleanArray(0 downto 0);
  signal place_1482_token : boolean;
  signal place_1483_preds : BooleanArray(0 downto 0);
  signal place_1483_succs : BooleanArray(0 downto 0);
  signal place_1483_token : boolean;
  signal place_1484_preds : BooleanArray(0 downto 0);
  signal place_1484_succs : BooleanArray(0 downto 0);
  signal place_1484_token : boolean;
  signal place_1485_preds : BooleanArray(0 downto 0);
  signal place_1485_succs : BooleanArray(0 downto 0);
  signal place_1485_token : boolean;
  signal place_1486_preds : BooleanArray(0 downto 0);
  signal place_1486_succs : BooleanArray(0 downto 0);
  signal place_1486_token : boolean;
  signal place_1487_preds : BooleanArray(0 downto 0);
  signal place_1487_succs : BooleanArray(0 downto 0);
  signal place_1487_token : boolean;
  signal place_1488_preds : BooleanArray(0 downto 0);
  signal place_1488_succs : BooleanArray(0 downto 0);
  signal place_1488_token : boolean;
  signal place_1489_preds : BooleanArray(0 downto 0);
  signal place_1489_succs : BooleanArray(0 downto 0);
  signal place_1489_token : boolean;
  signal place_1490_preds : BooleanArray(0 downto 0);
  signal place_1490_succs : BooleanArray(0 downto 0);
  signal place_1490_token : boolean;
  signal place_1491_preds : BooleanArray(0 downto 0);
  signal place_1491_succs : BooleanArray(0 downto 0);
  signal place_1491_token : boolean;
  signal place_1492_preds : BooleanArray(0 downto 0);
  signal place_1492_succs : BooleanArray(0 downto 0);
  signal place_1492_token : boolean;
  signal place_1493_preds : BooleanArray(0 downto 0);
  signal place_1493_succs : BooleanArray(0 downto 0);
  signal place_1493_token : boolean;
  signal place_1494_preds : BooleanArray(0 downto 0);
  signal place_1494_succs : BooleanArray(0 downto 0);
  signal place_1494_token : boolean;
  signal place_1495_preds : BooleanArray(0 downto 0);
  signal place_1495_succs : BooleanArray(0 downto 0);
  signal place_1495_token : boolean;
  signal place_1496_preds : BooleanArray(0 downto 0);
  signal place_1496_succs : BooleanArray(0 downto 0);
  signal place_1496_token : boolean;
  signal place_1497_preds : BooleanArray(0 downto 0);
  signal place_1497_succs : BooleanArray(0 downto 0);
  signal place_1497_token : boolean;
  signal place_1498_preds : BooleanArray(0 downto 0);
  signal place_1498_succs : BooleanArray(0 downto 0);
  signal place_1498_token : boolean;
  signal place_1499_preds : BooleanArray(0 downto 0);
  signal place_1499_succs : BooleanArray(0 downto 0);
  signal place_1499_token : boolean;
  signal place_1500_preds : BooleanArray(0 downto 0);
  signal place_1500_succs : BooleanArray(0 downto 0);
  signal place_1500_token : boolean;
  signal place_1501_preds : BooleanArray(0 downto 0);
  signal place_1501_succs : BooleanArray(0 downto 0);
  signal place_1501_token : boolean;
  signal place_1502_preds : BooleanArray(0 downto 0);
  signal place_1502_succs : BooleanArray(0 downto 0);
  signal place_1502_token : boolean;
  signal place_1503_preds : BooleanArray(0 downto 0);
  signal place_1503_succs : BooleanArray(0 downto 0);
  signal place_1503_token : boolean;
  signal place_1504_preds : BooleanArray(0 downto 0);
  signal place_1504_succs : BooleanArray(0 downto 0);
  signal place_1504_token : boolean;
  signal place_1505_preds : BooleanArray(0 downto 0);
  signal place_1505_succs : BooleanArray(0 downto 0);
  signal place_1505_token : boolean;
  signal place_1506_preds : BooleanArray(0 downto 0);
  signal place_1506_succs : BooleanArray(0 downto 0);
  signal place_1506_token : boolean;
  signal place_1507_preds : BooleanArray(0 downto 0);
  signal place_1507_succs : BooleanArray(0 downto 0);
  signal place_1507_token : boolean;
  signal place_1508_preds : BooleanArray(0 downto 0);
  signal place_1508_succs : BooleanArray(0 downto 0);
  signal place_1508_token : boolean;
  signal place_1509_preds : BooleanArray(0 downto 0);
  signal place_1509_succs : BooleanArray(0 downto 0);
  signal place_1509_token : boolean;
  signal place_1510_preds : BooleanArray(0 downto 0);
  signal place_1510_succs : BooleanArray(0 downto 0);
  signal place_1510_token : boolean;
  signal place_1511_preds : BooleanArray(0 downto 0);
  signal place_1511_succs : BooleanArray(0 downto 0);
  signal place_1511_token : boolean;
  signal place_1512_preds : BooleanArray(0 downto 0);
  signal place_1512_succs : BooleanArray(0 downto 0);
  signal place_1512_token : boolean;
  signal place_1513_preds : BooleanArray(0 downto 0);
  signal place_1513_succs : BooleanArray(0 downto 0);
  signal place_1513_token : boolean;
  signal place_1514_preds : BooleanArray(0 downto 0);
  signal place_1514_succs : BooleanArray(0 downto 0);
  signal place_1514_token : boolean;
  signal place_1515_preds : BooleanArray(0 downto 0);
  signal place_1515_succs : BooleanArray(0 downto 0);
  signal place_1515_token : boolean;
  signal place_1516_preds : BooleanArray(0 downto 0);
  signal place_1516_succs : BooleanArray(0 downto 0);
  signal place_1516_token : boolean;
  signal place_1517_preds : BooleanArray(0 downto 0);
  signal place_1517_succs : BooleanArray(0 downto 0);
  signal place_1517_token : boolean;
  signal place_1518_preds : BooleanArray(0 downto 0);
  signal place_1518_succs : BooleanArray(0 downto 0);
  signal place_1518_token : boolean;
  signal place_1519_preds : BooleanArray(0 downto 0);
  signal place_1519_succs : BooleanArray(0 downto 0);
  signal place_1519_token : boolean;
  signal place_1520_preds : BooleanArray(0 downto 0);
  signal place_1520_succs : BooleanArray(0 downto 0);
  signal place_1520_token : boolean;
  signal place_1521_preds : BooleanArray(0 downto 0);
  signal place_1521_succs : BooleanArray(0 downto 0);
  signal place_1521_token : boolean;
  signal place_1522_preds : BooleanArray(0 downto 0);
  signal place_1522_succs : BooleanArray(0 downto 0);
  signal place_1522_token : boolean;
  signal place_1523_preds : BooleanArray(0 downto 0);
  signal place_1523_succs : BooleanArray(0 downto 0);
  signal place_1523_token : boolean;
  signal place_1524_preds : BooleanArray(0 downto 0);
  signal place_1524_succs : BooleanArray(0 downto 0);
  signal place_1524_token : boolean;
  signal place_1525_preds : BooleanArray(0 downto 0);
  signal place_1525_succs : BooleanArray(0 downto 0);
  signal place_1525_token : boolean;
  signal place_1526_preds : BooleanArray(0 downto 0);
  signal place_1526_succs : BooleanArray(0 downto 0);
  signal place_1526_token : boolean;
  signal place_1527_preds : BooleanArray(0 downto 0);
  signal place_1527_succs : BooleanArray(0 downto 0);
  signal place_1527_token : boolean;
  signal place_1528_preds : BooleanArray(0 downto 0);
  signal place_1528_succs : BooleanArray(0 downto 0);
  signal place_1528_token : boolean;
  signal place_1529_preds : BooleanArray(0 downto 0);
  signal place_1529_succs : BooleanArray(0 downto 0);
  signal place_1529_token : boolean;
  signal place_1530_preds : BooleanArray(0 downto 0);
  signal place_1530_succs : BooleanArray(0 downto 0);
  signal place_1530_token : boolean;
  signal place_1531_preds : BooleanArray(0 downto 0);
  signal place_1531_succs : BooleanArray(0 downto 0);
  signal place_1531_token : boolean;
  signal place_1532_preds : BooleanArray(0 downto 0);
  signal place_1532_succs : BooleanArray(0 downto 0);
  signal place_1532_token : boolean;
  signal place_1533_preds : BooleanArray(0 downto 0);
  signal place_1533_succs : BooleanArray(0 downto 0);
  signal place_1533_token : boolean;
  signal place_1534_preds : BooleanArray(0 downto 0);
  signal place_1534_succs : BooleanArray(0 downto 0);
  signal place_1534_token : boolean;
  signal place_1535_preds : BooleanArray(0 downto 0);
  signal place_1535_succs : BooleanArray(0 downto 0);
  signal place_1535_token : boolean;
  signal place_1536_preds : BooleanArray(0 downto 0);
  signal place_1536_succs : BooleanArray(0 downto 0);
  signal place_1536_token : boolean;
  signal place_1537_preds : BooleanArray(0 downto 0);
  signal place_1537_succs : BooleanArray(0 downto 0);
  signal place_1537_token : boolean;
  signal place_1538_preds : BooleanArray(0 downto 0);
  signal place_1538_succs : BooleanArray(0 downto 0);
  signal place_1538_token : boolean;
  signal place_1539_preds : BooleanArray(0 downto 0);
  signal place_1539_succs : BooleanArray(0 downto 0);
  signal place_1539_token : boolean;
  signal place_1540_preds : BooleanArray(0 downto 0);
  signal place_1540_succs : BooleanArray(0 downto 0);
  signal place_1540_token : boolean;
  signal place_1541_preds : BooleanArray(0 downto 0);
  signal place_1541_succs : BooleanArray(0 downto 0);
  signal place_1541_token : boolean;
  signal place_1542_preds : BooleanArray(0 downto 0);
  signal place_1542_succs : BooleanArray(0 downto 0);
  signal place_1542_token : boolean;
  signal place_1543_preds : BooleanArray(0 downto 0);
  signal place_1543_succs : BooleanArray(0 downto 0);
  signal place_1543_token : boolean;
  signal place_1544_preds : BooleanArray(0 downto 0);
  signal place_1544_succs : BooleanArray(0 downto 0);
  signal place_1544_token : boolean;
  signal place_1545_preds : BooleanArray(0 downto 0);
  signal place_1545_succs : BooleanArray(0 downto 0);
  signal place_1545_token : boolean;
  signal place_1546_preds : BooleanArray(0 downto 0);
  signal place_1546_succs : BooleanArray(0 downto 0);
  signal place_1546_token : boolean;
  signal place_1547_preds : BooleanArray(0 downto 0);
  signal place_1547_succs : BooleanArray(0 downto 0);
  signal place_1547_token : boolean;
  signal place_1548_preds : BooleanArray(0 downto 0);
  signal place_1548_succs : BooleanArray(0 downto 0);
  signal place_1548_token : boolean;
  signal place_1549_preds : BooleanArray(0 downto 0);
  signal place_1549_succs : BooleanArray(0 downto 0);
  signal place_1549_token : boolean;
  signal place_1550_preds : BooleanArray(0 downto 0);
  signal place_1550_succs : BooleanArray(0 downto 0);
  signal place_1550_token : boolean;
  signal place_1551_preds : BooleanArray(0 downto 0);
  signal place_1551_succs : BooleanArray(0 downto 0);
  signal place_1551_token : boolean;
  signal place_1552_preds : BooleanArray(0 downto 0);
  signal place_1552_succs : BooleanArray(0 downto 0);
  signal place_1552_token : boolean;
  signal place_1553_preds : BooleanArray(0 downto 0);
  signal place_1553_succs : BooleanArray(0 downto 0);
  signal place_1553_token : boolean;

  signal transition_1_symbol_out : boolean;
  signal transition_1_preds : BooleanArray(0 downto 0);
  signal transition_2_symbol_out : boolean;
  signal transition_2_preds : BooleanArray(0 downto 0);
  signal transition_3_symbol_out : boolean;
  signal transition_3_preds : BooleanArray(0 downto 0);
  signal transition_4_symbol_out : boolean;
  signal transition_4_preds : BooleanArray(1 downto 0);
  signal transition_6_symbol_out : boolean;
  signal transition_6_preds : BooleanArray(0 downto 0);
  signal transition_7_symbol_out : boolean;
  signal transition_7_preds : BooleanArray(0 downto 0);
  signal transition_8_symbol_out : boolean;
  signal transition_8_preds : BooleanArray(0 downto 0);
  signal transition_9_symbol_out : boolean;
  signal transition_9_preds : BooleanArray(0 downto 0);
  signal transition_10_symbol_out : boolean;
  signal transition_10_preds : BooleanArray(0 downto 0);
  signal transition_11_symbol_out : boolean;
  signal transition_11_preds : BooleanArray(0 downto 0);
  signal transition_15_symbol_out : boolean;
  signal transition_15_preds : BooleanArray(0 downto 0);
  signal transition_16_symbol_out : boolean;
  signal transition_16_preds : BooleanArray(0 downto 0);
  signal transition_17_symbol_out : boolean;
  signal transition_17_preds : BooleanArray(0 downto 0);
  signal transition_18_symbol_out : boolean;
  signal transition_18_preds : BooleanArray(0 downto 0);
  signal transition_22_symbol_out : boolean;
  signal transition_22_preds : BooleanArray(0 downto 0);
  signal transition_23_symbol_out : boolean;
  signal transition_23_preds : BooleanArray(0 downto 0);
  signal transition_24_symbol_out : boolean;
  signal transition_24_preds : BooleanArray(0 downto 0);
  signal transition_25_symbol_out : boolean;
  signal transition_25_preds : BooleanArray(0 downto 0);
  signal transition_29_symbol_out : boolean;
  signal transition_29_preds : BooleanArray(1 downto 0);
  signal transition_30_symbol_out : boolean;
  signal transition_30_preds : BooleanArray(0 downto 0);
  signal transition_31_symbol_out : boolean;
  signal transition_31_preds : BooleanArray(0 downto 0);
  signal transition_32_symbol_out : boolean;
  signal transition_32_preds : BooleanArray(0 downto 0);
  signal transition_33_symbol_out : boolean;
  signal transition_33_preds : BooleanArray(0 downto 0);
  signal transition_37_symbol_out : boolean;
  signal transition_37_preds : BooleanArray(0 downto 0);
  signal transition_38_symbol_out : boolean;
  signal transition_38_preds : BooleanArray(0 downto 0);
  signal transition_39_symbol_out : boolean;
  signal transition_39_preds : BooleanArray(0 downto 0);
  signal transition_40_symbol_out : boolean;
  signal transition_40_preds : BooleanArray(0 downto 0);
  signal transition_44_symbol_out : boolean;
  signal transition_44_preds : BooleanArray(1 downto 0);
  signal transition_45_symbol_out : boolean;
  signal transition_45_preds : BooleanArray(0 downto 0);
  signal transition_46_symbol_out : boolean;
  signal transition_46_preds : BooleanArray(0 downto 0);
  signal transition_47_symbol_out : boolean;
  signal transition_47_preds : BooleanArray(0 downto 0);
  signal transition_48_symbol_out : boolean;
  signal transition_48_preds : BooleanArray(0 downto 0);
  signal transition_53_symbol_out : boolean;
  signal transition_53_preds : BooleanArray(0 downto 0);
  signal transition_54_symbol_out : boolean;
  signal transition_54_preds : BooleanArray(0 downto 0);
  signal transition_55_symbol_out : boolean;
  signal transition_55_preds : BooleanArray(1 downto 0);
  signal transition_57_symbol_out : boolean;
  signal transition_57_preds : BooleanArray(0 downto 0);
  signal transition_58_symbol_out : boolean;
  signal transition_58_preds : BooleanArray(0 downto 0);
  signal transition_59_symbol_out : boolean;
  signal transition_59_preds : BooleanArray(0 downto 0);
  signal transition_60_symbol_out : boolean;
  signal transition_60_preds : BooleanArray(0 downto 0);
  signal transition_61_symbol_out : boolean;
  signal transition_61_preds : BooleanArray(0 downto 0);
  signal transition_62_symbol_out : boolean;
  signal transition_62_preds : BooleanArray(0 downto 0);
  signal transition_63_symbol_out : boolean;
  signal transition_63_preds : BooleanArray(0 downto 0);
  signal transition_67_symbol_out : boolean;
  signal transition_67_preds : BooleanArray(0 downto 0);
  signal transition_68_symbol_out : boolean;
  signal transition_68_preds : BooleanArray(0 downto 0);
  signal transition_69_symbol_out : boolean;
  signal transition_69_preds : BooleanArray(0 downto 0);
  signal transition_70_symbol_out : boolean;
  signal transition_70_preds : BooleanArray(0 downto 0);
  signal transition_74_symbol_out : boolean;
  signal transition_74_preds : BooleanArray(0 downto 0);
  signal transition_75_symbol_out : boolean;
  signal transition_75_preds : BooleanArray(0 downto 0);
  signal transition_76_symbol_out : boolean;
  signal transition_76_preds : BooleanArray(0 downto 0);
  signal transition_77_symbol_out : boolean;
  signal transition_77_preds : BooleanArray(0 downto 0);
  signal transition_81_symbol_out : boolean;
  signal transition_81_preds : BooleanArray(1 downto 0);
  signal transition_82_symbol_out : boolean;
  signal transition_82_preds : BooleanArray(0 downto 0);
  signal transition_83_symbol_out : boolean;
  signal transition_83_preds : BooleanArray(0 downto 0);
  signal transition_84_symbol_out : boolean;
  signal transition_84_preds : BooleanArray(0 downto 0);
  signal transition_85_symbol_out : boolean;
  signal transition_85_preds : BooleanArray(0 downto 0);
  signal transition_89_symbol_out : boolean;
  signal transition_89_preds : BooleanArray(0 downto 0);
  signal transition_90_symbol_out : boolean;
  signal transition_90_preds : BooleanArray(0 downto 0);
  signal transition_91_symbol_out : boolean;
  signal transition_91_preds : BooleanArray(0 downto 0);
  signal transition_92_symbol_out : boolean;
  signal transition_92_preds : BooleanArray(0 downto 0);
  signal transition_96_symbol_out : boolean;
  signal transition_96_preds : BooleanArray(1 downto 0);
  signal transition_97_symbol_out : boolean;
  signal transition_97_preds : BooleanArray(0 downto 0);
  signal transition_98_symbol_out : boolean;
  signal transition_98_preds : BooleanArray(0 downto 0);
  signal transition_99_symbol_out : boolean;
  signal transition_99_preds : BooleanArray(0 downto 0);
  signal transition_100_symbol_out : boolean;
  signal transition_100_preds : BooleanArray(0 downto 0);
  signal transition_105_symbol_out : boolean;
  signal transition_105_preds : BooleanArray(0 downto 0);
  signal transition_106_symbol_out : boolean;
  signal transition_106_preds : BooleanArray(0 downto 0);
  signal transition_107_symbol_out : boolean;
  signal transition_107_preds : BooleanArray(1 downto 0);
  signal transition_109_symbol_out : boolean;
  signal transition_109_preds : BooleanArray(0 downto 0);
  signal transition_110_symbol_out : boolean;
  signal transition_110_preds : BooleanArray(0 downto 0);
  signal transition_111_symbol_out : boolean;
  signal transition_111_preds : BooleanArray(0 downto 0);
  signal transition_112_symbol_out : boolean;
  signal transition_112_preds : BooleanArray(0 downto 0);
  signal transition_113_symbol_out : boolean;
  signal transition_113_preds : BooleanArray(0 downto 0);
  signal transition_114_symbol_out : boolean;
  signal transition_114_preds : BooleanArray(0 downto 0);
  signal transition_115_symbol_out : boolean;
  signal transition_115_preds : BooleanArray(0 downto 0);
  signal transition_119_symbol_out : boolean;
  signal transition_119_preds : BooleanArray(1 downto 0);
  signal transition_120_symbol_out : boolean;
  signal transition_120_preds : BooleanArray(0 downto 0);
  signal transition_121_symbol_out : boolean;
  signal transition_121_preds : BooleanArray(0 downto 0);
  signal transition_122_symbol_out : boolean;
  signal transition_122_preds : BooleanArray(0 downto 0);
  signal transition_123_symbol_out : boolean;
  signal transition_123_preds : BooleanArray(0 downto 0);
  signal transition_124_symbol_out : boolean;
  signal transition_124_preds : BooleanArray(0 downto 0);
  signal transition_128_symbol_out : boolean;
  signal transition_128_preds : BooleanArray(0 downto 0);
  signal transition_129_symbol_out : boolean;
  signal transition_129_preds : BooleanArray(0 downto 0);
  signal transition_130_symbol_out : boolean;
  signal transition_130_preds : BooleanArray(0 downto 0);
  signal transition_131_symbol_out : boolean;
  signal transition_131_preds : BooleanArray(0 downto 0);
  signal transition_135_symbol_out : boolean;
  signal transition_135_preds : BooleanArray(0 downto 0);
  signal transition_136_symbol_out : boolean;
  signal transition_136_preds : BooleanArray(0 downto 0);
  signal transition_137_symbol_out : boolean;
  signal transition_137_preds : BooleanArray(0 downto 0);
  signal transition_138_symbol_out : boolean;
  signal transition_138_preds : BooleanArray(0 downto 0);
  signal transition_142_symbol_out : boolean;
  signal transition_142_preds : BooleanArray(1 downto 0);
  signal transition_143_symbol_out : boolean;
  signal transition_143_preds : BooleanArray(0 downto 0);
  signal transition_144_symbol_out : boolean;
  signal transition_144_preds : BooleanArray(0 downto 0);
  signal transition_145_symbol_out : boolean;
  signal transition_145_preds : BooleanArray(0 downto 0);
  signal transition_146_symbol_out : boolean;
  signal transition_146_preds : BooleanArray(0 downto 0);
  signal transition_150_symbol_out : boolean;
  signal transition_150_preds : BooleanArray(0 downto 0);
  signal transition_151_symbol_out : boolean;
  signal transition_151_preds : BooleanArray(0 downto 0);
  signal transition_152_symbol_out : boolean;
  signal transition_152_preds : BooleanArray(0 downto 0);
  signal transition_153_symbol_out : boolean;
  signal transition_153_preds : BooleanArray(0 downto 0);
  signal transition_157_symbol_out : boolean;
  signal transition_157_preds : BooleanArray(1 downto 0);
  signal transition_158_symbol_out : boolean;
  signal transition_158_preds : BooleanArray(0 downto 0);
  signal transition_159_symbol_out : boolean;
  signal transition_159_preds : BooleanArray(0 downto 0);
  signal transition_160_symbol_out : boolean;
  signal transition_160_preds : BooleanArray(0 downto 0);
  signal transition_161_symbol_out : boolean;
  signal transition_161_preds : BooleanArray(0 downto 0);
  signal transition_166_symbol_out : boolean;
  signal transition_166_preds : BooleanArray(0 downto 0);
  signal transition_167_symbol_out : boolean;
  signal transition_167_preds : BooleanArray(0 downto 0);
  signal transition_168_symbol_out : boolean;
  signal transition_168_preds : BooleanArray(1 downto 0);
  signal transition_169_symbol_out : boolean;
  signal transition_169_preds : BooleanArray(0 downto 0);
  signal transition_170_symbol_out : boolean;
  signal transition_170_preds : BooleanArray(0 downto 0);
  signal transition_171_symbol_out : boolean;
  signal transition_171_preds : BooleanArray(0 downto 0);
  signal transition_172_symbol_out : boolean;
  signal transition_172_preds : BooleanArray(0 downto 0);
  signal transition_173_symbol_out : boolean;
  signal transition_173_preds : BooleanArray(0 downto 0);
  signal transition_177_symbol_out : boolean;
  signal transition_177_preds : BooleanArray(0 downto 0);
  signal transition_178_symbol_out : boolean;
  signal transition_178_preds : BooleanArray(0 downto 0);
  signal transition_179_symbol_out : boolean;
  signal transition_179_preds : BooleanArray(0 downto 0);
  signal transition_180_symbol_out : boolean;
  signal transition_180_preds : BooleanArray(0 downto 0);
  signal transition_184_symbol_out : boolean;
  signal transition_184_preds : BooleanArray(0 downto 0);
  signal transition_185_symbol_out : boolean;
  signal transition_185_preds : BooleanArray(0 downto 0);
  signal transition_186_symbol_out : boolean;
  signal transition_186_preds : BooleanArray(0 downto 0);
  signal transition_187_symbol_out : boolean;
  signal transition_187_preds : BooleanArray(0 downto 0);
  signal transition_191_symbol_out : boolean;
  signal transition_191_preds : BooleanArray(1 downto 0);
  signal transition_192_symbol_out : boolean;
  signal transition_192_preds : BooleanArray(0 downto 0);
  signal transition_193_symbol_out : boolean;
  signal transition_193_preds : BooleanArray(0 downto 0);
  signal transition_194_symbol_out : boolean;
  signal transition_194_preds : BooleanArray(0 downto 0);
  signal transition_195_symbol_out : boolean;
  signal transition_195_preds : BooleanArray(0 downto 0);
  signal transition_199_symbol_out : boolean;
  signal transition_199_preds : BooleanArray(0 downto 0);
  signal transition_200_symbol_out : boolean;
  signal transition_200_preds : BooleanArray(0 downto 0);
  signal transition_201_symbol_out : boolean;
  signal transition_201_preds : BooleanArray(0 downto 0);
  signal transition_202_symbol_out : boolean;
  signal transition_202_preds : BooleanArray(0 downto 0);
  signal transition_206_symbol_out : boolean;
  signal transition_206_preds : BooleanArray(1 downto 0);
  signal transition_207_symbol_out : boolean;
  signal transition_207_preds : BooleanArray(0 downto 0);
  signal transition_208_symbol_out : boolean;
  signal transition_208_preds : BooleanArray(0 downto 0);
  signal transition_209_symbol_out : boolean;
  signal transition_209_preds : BooleanArray(0 downto 0);
  signal transition_210_symbol_out : boolean;
  signal transition_210_preds : BooleanArray(0 downto 0);
  signal transition_215_symbol_out : boolean;
  signal transition_215_preds : BooleanArray(0 downto 0);
  signal transition_216_symbol_out : boolean;
  signal transition_216_preds : BooleanArray(0 downto 0);
  signal transition_217_symbol_out : boolean;
  signal transition_217_preds : BooleanArray(1 downto 0);
  signal transition_219_symbol_out : boolean;
  signal transition_219_preds : BooleanArray(0 downto 0);
  signal transition_220_symbol_out : boolean;
  signal transition_220_preds : BooleanArray(0 downto 0);
  signal transition_221_symbol_out : boolean;
  signal transition_221_preds : BooleanArray(0 downto 0);
  signal transition_222_symbol_out : boolean;
  signal transition_222_preds : BooleanArray(0 downto 0);
  signal transition_223_symbol_out : boolean;
  signal transition_223_preds : BooleanArray(0 downto 0);
  signal transition_224_symbol_out : boolean;
  signal transition_224_preds : BooleanArray(0 downto 0);
  signal transition_225_symbol_out : boolean;
  signal transition_225_preds : BooleanArray(0 downto 0);
  signal transition_229_symbol_out : boolean;
  signal transition_229_preds : BooleanArray(0 downto 0);
  signal transition_230_symbol_out : boolean;
  signal transition_230_preds : BooleanArray(0 downto 0);
  signal transition_231_symbol_out : boolean;
  signal transition_231_preds : BooleanArray(0 downto 0);
  signal transition_232_symbol_out : boolean;
  signal transition_232_preds : BooleanArray(0 downto 0);
  signal transition_236_symbol_out : boolean;
  signal transition_236_preds : BooleanArray(0 downto 0);
  signal transition_237_symbol_out : boolean;
  signal transition_237_preds : BooleanArray(0 downto 0);
  signal transition_238_symbol_out : boolean;
  signal transition_238_preds : BooleanArray(0 downto 0);
  signal transition_239_symbol_out : boolean;
  signal transition_239_preds : BooleanArray(0 downto 0);
  signal transition_243_symbol_out : boolean;
  signal transition_243_preds : BooleanArray(1 downto 0);
  signal transition_244_symbol_out : boolean;
  signal transition_244_preds : BooleanArray(0 downto 0);
  signal transition_245_symbol_out : boolean;
  signal transition_245_preds : BooleanArray(0 downto 0);
  signal transition_246_symbol_out : boolean;
  signal transition_246_preds : BooleanArray(0 downto 0);
  signal transition_247_symbol_out : boolean;
  signal transition_247_preds : BooleanArray(0 downto 0);
  signal transition_251_symbol_out : boolean;
  signal transition_251_preds : BooleanArray(0 downto 0);
  signal transition_252_symbol_out : boolean;
  signal transition_252_preds : BooleanArray(0 downto 0);
  signal transition_253_symbol_out : boolean;
  signal transition_253_preds : BooleanArray(0 downto 0);
  signal transition_254_symbol_out : boolean;
  signal transition_254_preds : BooleanArray(0 downto 0);
  signal transition_258_symbol_out : boolean;
  signal transition_258_preds : BooleanArray(1 downto 0);
  signal transition_259_symbol_out : boolean;
  signal transition_259_preds : BooleanArray(0 downto 0);
  signal transition_260_symbol_out : boolean;
  signal transition_260_preds : BooleanArray(0 downto 0);
  signal transition_261_symbol_out : boolean;
  signal transition_261_preds : BooleanArray(0 downto 0);
  signal transition_262_symbol_out : boolean;
  signal transition_262_preds : BooleanArray(0 downto 0);
  signal transition_267_symbol_out : boolean;
  signal transition_267_preds : BooleanArray(0 downto 0);
  signal transition_268_symbol_out : boolean;
  signal transition_268_preds : BooleanArray(0 downto 0);
  signal transition_269_symbol_out : boolean;
  signal transition_269_preds : BooleanArray(1 downto 0);
  signal transition_271_symbol_out : boolean;
  signal transition_271_preds : BooleanArray(0 downto 0);
  signal transition_272_symbol_out : boolean;
  signal transition_272_preds : BooleanArray(0 downto 0);
  signal transition_273_symbol_out : boolean;
  signal transition_273_preds : BooleanArray(0 downto 0);
  signal transition_274_symbol_out : boolean;
  signal transition_274_preds : BooleanArray(0 downto 0);
  signal transition_275_symbol_out : boolean;
  signal transition_275_preds : BooleanArray(0 downto 0);
  signal transition_276_symbol_out : boolean;
  signal transition_276_preds : BooleanArray(0 downto 0);
  signal transition_277_symbol_out : boolean;
  signal transition_277_preds : BooleanArray(0 downto 0);
  signal transition_281_symbol_out : boolean;
  signal transition_281_preds : BooleanArray(1 downto 0);
  signal transition_282_symbol_out : boolean;
  signal transition_282_preds : BooleanArray(0 downto 0);
  signal transition_283_symbol_out : boolean;
  signal transition_283_preds : BooleanArray(0 downto 0);
  signal transition_284_symbol_out : boolean;
  signal transition_284_preds : BooleanArray(0 downto 0);
  signal transition_285_symbol_out : boolean;
  signal transition_285_preds : BooleanArray(0 downto 0);
  signal transition_286_symbol_out : boolean;
  signal transition_286_preds : BooleanArray(0 downto 0);
  signal transition_290_symbol_out : boolean;
  signal transition_290_preds : BooleanArray(0 downto 0);
  signal transition_291_symbol_out : boolean;
  signal transition_291_preds : BooleanArray(0 downto 0);
  signal transition_292_symbol_out : boolean;
  signal transition_292_preds : BooleanArray(0 downto 0);
  signal transition_293_symbol_out : boolean;
  signal transition_293_preds : BooleanArray(0 downto 0);
  signal transition_297_symbol_out : boolean;
  signal transition_297_preds : BooleanArray(0 downto 0);
  signal transition_298_symbol_out : boolean;
  signal transition_298_preds : BooleanArray(0 downto 0);
  signal transition_299_symbol_out : boolean;
  signal transition_299_preds : BooleanArray(0 downto 0);
  signal transition_300_symbol_out : boolean;
  signal transition_300_preds : BooleanArray(0 downto 0);
  signal transition_304_symbol_out : boolean;
  signal transition_304_preds : BooleanArray(1 downto 0);
  signal transition_305_symbol_out : boolean;
  signal transition_305_preds : BooleanArray(0 downto 0);
  signal transition_306_symbol_out : boolean;
  signal transition_306_preds : BooleanArray(0 downto 0);
  signal transition_307_symbol_out : boolean;
  signal transition_307_preds : BooleanArray(0 downto 0);
  signal transition_308_symbol_out : boolean;
  signal transition_308_preds : BooleanArray(0 downto 0);
  signal transition_312_symbol_out : boolean;
  signal transition_312_preds : BooleanArray(0 downto 0);
  signal transition_313_symbol_out : boolean;
  signal transition_313_preds : BooleanArray(0 downto 0);
  signal transition_314_symbol_out : boolean;
  signal transition_314_preds : BooleanArray(0 downto 0);
  signal transition_315_symbol_out : boolean;
  signal transition_315_preds : BooleanArray(0 downto 0);
  signal transition_319_symbol_out : boolean;
  signal transition_319_preds : BooleanArray(1 downto 0);
  signal transition_320_symbol_out : boolean;
  signal transition_320_preds : BooleanArray(0 downto 0);
  signal transition_321_symbol_out : boolean;
  signal transition_321_preds : BooleanArray(0 downto 0);
  signal transition_322_symbol_out : boolean;
  signal transition_322_preds : BooleanArray(0 downto 0);
  signal transition_323_symbol_out : boolean;
  signal transition_323_preds : BooleanArray(0 downto 0);
  signal transition_328_symbol_out : boolean;
  signal transition_328_preds : BooleanArray(0 downto 0);
  signal transition_329_symbol_out : boolean;
  signal transition_329_preds : BooleanArray(0 downto 0);
  signal transition_330_symbol_out : boolean;
  signal transition_330_preds : BooleanArray(1 downto 0);
  signal transition_331_symbol_out : boolean;
  signal transition_331_preds : BooleanArray(0 downto 0);
  signal transition_332_symbol_out : boolean;
  signal transition_332_preds : BooleanArray(0 downto 0);
  signal transition_333_symbol_out : boolean;
  signal transition_333_preds : BooleanArray(0 downto 0);
  signal transition_334_symbol_out : boolean;
  signal transition_334_preds : BooleanArray(0 downto 0);
  signal transition_335_symbol_out : boolean;
  signal transition_335_preds : BooleanArray(0 downto 0);
  signal transition_339_symbol_out : boolean;
  signal transition_339_preds : BooleanArray(0 downto 0);
  signal transition_340_symbol_out : boolean;
  signal transition_340_preds : BooleanArray(0 downto 0);
  signal transition_341_symbol_out : boolean;
  signal transition_341_preds : BooleanArray(0 downto 0);
  signal transition_342_symbol_out : boolean;
  signal transition_342_preds : BooleanArray(0 downto 0);
  signal transition_346_symbol_out : boolean;
  signal transition_346_preds : BooleanArray(0 downto 0);
  signal transition_347_symbol_out : boolean;
  signal transition_347_preds : BooleanArray(0 downto 0);
  signal transition_348_symbol_out : boolean;
  signal transition_348_preds : BooleanArray(0 downto 0);
  signal transition_349_symbol_out : boolean;
  signal transition_349_preds : BooleanArray(0 downto 0);
  signal transition_353_symbol_out : boolean;
  signal transition_353_preds : BooleanArray(1 downto 0);
  signal transition_354_symbol_out : boolean;
  signal transition_354_preds : BooleanArray(0 downto 0);
  signal transition_355_symbol_out : boolean;
  signal transition_355_preds : BooleanArray(0 downto 0);
  signal transition_356_symbol_out : boolean;
  signal transition_356_preds : BooleanArray(0 downto 0);
  signal transition_357_symbol_out : boolean;
  signal transition_357_preds : BooleanArray(0 downto 0);
  signal transition_361_symbol_out : boolean;
  signal transition_361_preds : BooleanArray(0 downto 0);
  signal transition_362_symbol_out : boolean;
  signal transition_362_preds : BooleanArray(0 downto 0);
  signal transition_363_symbol_out : boolean;
  signal transition_363_preds : BooleanArray(0 downto 0);
  signal transition_364_symbol_out : boolean;
  signal transition_364_preds : BooleanArray(0 downto 0);
  signal transition_368_symbol_out : boolean;
  signal transition_368_preds : BooleanArray(1 downto 0);
  signal transition_369_symbol_out : boolean;
  signal transition_369_preds : BooleanArray(0 downto 0);
  signal transition_370_symbol_out : boolean;
  signal transition_370_preds : BooleanArray(0 downto 0);
  signal transition_371_symbol_out : boolean;
  signal transition_371_preds : BooleanArray(0 downto 0);
  signal transition_372_symbol_out : boolean;
  signal transition_372_preds : BooleanArray(0 downto 0);
  signal transition_377_symbol_out : boolean;
  signal transition_377_preds : BooleanArray(0 downto 0);
  signal transition_378_symbol_out : boolean;
  signal transition_378_preds : BooleanArray(0 downto 0);
  signal transition_379_symbol_out : boolean;
  signal transition_379_preds : BooleanArray(1 downto 0);
  signal transition_381_symbol_out : boolean;
  signal transition_381_preds : BooleanArray(0 downto 0);
  signal transition_382_symbol_out : boolean;
  signal transition_382_preds : BooleanArray(0 downto 0);
  signal transition_383_symbol_out : boolean;
  signal transition_383_preds : BooleanArray(0 downto 0);
  signal transition_384_symbol_out : boolean;
  signal transition_384_preds : BooleanArray(0 downto 0);
  signal transition_385_symbol_out : boolean;
  signal transition_385_preds : BooleanArray(0 downto 0);
  signal transition_386_symbol_out : boolean;
  signal transition_386_preds : BooleanArray(0 downto 0);
  signal transition_387_symbol_out : boolean;
  signal transition_387_preds : BooleanArray(0 downto 0);
  signal transition_391_symbol_out : boolean;
  signal transition_391_preds : BooleanArray(0 downto 0);
  signal transition_392_symbol_out : boolean;
  signal transition_392_preds : BooleanArray(0 downto 0);
  signal transition_393_symbol_out : boolean;
  signal transition_393_preds : BooleanArray(0 downto 0);
  signal transition_394_symbol_out : boolean;
  signal transition_394_preds : BooleanArray(0 downto 0);
  signal transition_398_symbol_out : boolean;
  signal transition_398_preds : BooleanArray(0 downto 0);
  signal transition_399_symbol_out : boolean;
  signal transition_399_preds : BooleanArray(0 downto 0);
  signal transition_400_symbol_out : boolean;
  signal transition_400_preds : BooleanArray(0 downto 0);
  signal transition_401_symbol_out : boolean;
  signal transition_401_preds : BooleanArray(0 downto 0);
  signal transition_405_symbol_out : boolean;
  signal transition_405_preds : BooleanArray(1 downto 0);
  signal transition_406_symbol_out : boolean;
  signal transition_406_preds : BooleanArray(0 downto 0);
  signal transition_407_symbol_out : boolean;
  signal transition_407_preds : BooleanArray(0 downto 0);
  signal transition_408_symbol_out : boolean;
  signal transition_408_preds : BooleanArray(0 downto 0);
  signal transition_409_symbol_out : boolean;
  signal transition_409_preds : BooleanArray(0 downto 0);
  signal transition_413_symbol_out : boolean;
  signal transition_413_preds : BooleanArray(0 downto 0);
  signal transition_414_symbol_out : boolean;
  signal transition_414_preds : BooleanArray(0 downto 0);
  signal transition_415_symbol_out : boolean;
  signal transition_415_preds : BooleanArray(0 downto 0);
  signal transition_416_symbol_out : boolean;
  signal transition_416_preds : BooleanArray(0 downto 0);
  signal transition_420_symbol_out : boolean;
  signal transition_420_preds : BooleanArray(1 downto 0);
  signal transition_421_symbol_out : boolean;
  signal transition_421_preds : BooleanArray(0 downto 0);
  signal transition_422_symbol_out : boolean;
  signal transition_422_preds : BooleanArray(0 downto 0);
  signal transition_423_symbol_out : boolean;
  signal transition_423_preds : BooleanArray(0 downto 0);
  signal transition_424_symbol_out : boolean;
  signal transition_424_preds : BooleanArray(0 downto 0);
  signal transition_429_symbol_out : boolean;
  signal transition_429_preds : BooleanArray(0 downto 0);
  signal transition_430_symbol_out : boolean;
  signal transition_430_preds : BooleanArray(0 downto 0);
  signal transition_431_symbol_out : boolean;
  signal transition_431_preds : BooleanArray(1 downto 0);
  signal transition_433_symbol_out : boolean;
  signal transition_433_preds : BooleanArray(0 downto 0);
  signal transition_434_symbol_out : boolean;
  signal transition_434_preds : BooleanArray(0 downto 0);
  signal transition_435_symbol_out : boolean;
  signal transition_435_preds : BooleanArray(0 downto 0);
  signal transition_436_symbol_out : boolean;
  signal transition_436_preds : BooleanArray(0 downto 0);
  signal transition_437_symbol_out : boolean;
  signal transition_437_preds : BooleanArray(0 downto 0);
  signal transition_438_symbol_out : boolean;
  signal transition_438_preds : BooleanArray(0 downto 0);
  signal transition_439_symbol_out : boolean;
  signal transition_439_preds : BooleanArray(0 downto 0);
  signal transition_443_symbol_out : boolean;
  signal transition_443_preds : BooleanArray(1 downto 0);
  signal transition_444_symbol_out : boolean;
  signal transition_444_preds : BooleanArray(0 downto 0);
  signal transition_445_symbol_out : boolean;
  signal transition_445_preds : BooleanArray(0 downto 0);
  signal transition_446_symbol_out : boolean;
  signal transition_446_preds : BooleanArray(0 downto 0);
  signal transition_447_symbol_out : boolean;
  signal transition_447_preds : BooleanArray(0 downto 0);
  signal transition_448_symbol_out : boolean;
  signal transition_448_preds : BooleanArray(0 downto 0);
  signal transition_452_symbol_out : boolean;
  signal transition_452_preds : BooleanArray(0 downto 0);
  signal transition_453_symbol_out : boolean;
  signal transition_453_preds : BooleanArray(0 downto 0);
  signal transition_454_symbol_out : boolean;
  signal transition_454_preds : BooleanArray(0 downto 0);
  signal transition_455_symbol_out : boolean;
  signal transition_455_preds : BooleanArray(0 downto 0);
  signal transition_459_symbol_out : boolean;
  signal transition_459_preds : BooleanArray(0 downto 0);
  signal transition_460_symbol_out : boolean;
  signal transition_460_preds : BooleanArray(0 downto 0);
  signal transition_461_symbol_out : boolean;
  signal transition_461_preds : BooleanArray(0 downto 0);
  signal transition_462_symbol_out : boolean;
  signal transition_462_preds : BooleanArray(0 downto 0);
  signal transition_466_symbol_out : boolean;
  signal transition_466_preds : BooleanArray(1 downto 0);
  signal transition_467_symbol_out : boolean;
  signal transition_467_preds : BooleanArray(0 downto 0);
  signal transition_468_symbol_out : boolean;
  signal transition_468_preds : BooleanArray(0 downto 0);
  signal transition_469_symbol_out : boolean;
  signal transition_469_preds : BooleanArray(0 downto 0);
  signal transition_470_symbol_out : boolean;
  signal transition_470_preds : BooleanArray(0 downto 0);
  signal transition_474_symbol_out : boolean;
  signal transition_474_preds : BooleanArray(0 downto 0);
  signal transition_475_symbol_out : boolean;
  signal transition_475_preds : BooleanArray(0 downto 0);
  signal transition_476_symbol_out : boolean;
  signal transition_476_preds : BooleanArray(0 downto 0);
  signal transition_477_symbol_out : boolean;
  signal transition_477_preds : BooleanArray(0 downto 0);
  signal transition_481_symbol_out : boolean;
  signal transition_481_preds : BooleanArray(1 downto 0);
  signal transition_482_symbol_out : boolean;
  signal transition_482_preds : BooleanArray(0 downto 0);
  signal transition_483_symbol_out : boolean;
  signal transition_483_preds : BooleanArray(0 downto 0);
  signal transition_484_symbol_out : boolean;
  signal transition_484_preds : BooleanArray(0 downto 0);
  signal transition_485_symbol_out : boolean;
  signal transition_485_preds : BooleanArray(0 downto 0);
  signal transition_490_symbol_out : boolean;
  signal transition_490_preds : BooleanArray(0 downto 0);
  signal transition_491_symbol_out : boolean;
  signal transition_491_preds : BooleanArray(0 downto 0);
  signal transition_492_symbol_out : boolean;
  signal transition_492_preds : BooleanArray(1 downto 0);
  signal transition_493_symbol_out : boolean;
  signal transition_493_preds : BooleanArray(0 downto 0);
  signal transition_494_symbol_out : boolean;
  signal transition_494_preds : BooleanArray(0 downto 0);
  signal transition_495_symbol_out : boolean;
  signal transition_495_preds : BooleanArray(0 downto 0);
  signal transition_496_symbol_out : boolean;
  signal transition_496_preds : BooleanArray(0 downto 0);
  signal transition_500_symbol_out : boolean;
  signal transition_500_preds : BooleanArray(1 downto 0);
  signal transition_501_symbol_out : boolean;
  signal transition_501_preds : BooleanArray(0 downto 0);
  signal transition_502_symbol_out : boolean;
  signal transition_502_preds : BooleanArray(0 downto 0);
  signal transition_503_symbol_out : boolean;
  signal transition_503_preds : BooleanArray(0 downto 0);
  signal transition_504_symbol_out : boolean;
  signal transition_504_preds : BooleanArray(0 downto 0);
  signal transition_508_symbol_out : boolean;
  signal transition_508_preds : BooleanArray(0 downto 0);
  signal transition_509_symbol_out : boolean;
  signal transition_509_preds : BooleanArray(0 downto 0);
  signal transition_510_symbol_out : boolean;
  signal transition_510_preds : BooleanArray(0 downto 0);
  signal transition_511_symbol_out : boolean;
  signal transition_511_preds : BooleanArray(0 downto 0);
  signal transition_515_symbol_out : boolean;
  signal transition_515_preds : BooleanArray(0 downto 0);
  signal transition_516_symbol_out : boolean;
  signal transition_516_preds : BooleanArray(0 downto 0);
  signal transition_517_symbol_out : boolean;
  signal transition_517_preds : BooleanArray(0 downto 0);
  signal transition_518_symbol_out : boolean;
  signal transition_518_preds : BooleanArray(0 downto 0);
  signal transition_522_symbol_out : boolean;
  signal transition_522_preds : BooleanArray(0 downto 0);
  signal transition_523_symbol_out : boolean;
  signal transition_523_preds : BooleanArray(0 downto 0);
  signal transition_524_symbol_out : boolean;
  signal transition_524_preds : BooleanArray(0 downto 0);
  signal transition_525_symbol_out : boolean;
  signal transition_525_preds : BooleanArray(0 downto 0);
  signal transition_529_symbol_out : boolean;
  signal transition_529_preds : BooleanArray(1 downto 0);
  signal transition_530_symbol_out : boolean;
  signal transition_530_preds : BooleanArray(0 downto 0);
  signal transition_531_symbol_out : boolean;
  signal transition_531_preds : BooleanArray(0 downto 0);
  signal transition_532_symbol_out : boolean;
  signal transition_532_preds : BooleanArray(0 downto 0);
  signal transition_533_symbol_out : boolean;
  signal transition_533_preds : BooleanArray(0 downto 0);
  signal transition_537_symbol_out : boolean;
  signal transition_537_preds : BooleanArray(0 downto 0);
  signal transition_538_symbol_out : boolean;
  signal transition_538_preds : BooleanArray(0 downto 0);
  signal transition_539_symbol_out : boolean;
  signal transition_539_preds : BooleanArray(0 downto 0);
  signal transition_540_symbol_out : boolean;
  signal transition_540_preds : BooleanArray(0 downto 0);
  signal transition_544_symbol_out : boolean;
  signal transition_544_preds : BooleanArray(1 downto 0);
  signal transition_545_symbol_out : boolean;
  signal transition_545_preds : BooleanArray(0 downto 0);
  signal transition_546_symbol_out : boolean;
  signal transition_546_preds : BooleanArray(0 downto 0);
  signal transition_547_symbol_out : boolean;
  signal transition_547_preds : BooleanArray(0 downto 0);
  signal transition_548_symbol_out : boolean;
  signal transition_548_preds : BooleanArray(0 downto 0);
  signal transition_553_symbol_out : boolean;
  signal transition_553_preds : BooleanArray(0 downto 0);
  signal transition_554_symbol_out : boolean;
  signal transition_554_preds : BooleanArray(0 downto 0);
  signal transition_555_symbol_out : boolean;
  signal transition_555_preds : BooleanArray(2 downto 0);
  signal transition_556_symbol_out : boolean;
  signal transition_556_preds : BooleanArray(0 downto 0);
  signal transition_557_symbol_out : boolean;
  signal transition_557_preds : BooleanArray(0 downto 0);
  signal transition_558_symbol_out : boolean;
  signal transition_558_preds : BooleanArray(0 downto 0);
  signal transition_559_symbol_out : boolean;
  signal transition_559_preds : BooleanArray(0 downto 0);
  signal transition_563_symbol_out : boolean;
  signal transition_563_preds : BooleanArray(1 downto 0);
  signal transition_564_symbol_out : boolean;
  signal transition_564_preds : BooleanArray(0 downto 0);
  signal transition_565_symbol_out : boolean;
  signal transition_565_preds : BooleanArray(0 downto 0);
  signal transition_566_symbol_out : boolean;
  signal transition_566_preds : BooleanArray(0 downto 0);
  signal transition_567_symbol_out : boolean;
  signal transition_567_preds : BooleanArray(0 downto 0);
  signal transition_571_symbol_out : boolean;
  signal transition_571_preds : BooleanArray(0 downto 0);
  signal transition_572_symbol_out : boolean;
  signal transition_572_preds : BooleanArray(0 downto 0);
  signal transition_573_symbol_out : boolean;
  signal transition_573_preds : BooleanArray(0 downto 0);
  signal transition_574_symbol_out : boolean;
  signal transition_574_preds : BooleanArray(0 downto 0);
  signal transition_578_symbol_out : boolean;
  signal transition_578_preds : BooleanArray(0 downto 0);
  signal transition_579_symbol_out : boolean;
  signal transition_579_preds : BooleanArray(0 downto 0);
  signal transition_580_symbol_out : boolean;
  signal transition_580_preds : BooleanArray(0 downto 0);
  signal transition_581_symbol_out : boolean;
  signal transition_581_preds : BooleanArray(0 downto 0);
  signal transition_585_symbol_out : boolean;
  signal transition_585_preds : BooleanArray(0 downto 0);
  signal transition_586_symbol_out : boolean;
  signal transition_586_preds : BooleanArray(0 downto 0);
  signal transition_587_symbol_out : boolean;
  signal transition_587_preds : BooleanArray(0 downto 0);
  signal transition_588_symbol_out : boolean;
  signal transition_588_preds : BooleanArray(0 downto 0);
  signal transition_592_symbol_out : boolean;
  signal transition_592_preds : BooleanArray(1 downto 0);
  signal transition_593_symbol_out : boolean;
  signal transition_593_preds : BooleanArray(0 downto 0);
  signal transition_594_symbol_out : boolean;
  signal transition_594_preds : BooleanArray(0 downto 0);
  signal transition_595_symbol_out : boolean;
  signal transition_595_preds : BooleanArray(0 downto 0);
  signal transition_596_symbol_out : boolean;
  signal transition_596_preds : BooleanArray(0 downto 0);
  signal transition_600_symbol_out : boolean;
  signal transition_600_preds : BooleanArray(0 downto 0);
  signal transition_601_symbol_out : boolean;
  signal transition_601_preds : BooleanArray(0 downto 0);
  signal transition_602_symbol_out : boolean;
  signal transition_602_preds : BooleanArray(0 downto 0);
  signal transition_603_symbol_out : boolean;
  signal transition_603_preds : BooleanArray(0 downto 0);
  signal transition_607_symbol_out : boolean;
  signal transition_607_preds : BooleanArray(1 downto 0);
  signal transition_608_symbol_out : boolean;
  signal transition_608_preds : BooleanArray(0 downto 0);
  signal transition_609_symbol_out : boolean;
  signal transition_609_preds : BooleanArray(0 downto 0);
  signal transition_610_symbol_out : boolean;
  signal transition_610_preds : BooleanArray(0 downto 0);
  signal transition_611_symbol_out : boolean;
  signal transition_611_preds : BooleanArray(0 downto 0);
  signal transition_616_symbol_out : boolean;
  signal transition_616_preds : BooleanArray(0 downto 0);
  signal transition_617_symbol_out : boolean;
  signal transition_617_preds : BooleanArray(0 downto 0);
  signal transition_618_symbol_out : boolean;
  signal transition_618_preds : BooleanArray(2 downto 0);
  signal transition_619_symbol_out : boolean;
  signal transition_619_preds : BooleanArray(0 downto 0);
  signal transition_620_symbol_out : boolean;
  signal transition_620_preds : BooleanArray(0 downto 0);
  signal transition_621_symbol_out : boolean;
  signal transition_621_preds : BooleanArray(0 downto 0);
  signal transition_622_symbol_out : boolean;
  signal transition_622_preds : BooleanArray(0 downto 0);
  signal transition_626_symbol_out : boolean;
  signal transition_626_preds : BooleanArray(1 downto 0);
  signal transition_627_symbol_out : boolean;
  signal transition_627_preds : BooleanArray(0 downto 0);
  signal transition_628_symbol_out : boolean;
  signal transition_628_preds : BooleanArray(0 downto 0);
  signal transition_629_symbol_out : boolean;
  signal transition_629_preds : BooleanArray(0 downto 0);
  signal transition_630_symbol_out : boolean;
  signal transition_630_preds : BooleanArray(0 downto 0);
  signal transition_634_symbol_out : boolean;
  signal transition_634_preds : BooleanArray(0 downto 0);
  signal transition_635_symbol_out : boolean;
  signal transition_635_preds : BooleanArray(0 downto 0);
  signal transition_636_symbol_out : boolean;
  signal transition_636_preds : BooleanArray(0 downto 0);
  signal transition_637_symbol_out : boolean;
  signal transition_637_preds : BooleanArray(0 downto 0);
  signal transition_641_symbol_out : boolean;
  signal transition_641_preds : BooleanArray(0 downto 0);
  signal transition_642_symbol_out : boolean;
  signal transition_642_preds : BooleanArray(0 downto 0);
  signal transition_643_symbol_out : boolean;
  signal transition_643_preds : BooleanArray(0 downto 0);
  signal transition_644_symbol_out : boolean;
  signal transition_644_preds : BooleanArray(0 downto 0);
  signal transition_648_symbol_out : boolean;
  signal transition_648_preds : BooleanArray(0 downto 0);
  signal transition_649_symbol_out : boolean;
  signal transition_649_preds : BooleanArray(0 downto 0);
  signal transition_650_symbol_out : boolean;
  signal transition_650_preds : BooleanArray(0 downto 0);
  signal transition_651_symbol_out : boolean;
  signal transition_651_preds : BooleanArray(0 downto 0);
  signal transition_655_symbol_out : boolean;
  signal transition_655_preds : BooleanArray(1 downto 0);
  signal transition_656_symbol_out : boolean;
  signal transition_656_preds : BooleanArray(0 downto 0);
  signal transition_657_symbol_out : boolean;
  signal transition_657_preds : BooleanArray(0 downto 0);
  signal transition_658_symbol_out : boolean;
  signal transition_658_preds : BooleanArray(0 downto 0);
  signal transition_659_symbol_out : boolean;
  signal transition_659_preds : BooleanArray(0 downto 0);
  signal transition_663_symbol_out : boolean;
  signal transition_663_preds : BooleanArray(0 downto 0);
  signal transition_664_symbol_out : boolean;
  signal transition_664_preds : BooleanArray(0 downto 0);
  signal transition_665_symbol_out : boolean;
  signal transition_665_preds : BooleanArray(0 downto 0);
  signal transition_666_symbol_out : boolean;
  signal transition_666_preds : BooleanArray(0 downto 0);
  signal transition_670_symbol_out : boolean;
  signal transition_670_preds : BooleanArray(1 downto 0);
  signal transition_671_symbol_out : boolean;
  signal transition_671_preds : BooleanArray(0 downto 0);
  signal transition_672_symbol_out : boolean;
  signal transition_672_preds : BooleanArray(0 downto 0);
  signal transition_673_symbol_out : boolean;
  signal transition_673_preds : BooleanArray(0 downto 0);
  signal transition_674_symbol_out : boolean;
  signal transition_674_preds : BooleanArray(0 downto 0);
  signal transition_679_symbol_out : boolean;
  signal transition_679_preds : BooleanArray(0 downto 0);
  signal transition_680_symbol_out : boolean;
  signal transition_680_preds : BooleanArray(0 downto 0);
  signal transition_681_symbol_out : boolean;
  signal transition_681_preds : BooleanArray(2 downto 0);
  signal transition_682_symbol_out : boolean;
  signal transition_682_preds : BooleanArray(0 downto 0);
  signal transition_683_symbol_out : boolean;
  signal transition_683_preds : BooleanArray(0 downto 0);
  signal transition_684_symbol_out : boolean;
  signal transition_684_preds : BooleanArray(0 downto 0);
  signal transition_685_symbol_out : boolean;
  signal transition_685_preds : BooleanArray(0 downto 0);
  signal transition_686_symbol_out : boolean;
  signal transition_686_preds : BooleanArray(0 downto 0);
  signal transition_690_symbol_out : boolean;
  signal transition_690_preds : BooleanArray(0 downto 0);
  signal transition_691_symbol_out : boolean;
  signal transition_691_preds : BooleanArray(0 downto 0);
  signal transition_692_symbol_out : boolean;
  signal transition_692_preds : BooleanArray(0 downto 0);
  signal transition_693_symbol_out : boolean;
  signal transition_693_preds : BooleanArray(0 downto 0);
  signal transition_697_symbol_out : boolean;
  signal transition_697_preds : BooleanArray(0 downto 0);
  signal transition_698_symbol_out : boolean;
  signal transition_698_preds : BooleanArray(0 downto 0);
  signal transition_699_symbol_out : boolean;
  signal transition_699_preds : BooleanArray(0 downto 0);
  signal transition_700_symbol_out : boolean;
  signal transition_700_preds : BooleanArray(0 downto 0);
  signal transition_704_symbol_out : boolean;
  signal transition_704_preds : BooleanArray(1 downto 0);
  signal transition_705_symbol_out : boolean;
  signal transition_705_preds : BooleanArray(0 downto 0);
  signal transition_706_symbol_out : boolean;
  signal transition_706_preds : BooleanArray(0 downto 0);
  signal transition_707_symbol_out : boolean;
  signal transition_707_preds : BooleanArray(0 downto 0);
  signal transition_708_symbol_out : boolean;
  signal transition_708_preds : BooleanArray(0 downto 0);
  signal transition_712_symbol_out : boolean;
  signal transition_712_preds : BooleanArray(0 downto 0);
  signal transition_713_symbol_out : boolean;
  signal transition_713_preds : BooleanArray(0 downto 0);
  signal transition_714_symbol_out : boolean;
  signal transition_714_preds : BooleanArray(0 downto 0);
  signal transition_715_symbol_out : boolean;
  signal transition_715_preds : BooleanArray(0 downto 0);
  signal transition_719_symbol_out : boolean;
  signal transition_719_preds : BooleanArray(1 downto 0);
  signal transition_720_symbol_out : boolean;
  signal transition_720_preds : BooleanArray(0 downto 0);
  signal transition_721_symbol_out : boolean;
  signal transition_721_preds : BooleanArray(0 downto 0);
  signal transition_722_symbol_out : boolean;
  signal transition_722_preds : BooleanArray(0 downto 0);
  signal transition_723_symbol_out : boolean;
  signal transition_723_preds : BooleanArray(0 downto 0);
  signal transition_728_symbol_out : boolean;
  signal transition_728_preds : BooleanArray(0 downto 0);
  signal transition_729_symbol_out : boolean;
  signal transition_729_preds : BooleanArray(0 downto 0);
  signal transition_730_symbol_out : boolean;
  signal transition_730_preds : BooleanArray(1 downto 0);
  signal transition_732_symbol_out : boolean;
  signal transition_732_preds : BooleanArray(0 downto 0);
  signal transition_733_symbol_out : boolean;
  signal transition_733_preds : BooleanArray(0 downto 0);
  signal transition_734_symbol_out : boolean;
  signal transition_734_preds : BooleanArray(0 downto 0);
  signal transition_735_symbol_out : boolean;
  signal transition_735_preds : BooleanArray(0 downto 0);
  signal transition_736_symbol_out : boolean;
  signal transition_736_preds : BooleanArray(0 downto 0);
  signal transition_737_symbol_out : boolean;
  signal transition_737_preds : BooleanArray(0 downto 0);
  signal transition_741_symbol_out : boolean;
  signal transition_741_preds : BooleanArray(0 downto 0);
  signal transition_742_symbol_out : boolean;
  signal transition_742_preds : BooleanArray(0 downto 0);
  signal transition_743_symbol_out : boolean;
  signal transition_743_preds : BooleanArray(0 downto 0);
  signal transition_744_symbol_out : boolean;
  signal transition_744_preds : BooleanArray(0 downto 0);
  signal transition_748_symbol_out : boolean;
  signal transition_748_preds : BooleanArray(0 downto 0);
  signal transition_749_symbol_out : boolean;
  signal transition_749_preds : BooleanArray(0 downto 0);
  signal transition_750_symbol_out : boolean;
  signal transition_750_preds : BooleanArray(0 downto 0);
  signal transition_751_symbol_out : boolean;
  signal transition_751_preds : BooleanArray(0 downto 0);
  signal transition_755_symbol_out : boolean;
  signal transition_755_preds : BooleanArray(1 downto 0);
  signal transition_756_symbol_out : boolean;
  signal transition_756_preds : BooleanArray(0 downto 0);
  signal transition_757_symbol_out : boolean;
  signal transition_757_preds : BooleanArray(0 downto 0);
  signal transition_758_symbol_out : boolean;
  signal transition_758_preds : BooleanArray(0 downto 0);
  signal transition_759_symbol_out : boolean;
  signal transition_759_preds : BooleanArray(0 downto 0);
  signal transition_763_symbol_out : boolean;
  signal transition_763_preds : BooleanArray(0 downto 0);
  signal transition_764_symbol_out : boolean;
  signal transition_764_preds : BooleanArray(0 downto 0);
  signal transition_765_symbol_out : boolean;
  signal transition_765_preds : BooleanArray(0 downto 0);
  signal transition_766_symbol_out : boolean;
  signal transition_766_preds : BooleanArray(0 downto 0);
  signal transition_770_symbol_out : boolean;
  signal transition_770_preds : BooleanArray(1 downto 0);
  signal transition_771_symbol_out : boolean;
  signal transition_771_preds : BooleanArray(0 downto 0);
  signal transition_772_symbol_out : boolean;
  signal transition_772_preds : BooleanArray(0 downto 0);
  signal transition_773_symbol_out : boolean;
  signal transition_773_preds : BooleanArray(0 downto 0);
  signal transition_774_symbol_out : boolean;
  signal transition_774_preds : BooleanArray(0 downto 0);
  signal transition_779_symbol_out : boolean;
  signal transition_779_preds : BooleanArray(0 downto 0);
  signal transition_780_symbol_out : boolean;
  signal transition_780_preds : BooleanArray(0 downto 0);
  signal transition_781_symbol_out : boolean;
  signal transition_781_preds : BooleanArray(1 downto 0);
  signal transition_783_symbol_out : boolean;
  signal transition_783_preds : BooleanArray(0 downto 0);
  signal transition_784_symbol_out : boolean;
  signal transition_784_preds : BooleanArray(0 downto 0);
  signal transition_785_symbol_out : boolean;
  signal transition_785_preds : BooleanArray(0 downto 0);
  signal transition_786_symbol_out : boolean;
  signal transition_786_preds : BooleanArray(0 downto 0);
  signal transition_787_symbol_out : boolean;
  signal transition_787_preds : BooleanArray(0 downto 0);
  signal transition_788_symbol_out : boolean;
  signal transition_788_preds : BooleanArray(0 downto 0);
  signal transition_792_symbol_out : boolean;
  signal transition_792_preds : BooleanArray(1 downto 0);
  signal transition_793_symbol_out : boolean;
  signal transition_793_preds : BooleanArray(0 downto 0);
  signal transition_794_symbol_out : boolean;
  signal transition_794_preds : BooleanArray(0 downto 0);
  signal transition_795_symbol_out : boolean;
  signal transition_795_preds : BooleanArray(0 downto 0);
  signal transition_796_symbol_out : boolean;
  signal transition_796_preds : BooleanArray(0 downto 0);
  signal transition_800_symbol_out : boolean;
  signal transition_800_preds : BooleanArray(0 downto 0);
  signal transition_801_symbol_out : boolean;
  signal transition_801_preds : BooleanArray(0 downto 0);
  signal transition_802_symbol_out : boolean;
  signal transition_802_preds : BooleanArray(0 downto 0);
  signal transition_803_symbol_out : boolean;
  signal transition_803_preds : BooleanArray(0 downto 0);
  signal transition_807_symbol_out : boolean;
  signal transition_807_preds : BooleanArray(0 downto 0);
  signal transition_808_symbol_out : boolean;
  signal transition_808_preds : BooleanArray(0 downto 0);
  signal transition_809_symbol_out : boolean;
  signal transition_809_preds : BooleanArray(0 downto 0);
  signal transition_810_symbol_out : boolean;
  signal transition_810_preds : BooleanArray(0 downto 0);
  signal transition_814_symbol_out : boolean;
  signal transition_814_preds : BooleanArray(0 downto 0);
  signal transition_815_symbol_out : boolean;
  signal transition_815_preds : BooleanArray(0 downto 0);
  signal transition_816_symbol_out : boolean;
  signal transition_816_preds : BooleanArray(0 downto 0);
  signal transition_817_symbol_out : boolean;
  signal transition_817_preds : BooleanArray(0 downto 0);
  signal transition_821_symbol_out : boolean;
  signal transition_821_preds : BooleanArray(1 downto 0);
  signal transition_822_symbol_out : boolean;
  signal transition_822_preds : BooleanArray(0 downto 0);
  signal transition_823_symbol_out : boolean;
  signal transition_823_preds : BooleanArray(0 downto 0);
  signal transition_824_symbol_out : boolean;
  signal transition_824_preds : BooleanArray(0 downto 0);
  signal transition_825_symbol_out : boolean;
  signal transition_825_preds : BooleanArray(0 downto 0);
  signal transition_829_symbol_out : boolean;
  signal transition_829_preds : BooleanArray(0 downto 0);
  signal transition_830_symbol_out : boolean;
  signal transition_830_preds : BooleanArray(0 downto 0);
  signal transition_831_symbol_out : boolean;
  signal transition_831_preds : BooleanArray(0 downto 0);
  signal transition_832_symbol_out : boolean;
  signal transition_832_preds : BooleanArray(0 downto 0);
  signal transition_836_symbol_out : boolean;
  signal transition_836_preds : BooleanArray(1 downto 0);
  signal transition_837_symbol_out : boolean;
  signal transition_837_preds : BooleanArray(0 downto 0);
  signal transition_838_symbol_out : boolean;
  signal transition_838_preds : BooleanArray(0 downto 0);
  signal transition_839_symbol_out : boolean;
  signal transition_839_preds : BooleanArray(0 downto 0);
  signal transition_840_symbol_out : boolean;
  signal transition_840_preds : BooleanArray(0 downto 0);
  signal transition_845_symbol_out : boolean;
  signal transition_845_preds : BooleanArray(0 downto 0);
  signal transition_846_symbol_out : boolean;
  signal transition_846_preds : BooleanArray(0 downto 0);
  signal transition_847_symbol_out : boolean;
  signal transition_847_preds : BooleanArray(1 downto 0);
  signal transition_848_symbol_out : boolean;
  signal transition_848_preds : BooleanArray(0 downto 0);
  signal transition_849_symbol_out : boolean;
  signal transition_849_preds : BooleanArray(0 downto 0);
  signal transition_850_symbol_out : boolean;
  signal transition_850_preds : BooleanArray(0 downto 0);
  signal transition_851_symbol_out : boolean;
  signal transition_851_preds : BooleanArray(0 downto 0);
  signal transition_852_symbol_out : boolean;
  signal transition_852_preds : BooleanArray(0 downto 0);
  signal transition_856_symbol_out : boolean;
  signal transition_856_preds : BooleanArray(0 downto 0);
  signal transition_857_symbol_out : boolean;
  signal transition_857_preds : BooleanArray(0 downto 0);
  signal transition_858_symbol_out : boolean;
  signal transition_858_preds : BooleanArray(0 downto 0);
  signal transition_859_symbol_out : boolean;
  signal transition_859_preds : BooleanArray(0 downto 0);
  signal transition_863_symbol_out : boolean;
  signal transition_863_preds : BooleanArray(0 downto 0);
  signal transition_864_symbol_out : boolean;
  signal transition_864_preds : BooleanArray(0 downto 0);
  signal transition_865_symbol_out : boolean;
  signal transition_865_preds : BooleanArray(0 downto 0);
  signal transition_866_symbol_out : boolean;
  signal transition_866_preds : BooleanArray(0 downto 0);
  signal transition_870_symbol_out : boolean;
  signal transition_870_preds : BooleanArray(1 downto 0);
  signal transition_871_symbol_out : boolean;
  signal transition_871_preds : BooleanArray(0 downto 0);
  signal transition_872_symbol_out : boolean;
  signal transition_872_preds : BooleanArray(0 downto 0);
  signal transition_873_symbol_out : boolean;
  signal transition_873_preds : BooleanArray(0 downto 0);
  signal transition_874_symbol_out : boolean;
  signal transition_874_preds : BooleanArray(0 downto 0);
  signal transition_878_symbol_out : boolean;
  signal transition_878_preds : BooleanArray(0 downto 0);
  signal transition_879_symbol_out : boolean;
  signal transition_879_preds : BooleanArray(0 downto 0);
  signal transition_880_symbol_out : boolean;
  signal transition_880_preds : BooleanArray(0 downto 0);
  signal transition_881_symbol_out : boolean;
  signal transition_881_preds : BooleanArray(0 downto 0);
  signal transition_885_symbol_out : boolean;
  signal transition_885_preds : BooleanArray(1 downto 0);
  signal transition_886_symbol_out : boolean;
  signal transition_886_preds : BooleanArray(0 downto 0);
  signal transition_887_symbol_out : boolean;
  signal transition_887_preds : BooleanArray(0 downto 0);
  signal transition_888_symbol_out : boolean;
  signal transition_888_preds : BooleanArray(0 downto 0);
  signal transition_889_symbol_out : boolean;
  signal transition_889_preds : BooleanArray(0 downto 0);
  signal transition_894_symbol_out : boolean;
  signal transition_894_preds : BooleanArray(0 downto 0);
  signal transition_895_symbol_out : boolean;
  signal transition_895_preds : BooleanArray(0 downto 0);
  signal transition_896_symbol_out : boolean;
  signal transition_896_preds : BooleanArray(1 downto 0);
  signal transition_898_symbol_out : boolean;
  signal transition_898_preds : BooleanArray(0 downto 0);
  signal transition_899_symbol_out : boolean;
  signal transition_899_preds : BooleanArray(0 downto 0);
  signal transition_900_symbol_out : boolean;
  signal transition_900_preds : BooleanArray(0 downto 0);
  signal transition_901_symbol_out : boolean;
  signal transition_901_preds : BooleanArray(0 downto 0);
  signal transition_902_symbol_out : boolean;
  signal transition_902_preds : BooleanArray(0 downto 0);
  signal transition_903_symbol_out : boolean;
  signal transition_903_preds : BooleanArray(0 downto 0);
  signal transition_907_symbol_out : boolean;
  signal transition_907_preds : BooleanArray(0 downto 0);
  signal transition_908_symbol_out : boolean;
  signal transition_908_preds : BooleanArray(0 downto 0);
  signal transition_909_symbol_out : boolean;
  signal transition_909_preds : BooleanArray(0 downto 0);
  signal transition_910_symbol_out : boolean;
  signal transition_910_preds : BooleanArray(0 downto 0);
  signal transition_914_symbol_out : boolean;
  signal transition_914_preds : BooleanArray(0 downto 0);
  signal transition_915_symbol_out : boolean;
  signal transition_915_preds : BooleanArray(0 downto 0);
  signal transition_916_symbol_out : boolean;
  signal transition_916_preds : BooleanArray(0 downto 0);
  signal transition_917_symbol_out : boolean;
  signal transition_917_preds : BooleanArray(0 downto 0);
  signal transition_921_symbol_out : boolean;
  signal transition_921_preds : BooleanArray(1 downto 0);
  signal transition_922_symbol_out : boolean;
  signal transition_922_preds : BooleanArray(0 downto 0);
  signal transition_923_symbol_out : boolean;
  signal transition_923_preds : BooleanArray(0 downto 0);
  signal transition_924_symbol_out : boolean;
  signal transition_924_preds : BooleanArray(0 downto 0);
  signal transition_925_symbol_out : boolean;
  signal transition_925_preds : BooleanArray(0 downto 0);
  signal transition_929_symbol_out : boolean;
  signal transition_929_preds : BooleanArray(0 downto 0);
  signal transition_930_symbol_out : boolean;
  signal transition_930_preds : BooleanArray(0 downto 0);
  signal transition_931_symbol_out : boolean;
  signal transition_931_preds : BooleanArray(0 downto 0);
  signal transition_932_symbol_out : boolean;
  signal transition_932_preds : BooleanArray(0 downto 0);
  signal transition_936_symbol_out : boolean;
  signal transition_936_preds : BooleanArray(1 downto 0);
  signal transition_937_symbol_out : boolean;
  signal transition_937_preds : BooleanArray(0 downto 0);
  signal transition_938_symbol_out : boolean;
  signal transition_938_preds : BooleanArray(0 downto 0);
  signal transition_939_symbol_out : boolean;
  signal transition_939_preds : BooleanArray(0 downto 0);
  signal transition_940_symbol_out : boolean;
  signal transition_940_preds : BooleanArray(0 downto 0);
  signal transition_945_symbol_out : boolean;
  signal transition_945_preds : BooleanArray(0 downto 0);
  signal transition_946_symbol_out : boolean;
  signal transition_946_preds : BooleanArray(0 downto 0);
  signal transition_947_symbol_out : boolean;
  signal transition_947_preds : BooleanArray(1 downto 0);
  signal transition_949_symbol_out : boolean;
  signal transition_949_preds : BooleanArray(0 downto 0);
  signal transition_950_symbol_out : boolean;
  signal transition_950_preds : BooleanArray(0 downto 0);
  signal transition_951_symbol_out : boolean;
  signal transition_951_preds : BooleanArray(0 downto 0);
  signal transition_952_symbol_out : boolean;
  signal transition_952_preds : BooleanArray(0 downto 0);
  signal transition_953_symbol_out : boolean;
  signal transition_953_preds : BooleanArray(0 downto 0);
  signal transition_954_symbol_out : boolean;
  signal transition_954_preds : BooleanArray(0 downto 0);
  signal transition_958_symbol_out : boolean;
  signal transition_958_preds : BooleanArray(1 downto 0);
  signal transition_959_symbol_out : boolean;
  signal transition_959_preds : BooleanArray(0 downto 0);
  signal transition_960_symbol_out : boolean;
  signal transition_960_preds : BooleanArray(0 downto 0);
  signal transition_961_symbol_out : boolean;
  signal transition_961_preds : BooleanArray(0 downto 0);
  signal transition_962_symbol_out : boolean;
  signal transition_962_preds : BooleanArray(0 downto 0);
  signal transition_966_symbol_out : boolean;
  signal transition_966_preds : BooleanArray(0 downto 0);
  signal transition_967_symbol_out : boolean;
  signal transition_967_preds : BooleanArray(0 downto 0);
  signal transition_968_symbol_out : boolean;
  signal transition_968_preds : BooleanArray(0 downto 0);
  signal transition_969_symbol_out : boolean;
  signal transition_969_preds : BooleanArray(0 downto 0);
  signal transition_973_symbol_out : boolean;
  signal transition_973_preds : BooleanArray(0 downto 0);
  signal transition_974_symbol_out : boolean;
  signal transition_974_preds : BooleanArray(0 downto 0);
  signal transition_975_symbol_out : boolean;
  signal transition_975_preds : BooleanArray(0 downto 0);
  signal transition_976_symbol_out : boolean;
  signal transition_976_preds : BooleanArray(0 downto 0);
  signal transition_980_symbol_out : boolean;
  signal transition_980_preds : BooleanArray(0 downto 0);
  signal transition_981_symbol_out : boolean;
  signal transition_981_preds : BooleanArray(0 downto 0);
  signal transition_982_symbol_out : boolean;
  signal transition_982_preds : BooleanArray(0 downto 0);
  signal transition_983_symbol_out : boolean;
  signal transition_983_preds : BooleanArray(0 downto 0);
  signal transition_987_symbol_out : boolean;
  signal transition_987_preds : BooleanArray(1 downto 0);
  signal transition_988_symbol_out : boolean;
  signal transition_988_preds : BooleanArray(0 downto 0);
  signal transition_989_symbol_out : boolean;
  signal transition_989_preds : BooleanArray(0 downto 0);
  signal transition_990_symbol_out : boolean;
  signal transition_990_preds : BooleanArray(0 downto 0);
  signal transition_991_symbol_out : boolean;
  signal transition_991_preds : BooleanArray(0 downto 0);
  signal transition_995_symbol_out : boolean;
  signal transition_995_preds : BooleanArray(0 downto 0);
  signal transition_996_symbol_out : boolean;
  signal transition_996_preds : BooleanArray(0 downto 0);
  signal transition_997_symbol_out : boolean;
  signal transition_997_preds : BooleanArray(0 downto 0);
  signal transition_998_symbol_out : boolean;
  signal transition_998_preds : BooleanArray(0 downto 0);
  signal transition_1002_symbol_out : boolean;
  signal transition_1002_preds : BooleanArray(1 downto 0);
  signal transition_1003_symbol_out : boolean;
  signal transition_1003_preds : BooleanArray(0 downto 0);
  signal transition_1004_symbol_out : boolean;
  signal transition_1004_preds : BooleanArray(0 downto 0);
  signal transition_1005_symbol_out : boolean;
  signal transition_1005_preds : BooleanArray(0 downto 0);
  signal transition_1006_symbol_out : boolean;
  signal transition_1006_preds : BooleanArray(0 downto 0);
  signal transition_1011_symbol_out : boolean;
  signal transition_1011_preds : BooleanArray(0 downto 0);
  signal transition_1012_symbol_out : boolean;
  signal transition_1012_preds : BooleanArray(0 downto 0);
  signal transition_1013_symbol_out : boolean;
  signal transition_1013_preds : BooleanArray(1 downto 0);
  signal transition_1014_symbol_out : boolean;
  signal transition_1014_preds : BooleanArray(0 downto 0);
  signal transition_1015_symbol_out : boolean;
  signal transition_1015_preds : BooleanArray(0 downto 0);
  signal transition_1016_symbol_out : boolean;
  signal transition_1016_preds : BooleanArray(0 downto 0);
  signal transition_1017_symbol_out : boolean;
  signal transition_1017_preds : BooleanArray(0 downto 0);
  signal transition_1018_symbol_out : boolean;
  signal transition_1018_preds : BooleanArray(0 downto 0);
  signal transition_1022_symbol_out : boolean;
  signal transition_1022_preds : BooleanArray(0 downto 0);
  signal transition_1023_symbol_out : boolean;
  signal transition_1023_preds : BooleanArray(0 downto 0);
  signal transition_1024_symbol_out : boolean;
  signal transition_1024_preds : BooleanArray(0 downto 0);
  signal transition_1025_symbol_out : boolean;
  signal transition_1025_preds : BooleanArray(0 downto 0);
  signal transition_1029_symbol_out : boolean;
  signal transition_1029_preds : BooleanArray(0 downto 0);
  signal transition_1030_symbol_out : boolean;
  signal transition_1030_preds : BooleanArray(0 downto 0);
  signal transition_1031_symbol_out : boolean;
  signal transition_1031_preds : BooleanArray(0 downto 0);
  signal transition_1032_symbol_out : boolean;
  signal transition_1032_preds : BooleanArray(0 downto 0);
  signal transition_1036_symbol_out : boolean;
  signal transition_1036_preds : BooleanArray(1 downto 0);
  signal transition_1037_symbol_out : boolean;
  signal transition_1037_preds : BooleanArray(0 downto 0);
  signal transition_1038_symbol_out : boolean;
  signal transition_1038_preds : BooleanArray(0 downto 0);
  signal transition_1039_symbol_out : boolean;
  signal transition_1039_preds : BooleanArray(0 downto 0);
  signal transition_1040_symbol_out : boolean;
  signal transition_1040_preds : BooleanArray(0 downto 0);
  signal transition_1044_symbol_out : boolean;
  signal transition_1044_preds : BooleanArray(0 downto 0);
  signal transition_1045_symbol_out : boolean;
  signal transition_1045_preds : BooleanArray(0 downto 0);
  signal transition_1046_symbol_out : boolean;
  signal transition_1046_preds : BooleanArray(0 downto 0);
  signal transition_1047_symbol_out : boolean;
  signal transition_1047_preds : BooleanArray(0 downto 0);
  signal transition_1051_symbol_out : boolean;
  signal transition_1051_preds : BooleanArray(1 downto 0);
  signal transition_1052_symbol_out : boolean;
  signal transition_1052_preds : BooleanArray(0 downto 0);
  signal transition_1053_symbol_out : boolean;
  signal transition_1053_preds : BooleanArray(0 downto 0);
  signal transition_1054_symbol_out : boolean;
  signal transition_1054_preds : BooleanArray(0 downto 0);
  signal transition_1055_symbol_out : boolean;
  signal transition_1055_preds : BooleanArray(0 downto 0);
  signal transition_1060_symbol_out : boolean;
  signal transition_1060_preds : BooleanArray(0 downto 0);
  signal transition_1061_symbol_out : boolean;
  signal transition_1061_preds : BooleanArray(0 downto 0);
  signal transition_1062_symbol_out : boolean;
  signal transition_1062_preds : BooleanArray(1 downto 0);
  signal transition_1064_symbol_out : boolean;
  signal transition_1064_preds : BooleanArray(0 downto 0);
  signal transition_1065_symbol_out : boolean;
  signal transition_1065_preds : BooleanArray(0 downto 0);
  signal transition_1066_symbol_out : boolean;
  signal transition_1066_preds : BooleanArray(0 downto 0);
  signal transition_1067_symbol_out : boolean;
  signal transition_1067_preds : BooleanArray(0 downto 0);
  signal transition_1068_symbol_out : boolean;
  signal transition_1068_preds : BooleanArray(0 downto 0);
  signal transition_1069_symbol_out : boolean;
  signal transition_1069_preds : BooleanArray(0 downto 0);
  signal transition_1073_symbol_out : boolean;
  signal transition_1073_preds : BooleanArray(0 downto 0);
  signal transition_1074_symbol_out : boolean;
  signal transition_1074_preds : BooleanArray(0 downto 0);
  signal transition_1075_symbol_out : boolean;
  signal transition_1075_preds : BooleanArray(0 downto 0);
  signal transition_1076_symbol_out : boolean;
  signal transition_1076_preds : BooleanArray(0 downto 0);
  signal transition_1080_symbol_out : boolean;
  signal transition_1080_preds : BooleanArray(0 downto 0);
  signal transition_1081_symbol_out : boolean;
  signal transition_1081_preds : BooleanArray(0 downto 0);
  signal transition_1082_symbol_out : boolean;
  signal transition_1082_preds : BooleanArray(0 downto 0);
  signal transition_1083_symbol_out : boolean;
  signal transition_1083_preds : BooleanArray(0 downto 0);
  signal transition_1087_symbol_out : boolean;
  signal transition_1087_preds : BooleanArray(1 downto 0);
  signal transition_1088_symbol_out : boolean;
  signal transition_1088_preds : BooleanArray(0 downto 0);
  signal transition_1089_symbol_out : boolean;
  signal transition_1089_preds : BooleanArray(0 downto 0);
  signal transition_1090_symbol_out : boolean;
  signal transition_1090_preds : BooleanArray(0 downto 0);
  signal transition_1091_symbol_out : boolean;
  signal transition_1091_preds : BooleanArray(0 downto 0);
  signal transition_1095_symbol_out : boolean;
  signal transition_1095_preds : BooleanArray(0 downto 0);
  signal transition_1096_symbol_out : boolean;
  signal transition_1096_preds : BooleanArray(0 downto 0);
  signal transition_1097_symbol_out : boolean;
  signal transition_1097_preds : BooleanArray(0 downto 0);
  signal transition_1098_symbol_out : boolean;
  signal transition_1098_preds : BooleanArray(0 downto 0);
  signal transition_1102_symbol_out : boolean;
  signal transition_1102_preds : BooleanArray(1 downto 0);
  signal transition_1103_symbol_out : boolean;
  signal transition_1103_preds : BooleanArray(0 downto 0);
  signal transition_1104_symbol_out : boolean;
  signal transition_1104_preds : BooleanArray(0 downto 0);
  signal transition_1105_symbol_out : boolean;
  signal transition_1105_preds : BooleanArray(0 downto 0);
  signal transition_1106_symbol_out : boolean;
  signal transition_1106_preds : BooleanArray(0 downto 0);
  signal transition_1111_symbol_out : boolean;
  signal transition_1111_preds : BooleanArray(0 downto 0);
  signal transition_1112_symbol_out : boolean;
  signal transition_1112_preds : BooleanArray(0 downto 0);
  signal transition_1113_symbol_out : boolean;
  signal transition_1113_preds : BooleanArray(1 downto 0);
  signal transition_1115_symbol_out : boolean;
  signal transition_1115_preds : BooleanArray(0 downto 0);
  signal transition_1116_symbol_out : boolean;
  signal transition_1116_preds : BooleanArray(0 downto 0);
  signal transition_1117_symbol_out : boolean;
  signal transition_1117_preds : BooleanArray(0 downto 0);
  signal transition_1118_symbol_out : boolean;
  signal transition_1118_preds : BooleanArray(0 downto 0);
  signal transition_1119_symbol_out : boolean;
  signal transition_1119_preds : BooleanArray(0 downto 0);
  signal transition_1120_symbol_out : boolean;
  signal transition_1120_preds : BooleanArray(0 downto 0);
  signal transition_1124_symbol_out : boolean;
  signal transition_1124_preds : BooleanArray(1 downto 0);
  signal transition_1125_symbol_out : boolean;
  signal transition_1125_preds : BooleanArray(0 downto 0);
  signal transition_1126_symbol_out : boolean;
  signal transition_1126_preds : BooleanArray(0 downto 0);
  signal transition_1127_symbol_out : boolean;
  signal transition_1127_preds : BooleanArray(0 downto 0);
  signal transition_1128_symbol_out : boolean;
  signal transition_1128_preds : BooleanArray(0 downto 0);
  signal transition_1132_symbol_out : boolean;
  signal transition_1132_preds : BooleanArray(0 downto 0);
  signal transition_1133_symbol_out : boolean;
  signal transition_1133_preds : BooleanArray(0 downto 0);
  signal transition_1134_symbol_out : boolean;
  signal transition_1134_preds : BooleanArray(0 downto 0);
  signal transition_1135_symbol_out : boolean;
  signal transition_1135_preds : BooleanArray(0 downto 0);
  signal transition_1139_symbol_out : boolean;
  signal transition_1139_preds : BooleanArray(0 downto 0);
  signal transition_1140_symbol_out : boolean;
  signal transition_1140_preds : BooleanArray(0 downto 0);
  signal transition_1141_symbol_out : boolean;
  signal transition_1141_preds : BooleanArray(0 downto 0);
  signal transition_1142_symbol_out : boolean;
  signal transition_1142_preds : BooleanArray(0 downto 0);
  signal transition_1146_symbol_out : boolean;
  signal transition_1146_preds : BooleanArray(0 downto 0);
  signal transition_1147_symbol_out : boolean;
  signal transition_1147_preds : BooleanArray(0 downto 0);
  signal transition_1148_symbol_out : boolean;
  signal transition_1148_preds : BooleanArray(0 downto 0);
  signal transition_1149_symbol_out : boolean;
  signal transition_1149_preds : BooleanArray(0 downto 0);
  signal transition_1153_symbol_out : boolean;
  signal transition_1153_preds : BooleanArray(1 downto 0);
  signal transition_1154_symbol_out : boolean;
  signal transition_1154_preds : BooleanArray(0 downto 0);
  signal transition_1155_symbol_out : boolean;
  signal transition_1155_preds : BooleanArray(0 downto 0);
  signal transition_1156_symbol_out : boolean;
  signal transition_1156_preds : BooleanArray(0 downto 0);
  signal transition_1157_symbol_out : boolean;
  signal transition_1157_preds : BooleanArray(0 downto 0);
  signal transition_1161_symbol_out : boolean;
  signal transition_1161_preds : BooleanArray(0 downto 0);
  signal transition_1162_symbol_out : boolean;
  signal transition_1162_preds : BooleanArray(0 downto 0);
  signal transition_1163_symbol_out : boolean;
  signal transition_1163_preds : BooleanArray(0 downto 0);
  signal transition_1164_symbol_out : boolean;
  signal transition_1164_preds : BooleanArray(0 downto 0);
  signal transition_1168_symbol_out : boolean;
  signal transition_1168_preds : BooleanArray(1 downto 0);
  signal transition_1169_symbol_out : boolean;
  signal transition_1169_preds : BooleanArray(0 downto 0);
  signal transition_1170_symbol_out : boolean;
  signal transition_1170_preds : BooleanArray(0 downto 0);
  signal transition_1171_symbol_out : boolean;
  signal transition_1171_preds : BooleanArray(0 downto 0);
  signal transition_1172_symbol_out : boolean;
  signal transition_1172_preds : BooleanArray(0 downto 0);
  signal transition_1177_symbol_out : boolean;
  signal transition_1177_preds : BooleanArray(0 downto 0);
  signal transition_1178_symbol_out : boolean;
  signal transition_1178_preds : BooleanArray(0 downto 0);
  signal transition_1179_symbol_out : boolean;
  signal transition_1179_preds : BooleanArray(1 downto 0);
  signal transition_1180_symbol_out : boolean;
  signal transition_1180_preds : BooleanArray(0 downto 0);
  signal transition_1181_symbol_out : boolean;
  signal transition_1181_preds : BooleanArray(0 downto 0);
  signal transition_1182_symbol_out : boolean;
  signal transition_1182_preds : BooleanArray(0 downto 0);
  signal transition_1183_symbol_out : boolean;
  signal transition_1183_preds : BooleanArray(0 downto 0);
  signal transition_1187_symbol_out : boolean;
  signal transition_1187_preds : BooleanArray(1 downto 0);
  signal transition_1188_symbol_out : boolean;
  signal transition_1188_preds : BooleanArray(0 downto 0);
  signal transition_1189_symbol_out : boolean;
  signal transition_1189_preds : BooleanArray(0 downto 0);
  signal transition_1190_symbol_out : boolean;
  signal transition_1190_preds : BooleanArray(0 downto 0);
  signal transition_1191_symbol_out : boolean;
  signal transition_1191_preds : BooleanArray(0 downto 0);
  signal transition_1195_symbol_out : boolean;
  signal transition_1195_preds : BooleanArray(1 downto 0);
  signal transition_1196_symbol_out : boolean;
  signal transition_1196_preds : BooleanArray(0 downto 0);
  signal transition_1197_symbol_out : boolean;
  signal transition_1197_preds : BooleanArray(0 downto 0);
  signal transition_1198_symbol_out : boolean;
  signal transition_1198_preds : BooleanArray(0 downto 0);
  signal transition_1199_symbol_out : boolean;
  signal transition_1199_preds : BooleanArray(0 downto 0);
  signal transition_1204_symbol_out : boolean;
  signal transition_1204_preds : BooleanArray(0 downto 0);
  signal transition_1205_symbol_out : boolean;
  signal transition_1205_preds : BooleanArray(0 downto 0);

begin
  place_0_preds(0) <= transition_2_symbol_out;
  place_0_succs(0) <= transition_1_symbol_out;
  place_0 : place
    generic map(marking => true)
    port map(
      preds => place_0_preds,
      succs => place_0_succs,
      token => place_0_token,
      clk   => clk,
      reset => reset);

  place_5_preds(0) <= transition_7_symbol_out;
  place_5_succs(0) <= transition_6_symbol_out;
  place_5 : place
    generic map(marking => false)
    port map(
      preds => place_5_preds,
      succs => place_5_succs,
      token => place_5_token,
      clk   => clk,
      reset => reset);

  place_12_preds(0) <= transition_8_symbol_out;
  place_12_succs(0) <= transition_9_symbol_out;
  place_12 : place
    generic map(marking => false)
    port map(
      preds => place_12_preds,
      succs => place_12_succs,
      token => place_12_token,
      clk   => clk,
      reset => reset);

  place_13_preds(0) <= transition_9_symbol_out;
  place_13_succs(0) <= transition_10_symbol_out;
  place_13 : place
    generic map(marking => false)
    port map(
      preds => place_13_preds,
      succs => place_13_succs,
      token => place_13_token,
      clk   => clk,
      reset => reset);

  place_14_preds(0) <= transition_10_symbol_out;
  place_14_succs(0) <= transition_11_symbol_out;
  place_14 : place
    generic map(marking => false)
    port map(
      preds => place_14_preds,
      succs => place_14_succs,
      token => place_14_token,
      clk   => clk,
      reset => reset);

  place_19_preds(0) <= transition_15_symbol_out;
  place_19_succs(0) <= transition_16_symbol_out;
  place_19 : place
    generic map(marking => false)
    port map(
      preds => place_19_preds,
      succs => place_19_succs,
      token => place_19_token,
      clk   => clk,
      reset => reset);

  place_20_preds(0) <= transition_16_symbol_out;
  place_20_succs(0) <= transition_17_symbol_out;
  place_20 : place
    generic map(marking => false)
    port map(
      preds => place_20_preds,
      succs => place_20_succs,
      token => place_20_token,
      clk   => clk,
      reset => reset);

  place_21_preds(0) <= transition_17_symbol_out;
  place_21_succs(0) <= transition_18_symbol_out;
  place_21 : place
    generic map(marking => false)
    port map(
      preds => place_21_preds,
      succs => place_21_succs,
      token => place_21_token,
      clk   => clk,
      reset => reset);

  place_26_preds(0) <= transition_22_symbol_out;
  place_26_succs(0) <= transition_23_symbol_out;
  place_26 : place
    generic map(marking => false)
    port map(
      preds => place_26_preds,
      succs => place_26_succs,
      token => place_26_token,
      clk   => clk,
      reset => reset);

  place_27_preds(0) <= transition_23_symbol_out;
  place_27_succs(0) <= transition_24_symbol_out;
  place_27 : place
    generic map(marking => false)
    port map(
      preds => place_27_preds,
      succs => place_27_succs,
      token => place_27_token,
      clk   => clk,
      reset => reset);

  place_28_preds(0) <= transition_24_symbol_out;
  place_28_succs(0) <= transition_25_symbol_out;
  place_28 : place
    generic map(marking => false)
    port map(
      preds => place_28_preds,
      succs => place_28_succs,
      token => place_28_token,
      clk   => clk,
      reset => reset);

  place_34_preds(0) <= transition_30_symbol_out;
  place_34_succs(0) <= transition_31_symbol_out;
  place_34 : place
    generic map(marking => false)
    port map(
      preds => place_34_preds,
      succs => place_34_succs,
      token => place_34_token,
      clk   => clk,
      reset => reset);

  place_35_preds(0) <= transition_31_symbol_out;
  place_35_succs(0) <= transition_32_symbol_out;
  place_35 : place
    generic map(marking => false)
    port map(
      preds => place_35_preds,
      succs => place_35_succs,
      token => place_35_token,
      clk   => clk,
      reset => reset);

  place_36_preds(0) <= transition_32_symbol_out;
  place_36_succs(0) <= transition_33_symbol_out;
  place_36 : place
    generic map(marking => false)
    port map(
      preds => place_36_preds,
      succs => place_36_succs,
      token => place_36_token,
      clk   => clk,
      reset => reset);

  place_41_preds(0) <= transition_37_symbol_out;
  place_41_succs(0) <= transition_38_symbol_out;
  place_41 : place
    generic map(marking => false)
    port map(
      preds => place_41_preds,
      succs => place_41_succs,
      token => place_41_token,
      clk   => clk,
      reset => reset);

  place_42_preds(0) <= transition_38_symbol_out;
  place_42_succs(0) <= transition_39_symbol_out;
  place_42 : place
    generic map(marking => false)
    port map(
      preds => place_42_preds,
      succs => place_42_succs,
      token => place_42_token,
      clk   => clk,
      reset => reset);

  place_43_preds(0) <= transition_39_symbol_out;
  place_43_succs(0) <= transition_40_symbol_out;
  place_43 : place
    generic map(marking => false)
    port map(
      preds => place_43_preds,
      succs => place_43_succs,
      token => place_43_token,
      clk   => clk,
      reset => reset);

  place_49_preds(0) <= transition_45_symbol_out;
  place_49_succs(0) <= transition_46_symbol_out;
  place_49 : place
    generic map(marking => false)
    port map(
      preds => place_49_preds,
      succs => place_49_succs,
      token => place_49_token,
      clk   => clk,
      reset => reset);

  place_50_preds(0) <= transition_46_symbol_out;
  place_50_succs(0) <= transition_47_symbol_out;
  place_50 : place
    generic map(marking => false)
    port map(
      preds => place_50_preds,
      succs => place_50_succs,
      token => place_50_token,
      clk   => clk,
      reset => reset);

  place_51_preds(0) <= transition_47_symbol_out;
  place_51_succs(0) <= transition_48_symbol_out;
  place_51 : place
    generic map(marking => false)
    port map(
      preds => place_51_preds,
      succs => place_51_succs,
      token => place_51_token,
      clk   => clk,
      reset => reset);

  place_52_preds(0) <= transition_54_symbol_out;
  place_52_succs(0) <= transition_53_symbol_out;
  place_52 : place
    generic map(marking => false)
    port map(
      preds => place_52_preds,
      succs => place_52_succs,
      token => place_52_token,
      clk   => clk,
      reset => reset);

  place_56_preds(0) <= transition_58_symbol_out;
  place_56_succs(0) <= transition_57_symbol_out;
  place_56 : place
    generic map(marking => false)
    port map(
      preds => place_56_preds,
      succs => place_56_succs,
      token => place_56_token,
      clk   => clk,
      reset => reset);

  place_64_preds(0) <= transition_60_symbol_out;
  place_64_succs(0) <= transition_61_symbol_out;
  place_64 : place
    generic map(marking => false)
    port map(
      preds => place_64_preds,
      succs => place_64_succs,
      token => place_64_token,
      clk   => clk,
      reset => reset);

  place_65_preds(0) <= transition_61_symbol_out;
  place_65_succs(0) <= transition_62_symbol_out;
  place_65 : place
    generic map(marking => false)
    port map(
      preds => place_65_preds,
      succs => place_65_succs,
      token => place_65_token,
      clk   => clk,
      reset => reset);

  place_66_preds(0) <= transition_62_symbol_out;
  place_66_succs(0) <= transition_63_symbol_out;
  place_66 : place
    generic map(marking => false)
    port map(
      preds => place_66_preds,
      succs => place_66_succs,
      token => place_66_token,
      clk   => clk,
      reset => reset);

  place_71_preds(0) <= transition_67_symbol_out;
  place_71_succs(0) <= transition_68_symbol_out;
  place_71 : place
    generic map(marking => false)
    port map(
      preds => place_71_preds,
      succs => place_71_succs,
      token => place_71_token,
      clk   => clk,
      reset => reset);

  place_72_preds(0) <= transition_68_symbol_out;
  place_72_succs(0) <= transition_69_symbol_out;
  place_72 : place
    generic map(marking => false)
    port map(
      preds => place_72_preds,
      succs => place_72_succs,
      token => place_72_token,
      clk   => clk,
      reset => reset);

  place_73_preds(0) <= transition_69_symbol_out;
  place_73_succs(0) <= transition_70_symbol_out;
  place_73 : place
    generic map(marking => false)
    port map(
      preds => place_73_preds,
      succs => place_73_succs,
      token => place_73_token,
      clk   => clk,
      reset => reset);

  place_78_preds(0) <= transition_74_symbol_out;
  place_78_succs(0) <= transition_75_symbol_out;
  place_78 : place
    generic map(marking => false)
    port map(
      preds => place_78_preds,
      succs => place_78_succs,
      token => place_78_token,
      clk   => clk,
      reset => reset);

  place_79_preds(0) <= transition_75_symbol_out;
  place_79_succs(0) <= transition_76_symbol_out;
  place_79 : place
    generic map(marking => false)
    port map(
      preds => place_79_preds,
      succs => place_79_succs,
      token => place_79_token,
      clk   => clk,
      reset => reset);

  place_80_preds(0) <= transition_76_symbol_out;
  place_80_succs(0) <= transition_77_symbol_out;
  place_80 : place
    generic map(marking => false)
    port map(
      preds => place_80_preds,
      succs => place_80_succs,
      token => place_80_token,
      clk   => clk,
      reset => reset);

  place_86_preds(0) <= transition_82_symbol_out;
  place_86_succs(0) <= transition_83_symbol_out;
  place_86 : place
    generic map(marking => false)
    port map(
      preds => place_86_preds,
      succs => place_86_succs,
      token => place_86_token,
      clk   => clk,
      reset => reset);

  place_87_preds(0) <= transition_83_symbol_out;
  place_87_succs(0) <= transition_84_symbol_out;
  place_87 : place
    generic map(marking => false)
    port map(
      preds => place_87_preds,
      succs => place_87_succs,
      token => place_87_token,
      clk   => clk,
      reset => reset);

  place_88_preds(0) <= transition_84_symbol_out;
  place_88_succs(0) <= transition_85_symbol_out;
  place_88 : place
    generic map(marking => false)
    port map(
      preds => place_88_preds,
      succs => place_88_succs,
      token => place_88_token,
      clk   => clk,
      reset => reset);

  place_93_preds(0) <= transition_89_symbol_out;
  place_93_succs(0) <= transition_90_symbol_out;
  place_93 : place
    generic map(marking => false)
    port map(
      preds => place_93_preds,
      succs => place_93_succs,
      token => place_93_token,
      clk   => clk,
      reset => reset);

  place_94_preds(0) <= transition_90_symbol_out;
  place_94_succs(0) <= transition_91_symbol_out;
  place_94 : place
    generic map(marking => false)
    port map(
      preds => place_94_preds,
      succs => place_94_succs,
      token => place_94_token,
      clk   => clk,
      reset => reset);

  place_95_preds(0) <= transition_91_symbol_out;
  place_95_succs(0) <= transition_92_symbol_out;
  place_95 : place
    generic map(marking => false)
    port map(
      preds => place_95_preds,
      succs => place_95_succs,
      token => place_95_token,
      clk   => clk,
      reset => reset);

  place_101_preds(0) <= transition_97_symbol_out;
  place_101_succs(0) <= transition_98_symbol_out;
  place_101 : place
    generic map(marking => false)
    port map(
      preds => place_101_preds,
      succs => place_101_succs,
      token => place_101_token,
      clk   => clk,
      reset => reset);

  place_102_preds(0) <= transition_98_symbol_out;
  place_102_succs(0) <= transition_99_symbol_out;
  place_102 : place
    generic map(marking => false)
    port map(
      preds => place_102_preds,
      succs => place_102_succs,
      token => place_102_token,
      clk   => clk,
      reset => reset);

  place_103_preds(0) <= transition_99_symbol_out;
  place_103_succs(0) <= transition_100_symbol_out;
  place_103 : place
    generic map(marking => false)
    port map(
      preds => place_103_preds,
      succs => place_103_succs,
      token => place_103_token,
      clk   => clk,
      reset => reset);

  place_104_preds(0) <= transition_106_symbol_out;
  place_104_succs(0) <= transition_105_symbol_out;
  place_104 : place
    generic map(marking => false)
    port map(
      preds => place_104_preds,
      succs => place_104_succs,
      token => place_104_token,
      clk   => clk,
      reset => reset);

  place_108_preds(0) <= transition_110_symbol_out;
  place_108_succs(0) <= transition_109_symbol_out;
  place_108 : place
    generic map(marking => false)
    port map(
      preds => place_108_preds,
      succs => place_108_succs,
      token => place_108_token,
      clk   => clk,
      reset => reset);

  place_116_preds(0) <= transition_112_symbol_out;
  place_116_succs(0) <= transition_113_symbol_out;
  place_116 : place
    generic map(marking => false)
    port map(
      preds => place_116_preds,
      succs => place_116_succs,
      token => place_116_token,
      clk   => clk,
      reset => reset);

  place_117_preds(0) <= transition_113_symbol_out;
  place_117_succs(0) <= transition_114_symbol_out;
  place_117 : place
    generic map(marking => false)
    port map(
      preds => place_117_preds,
      succs => place_117_succs,
      token => place_117_token,
      clk   => clk,
      reset => reset);

  place_118_preds(0) <= transition_114_symbol_out;
  place_118_succs(0) <= transition_115_symbol_out;
  place_118 : place
    generic map(marking => false)
    port map(
      preds => place_118_preds,
      succs => place_118_succs,
      token => place_118_token,
      clk   => clk,
      reset => reset);

  place_125_preds(0) <= transition_121_symbol_out;
  place_125_succs(0) <= transition_122_symbol_out;
  place_125 : place
    generic map(marking => false)
    port map(
      preds => place_125_preds,
      succs => place_125_succs,
      token => place_125_token,
      clk   => clk,
      reset => reset);

  place_126_preds(0) <= transition_122_symbol_out;
  place_126_succs(0) <= transition_123_symbol_out;
  place_126 : place
    generic map(marking => false)
    port map(
      preds => place_126_preds,
      succs => place_126_succs,
      token => place_126_token,
      clk   => clk,
      reset => reset);

  place_127_preds(0) <= transition_123_symbol_out;
  place_127_succs(0) <= transition_124_symbol_out;
  place_127 : place
    generic map(marking => false)
    port map(
      preds => place_127_preds,
      succs => place_127_succs,
      token => place_127_token,
      clk   => clk,
      reset => reset);

  place_132_preds(0) <= transition_128_symbol_out;
  place_132_succs(0) <= transition_129_symbol_out;
  place_132 : place
    generic map(marking => false)
    port map(
      preds => place_132_preds,
      succs => place_132_succs,
      token => place_132_token,
      clk   => clk,
      reset => reset);

  place_133_preds(0) <= transition_129_symbol_out;
  place_133_succs(0) <= transition_130_symbol_out;
  place_133 : place
    generic map(marking => false)
    port map(
      preds => place_133_preds,
      succs => place_133_succs,
      token => place_133_token,
      clk   => clk,
      reset => reset);

  place_134_preds(0) <= transition_130_symbol_out;
  place_134_succs(0) <= transition_131_symbol_out;
  place_134 : place
    generic map(marking => false)
    port map(
      preds => place_134_preds,
      succs => place_134_succs,
      token => place_134_token,
      clk   => clk,
      reset => reset);

  place_139_preds(0) <= transition_135_symbol_out;
  place_139_succs(0) <= transition_136_symbol_out;
  place_139 : place
    generic map(marking => false)
    port map(
      preds => place_139_preds,
      succs => place_139_succs,
      token => place_139_token,
      clk   => clk,
      reset => reset);

  place_140_preds(0) <= transition_136_symbol_out;
  place_140_succs(0) <= transition_137_symbol_out;
  place_140 : place
    generic map(marking => false)
    port map(
      preds => place_140_preds,
      succs => place_140_succs,
      token => place_140_token,
      clk   => clk,
      reset => reset);

  place_141_preds(0) <= transition_137_symbol_out;
  place_141_succs(0) <= transition_138_symbol_out;
  place_141 : place
    generic map(marking => false)
    port map(
      preds => place_141_preds,
      succs => place_141_succs,
      token => place_141_token,
      clk   => clk,
      reset => reset);

  place_147_preds(0) <= transition_143_symbol_out;
  place_147_succs(0) <= transition_144_symbol_out;
  place_147 : place
    generic map(marking => false)
    port map(
      preds => place_147_preds,
      succs => place_147_succs,
      token => place_147_token,
      clk   => clk,
      reset => reset);

  place_148_preds(0) <= transition_144_symbol_out;
  place_148_succs(0) <= transition_145_symbol_out;
  place_148 : place
    generic map(marking => false)
    port map(
      preds => place_148_preds,
      succs => place_148_succs,
      token => place_148_token,
      clk   => clk,
      reset => reset);

  place_149_preds(0) <= transition_145_symbol_out;
  place_149_succs(0) <= transition_146_symbol_out;
  place_149 : place
    generic map(marking => false)
    port map(
      preds => place_149_preds,
      succs => place_149_succs,
      token => place_149_token,
      clk   => clk,
      reset => reset);

  place_154_preds(0) <= transition_150_symbol_out;
  place_154_succs(0) <= transition_151_symbol_out;
  place_154 : place
    generic map(marking => false)
    port map(
      preds => place_154_preds,
      succs => place_154_succs,
      token => place_154_token,
      clk   => clk,
      reset => reset);

  place_155_preds(0) <= transition_151_symbol_out;
  place_155_succs(0) <= transition_152_symbol_out;
  place_155 : place
    generic map(marking => false)
    port map(
      preds => place_155_preds,
      succs => place_155_succs,
      token => place_155_token,
      clk   => clk,
      reset => reset);

  place_156_preds(0) <= transition_152_symbol_out;
  place_156_succs(0) <= transition_153_symbol_out;
  place_156 : place
    generic map(marking => false)
    port map(
      preds => place_156_preds,
      succs => place_156_succs,
      token => place_156_token,
      clk   => clk,
      reset => reset);

  place_162_preds(0) <= transition_158_symbol_out;
  place_162_succs(0) <= transition_159_symbol_out;
  place_162 : place
    generic map(marking => false)
    port map(
      preds => place_162_preds,
      succs => place_162_succs,
      token => place_162_token,
      clk   => clk,
      reset => reset);

  place_163_preds(0) <= transition_159_symbol_out;
  place_163_succs(0) <= transition_160_symbol_out;
  place_163 : place
    generic map(marking => false)
    port map(
      preds => place_163_preds,
      succs => place_163_succs,
      token => place_163_token,
      clk   => clk,
      reset => reset);

  place_164_preds(0) <= transition_160_symbol_out;
  place_164_succs(0) <= transition_161_symbol_out;
  place_164 : place
    generic map(marking => false)
    port map(
      preds => place_164_preds,
      succs => place_164_succs,
      token => place_164_token,
      clk   => clk,
      reset => reset);

  place_165_preds(0) <= transition_167_symbol_out;
  place_165_succs(0) <= transition_166_symbol_out;
  place_165 : place
    generic map(marking => false)
    port map(
      preds => place_165_preds,
      succs => place_165_succs,
      token => place_165_token,
      clk   => clk,
      reset => reset);

  place_174_preds(0) <= transition_170_symbol_out;
  place_174_succs(0) <= transition_171_symbol_out;
  place_174 : place
    generic map(marking => false)
    port map(
      preds => place_174_preds,
      succs => place_174_succs,
      token => place_174_token,
      clk   => clk,
      reset => reset);

  place_175_preds(0) <= transition_171_symbol_out;
  place_175_succs(0) <= transition_172_symbol_out;
  place_175 : place
    generic map(marking => false)
    port map(
      preds => place_175_preds,
      succs => place_175_succs,
      token => place_175_token,
      clk   => clk,
      reset => reset);

  place_176_preds(0) <= transition_172_symbol_out;
  place_176_succs(0) <= transition_173_symbol_out;
  place_176 : place
    generic map(marking => false)
    port map(
      preds => place_176_preds,
      succs => place_176_succs,
      token => place_176_token,
      clk   => clk,
      reset => reset);

  place_181_preds(0) <= transition_177_symbol_out;
  place_181_succs(0) <= transition_178_symbol_out;
  place_181 : place
    generic map(marking => false)
    port map(
      preds => place_181_preds,
      succs => place_181_succs,
      token => place_181_token,
      clk   => clk,
      reset => reset);

  place_182_preds(0) <= transition_178_symbol_out;
  place_182_succs(0) <= transition_179_symbol_out;
  place_182 : place
    generic map(marking => false)
    port map(
      preds => place_182_preds,
      succs => place_182_succs,
      token => place_182_token,
      clk   => clk,
      reset => reset);

  place_183_preds(0) <= transition_179_symbol_out;
  place_183_succs(0) <= transition_180_symbol_out;
  place_183 : place
    generic map(marking => false)
    port map(
      preds => place_183_preds,
      succs => place_183_succs,
      token => place_183_token,
      clk   => clk,
      reset => reset);

  place_188_preds(0) <= transition_184_symbol_out;
  place_188_succs(0) <= transition_185_symbol_out;
  place_188 : place
    generic map(marking => false)
    port map(
      preds => place_188_preds,
      succs => place_188_succs,
      token => place_188_token,
      clk   => clk,
      reset => reset);

  place_189_preds(0) <= transition_185_symbol_out;
  place_189_succs(0) <= transition_186_symbol_out;
  place_189 : place
    generic map(marking => false)
    port map(
      preds => place_189_preds,
      succs => place_189_succs,
      token => place_189_token,
      clk   => clk,
      reset => reset);

  place_190_preds(0) <= transition_186_symbol_out;
  place_190_succs(0) <= transition_187_symbol_out;
  place_190 : place
    generic map(marking => false)
    port map(
      preds => place_190_preds,
      succs => place_190_succs,
      token => place_190_token,
      clk   => clk,
      reset => reset);

  place_196_preds(0) <= transition_192_symbol_out;
  place_196_succs(0) <= transition_193_symbol_out;
  place_196 : place
    generic map(marking => false)
    port map(
      preds => place_196_preds,
      succs => place_196_succs,
      token => place_196_token,
      clk   => clk,
      reset => reset);

  place_197_preds(0) <= transition_193_symbol_out;
  place_197_succs(0) <= transition_194_symbol_out;
  place_197 : place
    generic map(marking => false)
    port map(
      preds => place_197_preds,
      succs => place_197_succs,
      token => place_197_token,
      clk   => clk,
      reset => reset);

  place_198_preds(0) <= transition_194_symbol_out;
  place_198_succs(0) <= transition_195_symbol_out;
  place_198 : place
    generic map(marking => false)
    port map(
      preds => place_198_preds,
      succs => place_198_succs,
      token => place_198_token,
      clk   => clk,
      reset => reset);

  place_203_preds(0) <= transition_199_symbol_out;
  place_203_succs(0) <= transition_200_symbol_out;
  place_203 : place
    generic map(marking => false)
    port map(
      preds => place_203_preds,
      succs => place_203_succs,
      token => place_203_token,
      clk   => clk,
      reset => reset);

  place_204_preds(0) <= transition_200_symbol_out;
  place_204_succs(0) <= transition_201_symbol_out;
  place_204 : place
    generic map(marking => false)
    port map(
      preds => place_204_preds,
      succs => place_204_succs,
      token => place_204_token,
      clk   => clk,
      reset => reset);

  place_205_preds(0) <= transition_201_symbol_out;
  place_205_succs(0) <= transition_202_symbol_out;
  place_205 : place
    generic map(marking => false)
    port map(
      preds => place_205_preds,
      succs => place_205_succs,
      token => place_205_token,
      clk   => clk,
      reset => reset);

  place_211_preds(0) <= transition_207_symbol_out;
  place_211_succs(0) <= transition_208_symbol_out;
  place_211 : place
    generic map(marking => false)
    port map(
      preds => place_211_preds,
      succs => place_211_succs,
      token => place_211_token,
      clk   => clk,
      reset => reset);

  place_212_preds(0) <= transition_208_symbol_out;
  place_212_succs(0) <= transition_209_symbol_out;
  place_212 : place
    generic map(marking => false)
    port map(
      preds => place_212_preds,
      succs => place_212_succs,
      token => place_212_token,
      clk   => clk,
      reset => reset);

  place_213_preds(0) <= transition_209_symbol_out;
  place_213_succs(0) <= transition_210_symbol_out;
  place_213 : place
    generic map(marking => false)
    port map(
      preds => place_213_preds,
      succs => place_213_succs,
      token => place_213_token,
      clk   => clk,
      reset => reset);

  place_214_preds(0) <= transition_216_symbol_out;
  place_214_succs(0) <= transition_215_symbol_out;
  place_214 : place
    generic map(marking => false)
    port map(
      preds => place_214_preds,
      succs => place_214_succs,
      token => place_214_token,
      clk   => clk,
      reset => reset);

  place_218_preds(0) <= transition_220_symbol_out;
  place_218_succs(0) <= transition_219_symbol_out;
  place_218 : place
    generic map(marking => false)
    port map(
      preds => place_218_preds,
      succs => place_218_succs,
      token => place_218_token,
      clk   => clk,
      reset => reset);

  place_226_preds(0) <= transition_222_symbol_out;
  place_226_succs(0) <= transition_223_symbol_out;
  place_226 : place
    generic map(marking => false)
    port map(
      preds => place_226_preds,
      succs => place_226_succs,
      token => place_226_token,
      clk   => clk,
      reset => reset);

  place_227_preds(0) <= transition_223_symbol_out;
  place_227_succs(0) <= transition_224_symbol_out;
  place_227 : place
    generic map(marking => false)
    port map(
      preds => place_227_preds,
      succs => place_227_succs,
      token => place_227_token,
      clk   => clk,
      reset => reset);

  place_228_preds(0) <= transition_224_symbol_out;
  place_228_succs(0) <= transition_225_symbol_out;
  place_228 : place
    generic map(marking => false)
    port map(
      preds => place_228_preds,
      succs => place_228_succs,
      token => place_228_token,
      clk   => clk,
      reset => reset);

  place_233_preds(0) <= transition_229_symbol_out;
  place_233_succs(0) <= transition_230_symbol_out;
  place_233 : place
    generic map(marking => false)
    port map(
      preds => place_233_preds,
      succs => place_233_succs,
      token => place_233_token,
      clk   => clk,
      reset => reset);

  place_234_preds(0) <= transition_230_symbol_out;
  place_234_succs(0) <= transition_231_symbol_out;
  place_234 : place
    generic map(marking => false)
    port map(
      preds => place_234_preds,
      succs => place_234_succs,
      token => place_234_token,
      clk   => clk,
      reset => reset);

  place_235_preds(0) <= transition_231_symbol_out;
  place_235_succs(0) <= transition_232_symbol_out;
  place_235 : place
    generic map(marking => false)
    port map(
      preds => place_235_preds,
      succs => place_235_succs,
      token => place_235_token,
      clk   => clk,
      reset => reset);

  place_240_preds(0) <= transition_236_symbol_out;
  place_240_succs(0) <= transition_237_symbol_out;
  place_240 : place
    generic map(marking => false)
    port map(
      preds => place_240_preds,
      succs => place_240_succs,
      token => place_240_token,
      clk   => clk,
      reset => reset);

  place_241_preds(0) <= transition_237_symbol_out;
  place_241_succs(0) <= transition_238_symbol_out;
  place_241 : place
    generic map(marking => false)
    port map(
      preds => place_241_preds,
      succs => place_241_succs,
      token => place_241_token,
      clk   => clk,
      reset => reset);

  place_242_preds(0) <= transition_238_symbol_out;
  place_242_succs(0) <= transition_239_symbol_out;
  place_242 : place
    generic map(marking => false)
    port map(
      preds => place_242_preds,
      succs => place_242_succs,
      token => place_242_token,
      clk   => clk,
      reset => reset);

  place_248_preds(0) <= transition_244_symbol_out;
  place_248_succs(0) <= transition_245_symbol_out;
  place_248 : place
    generic map(marking => false)
    port map(
      preds => place_248_preds,
      succs => place_248_succs,
      token => place_248_token,
      clk   => clk,
      reset => reset);

  place_249_preds(0) <= transition_245_symbol_out;
  place_249_succs(0) <= transition_246_symbol_out;
  place_249 : place
    generic map(marking => false)
    port map(
      preds => place_249_preds,
      succs => place_249_succs,
      token => place_249_token,
      clk   => clk,
      reset => reset);

  place_250_preds(0) <= transition_246_symbol_out;
  place_250_succs(0) <= transition_247_symbol_out;
  place_250 : place
    generic map(marking => false)
    port map(
      preds => place_250_preds,
      succs => place_250_succs,
      token => place_250_token,
      clk   => clk,
      reset => reset);

  place_255_preds(0) <= transition_251_symbol_out;
  place_255_succs(0) <= transition_252_symbol_out;
  place_255 : place
    generic map(marking => false)
    port map(
      preds => place_255_preds,
      succs => place_255_succs,
      token => place_255_token,
      clk   => clk,
      reset => reset);

  place_256_preds(0) <= transition_252_symbol_out;
  place_256_succs(0) <= transition_253_symbol_out;
  place_256 : place
    generic map(marking => false)
    port map(
      preds => place_256_preds,
      succs => place_256_succs,
      token => place_256_token,
      clk   => clk,
      reset => reset);

  place_257_preds(0) <= transition_253_symbol_out;
  place_257_succs(0) <= transition_254_symbol_out;
  place_257 : place
    generic map(marking => false)
    port map(
      preds => place_257_preds,
      succs => place_257_succs,
      token => place_257_token,
      clk   => clk,
      reset => reset);

  place_263_preds(0) <= transition_259_symbol_out;
  place_263_succs(0) <= transition_260_symbol_out;
  place_263 : place
    generic map(marking => false)
    port map(
      preds => place_263_preds,
      succs => place_263_succs,
      token => place_263_token,
      clk   => clk,
      reset => reset);

  place_264_preds(0) <= transition_260_symbol_out;
  place_264_succs(0) <= transition_261_symbol_out;
  place_264 : place
    generic map(marking => false)
    port map(
      preds => place_264_preds,
      succs => place_264_succs,
      token => place_264_token,
      clk   => clk,
      reset => reset);

  place_265_preds(0) <= transition_261_symbol_out;
  place_265_succs(0) <= transition_262_symbol_out;
  place_265 : place
    generic map(marking => false)
    port map(
      preds => place_265_preds,
      succs => place_265_succs,
      token => place_265_token,
      clk   => clk,
      reset => reset);

  place_266_preds(0) <= transition_268_symbol_out;
  place_266_succs(0) <= transition_267_symbol_out;
  place_266 : place
    generic map(marking => false)
    port map(
      preds => place_266_preds,
      succs => place_266_succs,
      token => place_266_token,
      clk   => clk,
      reset => reset);

  place_270_preds(0) <= transition_272_symbol_out;
  place_270_succs(0) <= transition_271_symbol_out;
  place_270 : place
    generic map(marking => false)
    port map(
      preds => place_270_preds,
      succs => place_270_succs,
      token => place_270_token,
      clk   => clk,
      reset => reset);

  place_278_preds(0) <= transition_274_symbol_out;
  place_278_succs(0) <= transition_275_symbol_out;
  place_278 : place
    generic map(marking => false)
    port map(
      preds => place_278_preds,
      succs => place_278_succs,
      token => place_278_token,
      clk   => clk,
      reset => reset);

  place_279_preds(0) <= transition_275_symbol_out;
  place_279_succs(0) <= transition_276_symbol_out;
  place_279 : place
    generic map(marking => false)
    port map(
      preds => place_279_preds,
      succs => place_279_succs,
      token => place_279_token,
      clk   => clk,
      reset => reset);

  place_280_preds(0) <= transition_276_symbol_out;
  place_280_succs(0) <= transition_277_symbol_out;
  place_280 : place
    generic map(marking => false)
    port map(
      preds => place_280_preds,
      succs => place_280_succs,
      token => place_280_token,
      clk   => clk,
      reset => reset);

  place_287_preds(0) <= transition_283_symbol_out;
  place_287_succs(0) <= transition_284_symbol_out;
  place_287 : place
    generic map(marking => false)
    port map(
      preds => place_287_preds,
      succs => place_287_succs,
      token => place_287_token,
      clk   => clk,
      reset => reset);

  place_288_preds(0) <= transition_284_symbol_out;
  place_288_succs(0) <= transition_285_symbol_out;
  place_288 : place
    generic map(marking => false)
    port map(
      preds => place_288_preds,
      succs => place_288_succs,
      token => place_288_token,
      clk   => clk,
      reset => reset);

  place_289_preds(0) <= transition_285_symbol_out;
  place_289_succs(0) <= transition_286_symbol_out;
  place_289 : place
    generic map(marking => false)
    port map(
      preds => place_289_preds,
      succs => place_289_succs,
      token => place_289_token,
      clk   => clk,
      reset => reset);

  place_294_preds(0) <= transition_290_symbol_out;
  place_294_succs(0) <= transition_291_symbol_out;
  place_294 : place
    generic map(marking => false)
    port map(
      preds => place_294_preds,
      succs => place_294_succs,
      token => place_294_token,
      clk   => clk,
      reset => reset);

  place_295_preds(0) <= transition_291_symbol_out;
  place_295_succs(0) <= transition_292_symbol_out;
  place_295 : place
    generic map(marking => false)
    port map(
      preds => place_295_preds,
      succs => place_295_succs,
      token => place_295_token,
      clk   => clk,
      reset => reset);

  place_296_preds(0) <= transition_292_symbol_out;
  place_296_succs(0) <= transition_293_symbol_out;
  place_296 : place
    generic map(marking => false)
    port map(
      preds => place_296_preds,
      succs => place_296_succs,
      token => place_296_token,
      clk   => clk,
      reset => reset);

  place_301_preds(0) <= transition_297_symbol_out;
  place_301_succs(0) <= transition_298_symbol_out;
  place_301 : place
    generic map(marking => false)
    port map(
      preds => place_301_preds,
      succs => place_301_succs,
      token => place_301_token,
      clk   => clk,
      reset => reset);

  place_302_preds(0) <= transition_298_symbol_out;
  place_302_succs(0) <= transition_299_symbol_out;
  place_302 : place
    generic map(marking => false)
    port map(
      preds => place_302_preds,
      succs => place_302_succs,
      token => place_302_token,
      clk   => clk,
      reset => reset);

  place_303_preds(0) <= transition_299_symbol_out;
  place_303_succs(0) <= transition_300_symbol_out;
  place_303 : place
    generic map(marking => false)
    port map(
      preds => place_303_preds,
      succs => place_303_succs,
      token => place_303_token,
      clk   => clk,
      reset => reset);

  place_309_preds(0) <= transition_305_symbol_out;
  place_309_succs(0) <= transition_306_symbol_out;
  place_309 : place
    generic map(marking => false)
    port map(
      preds => place_309_preds,
      succs => place_309_succs,
      token => place_309_token,
      clk   => clk,
      reset => reset);

  place_310_preds(0) <= transition_306_symbol_out;
  place_310_succs(0) <= transition_307_symbol_out;
  place_310 : place
    generic map(marking => false)
    port map(
      preds => place_310_preds,
      succs => place_310_succs,
      token => place_310_token,
      clk   => clk,
      reset => reset);

  place_311_preds(0) <= transition_307_symbol_out;
  place_311_succs(0) <= transition_308_symbol_out;
  place_311 : place
    generic map(marking => false)
    port map(
      preds => place_311_preds,
      succs => place_311_succs,
      token => place_311_token,
      clk   => clk,
      reset => reset);

  place_316_preds(0) <= transition_312_symbol_out;
  place_316_succs(0) <= transition_313_symbol_out;
  place_316 : place
    generic map(marking => false)
    port map(
      preds => place_316_preds,
      succs => place_316_succs,
      token => place_316_token,
      clk   => clk,
      reset => reset);

  place_317_preds(0) <= transition_313_symbol_out;
  place_317_succs(0) <= transition_314_symbol_out;
  place_317 : place
    generic map(marking => false)
    port map(
      preds => place_317_preds,
      succs => place_317_succs,
      token => place_317_token,
      clk   => clk,
      reset => reset);

  place_318_preds(0) <= transition_314_symbol_out;
  place_318_succs(0) <= transition_315_symbol_out;
  place_318 : place
    generic map(marking => false)
    port map(
      preds => place_318_preds,
      succs => place_318_succs,
      token => place_318_token,
      clk   => clk,
      reset => reset);

  place_324_preds(0) <= transition_320_symbol_out;
  place_324_succs(0) <= transition_321_symbol_out;
  place_324 : place
    generic map(marking => false)
    port map(
      preds => place_324_preds,
      succs => place_324_succs,
      token => place_324_token,
      clk   => clk,
      reset => reset);

  place_325_preds(0) <= transition_321_symbol_out;
  place_325_succs(0) <= transition_322_symbol_out;
  place_325 : place
    generic map(marking => false)
    port map(
      preds => place_325_preds,
      succs => place_325_succs,
      token => place_325_token,
      clk   => clk,
      reset => reset);

  place_326_preds(0) <= transition_322_symbol_out;
  place_326_succs(0) <= transition_323_symbol_out;
  place_326 : place
    generic map(marking => false)
    port map(
      preds => place_326_preds,
      succs => place_326_succs,
      token => place_326_token,
      clk   => clk,
      reset => reset);

  place_327_preds(0) <= transition_329_symbol_out;
  place_327_succs(0) <= transition_328_symbol_out;
  place_327 : place
    generic map(marking => false)
    port map(
      preds => place_327_preds,
      succs => place_327_succs,
      token => place_327_token,
      clk   => clk,
      reset => reset);

  place_336_preds(0) <= transition_332_symbol_out;
  place_336_succs(0) <= transition_333_symbol_out;
  place_336 : place
    generic map(marking => false)
    port map(
      preds => place_336_preds,
      succs => place_336_succs,
      token => place_336_token,
      clk   => clk,
      reset => reset);

  place_337_preds(0) <= transition_333_symbol_out;
  place_337_succs(0) <= transition_334_symbol_out;
  place_337 : place
    generic map(marking => false)
    port map(
      preds => place_337_preds,
      succs => place_337_succs,
      token => place_337_token,
      clk   => clk,
      reset => reset);

  place_338_preds(0) <= transition_334_symbol_out;
  place_338_succs(0) <= transition_335_symbol_out;
  place_338 : place
    generic map(marking => false)
    port map(
      preds => place_338_preds,
      succs => place_338_succs,
      token => place_338_token,
      clk   => clk,
      reset => reset);

  place_343_preds(0) <= transition_339_symbol_out;
  place_343_succs(0) <= transition_340_symbol_out;
  place_343 : place
    generic map(marking => false)
    port map(
      preds => place_343_preds,
      succs => place_343_succs,
      token => place_343_token,
      clk   => clk,
      reset => reset);

  place_344_preds(0) <= transition_340_symbol_out;
  place_344_succs(0) <= transition_341_symbol_out;
  place_344 : place
    generic map(marking => false)
    port map(
      preds => place_344_preds,
      succs => place_344_succs,
      token => place_344_token,
      clk   => clk,
      reset => reset);

  place_345_preds(0) <= transition_341_symbol_out;
  place_345_succs(0) <= transition_342_symbol_out;
  place_345 : place
    generic map(marking => false)
    port map(
      preds => place_345_preds,
      succs => place_345_succs,
      token => place_345_token,
      clk   => clk,
      reset => reset);

  place_350_preds(0) <= transition_346_symbol_out;
  place_350_succs(0) <= transition_347_symbol_out;
  place_350 : place
    generic map(marking => false)
    port map(
      preds => place_350_preds,
      succs => place_350_succs,
      token => place_350_token,
      clk   => clk,
      reset => reset);

  place_351_preds(0) <= transition_347_symbol_out;
  place_351_succs(0) <= transition_348_symbol_out;
  place_351 : place
    generic map(marking => false)
    port map(
      preds => place_351_preds,
      succs => place_351_succs,
      token => place_351_token,
      clk   => clk,
      reset => reset);

  place_352_preds(0) <= transition_348_symbol_out;
  place_352_succs(0) <= transition_349_symbol_out;
  place_352 : place
    generic map(marking => false)
    port map(
      preds => place_352_preds,
      succs => place_352_succs,
      token => place_352_token,
      clk   => clk,
      reset => reset);

  place_358_preds(0) <= transition_354_symbol_out;
  place_358_succs(0) <= transition_355_symbol_out;
  place_358 : place
    generic map(marking => false)
    port map(
      preds => place_358_preds,
      succs => place_358_succs,
      token => place_358_token,
      clk   => clk,
      reset => reset);

  place_359_preds(0) <= transition_355_symbol_out;
  place_359_succs(0) <= transition_356_symbol_out;
  place_359 : place
    generic map(marking => false)
    port map(
      preds => place_359_preds,
      succs => place_359_succs,
      token => place_359_token,
      clk   => clk,
      reset => reset);

  place_360_preds(0) <= transition_356_symbol_out;
  place_360_succs(0) <= transition_357_symbol_out;
  place_360 : place
    generic map(marking => false)
    port map(
      preds => place_360_preds,
      succs => place_360_succs,
      token => place_360_token,
      clk   => clk,
      reset => reset);

  place_365_preds(0) <= transition_361_symbol_out;
  place_365_succs(0) <= transition_362_symbol_out;
  place_365 : place
    generic map(marking => false)
    port map(
      preds => place_365_preds,
      succs => place_365_succs,
      token => place_365_token,
      clk   => clk,
      reset => reset);

  place_366_preds(0) <= transition_362_symbol_out;
  place_366_succs(0) <= transition_363_symbol_out;
  place_366 : place
    generic map(marking => false)
    port map(
      preds => place_366_preds,
      succs => place_366_succs,
      token => place_366_token,
      clk   => clk,
      reset => reset);

  place_367_preds(0) <= transition_363_symbol_out;
  place_367_succs(0) <= transition_364_symbol_out;
  place_367 : place
    generic map(marking => false)
    port map(
      preds => place_367_preds,
      succs => place_367_succs,
      token => place_367_token,
      clk   => clk,
      reset => reset);

  place_373_preds(0) <= transition_369_symbol_out;
  place_373_succs(0) <= transition_370_symbol_out;
  place_373 : place
    generic map(marking => false)
    port map(
      preds => place_373_preds,
      succs => place_373_succs,
      token => place_373_token,
      clk   => clk,
      reset => reset);

  place_374_preds(0) <= transition_370_symbol_out;
  place_374_succs(0) <= transition_371_symbol_out;
  place_374 : place
    generic map(marking => false)
    port map(
      preds => place_374_preds,
      succs => place_374_succs,
      token => place_374_token,
      clk   => clk,
      reset => reset);

  place_375_preds(0) <= transition_371_symbol_out;
  place_375_succs(0) <= transition_372_symbol_out;
  place_375 : place
    generic map(marking => false)
    port map(
      preds => place_375_preds,
      succs => place_375_succs,
      token => place_375_token,
      clk   => clk,
      reset => reset);

  place_376_preds(0) <= transition_378_symbol_out;
  place_376_succs(0) <= transition_377_symbol_out;
  place_376 : place
    generic map(marking => false)
    port map(
      preds => place_376_preds,
      succs => place_376_succs,
      token => place_376_token,
      clk   => clk,
      reset => reset);

  place_380_preds(0) <= transition_382_symbol_out;
  place_380_succs(0) <= transition_381_symbol_out;
  place_380 : place
    generic map(marking => false)
    port map(
      preds => place_380_preds,
      succs => place_380_succs,
      token => place_380_token,
      clk   => clk,
      reset => reset);

  place_388_preds(0) <= transition_384_symbol_out;
  place_388_succs(0) <= transition_385_symbol_out;
  place_388 : place
    generic map(marking => false)
    port map(
      preds => place_388_preds,
      succs => place_388_succs,
      token => place_388_token,
      clk   => clk,
      reset => reset);

  place_389_preds(0) <= transition_385_symbol_out;
  place_389_succs(0) <= transition_386_symbol_out;
  place_389 : place
    generic map(marking => false)
    port map(
      preds => place_389_preds,
      succs => place_389_succs,
      token => place_389_token,
      clk   => clk,
      reset => reset);

  place_390_preds(0) <= transition_386_symbol_out;
  place_390_succs(0) <= transition_387_symbol_out;
  place_390 : place
    generic map(marking => false)
    port map(
      preds => place_390_preds,
      succs => place_390_succs,
      token => place_390_token,
      clk   => clk,
      reset => reset);

  place_395_preds(0) <= transition_391_symbol_out;
  place_395_succs(0) <= transition_392_symbol_out;
  place_395 : place
    generic map(marking => false)
    port map(
      preds => place_395_preds,
      succs => place_395_succs,
      token => place_395_token,
      clk   => clk,
      reset => reset);

  place_396_preds(0) <= transition_392_symbol_out;
  place_396_succs(0) <= transition_393_symbol_out;
  place_396 : place
    generic map(marking => false)
    port map(
      preds => place_396_preds,
      succs => place_396_succs,
      token => place_396_token,
      clk   => clk,
      reset => reset);

  place_397_preds(0) <= transition_393_symbol_out;
  place_397_succs(0) <= transition_394_symbol_out;
  place_397 : place
    generic map(marking => false)
    port map(
      preds => place_397_preds,
      succs => place_397_succs,
      token => place_397_token,
      clk   => clk,
      reset => reset);

  place_402_preds(0) <= transition_398_symbol_out;
  place_402_succs(0) <= transition_399_symbol_out;
  place_402 : place
    generic map(marking => false)
    port map(
      preds => place_402_preds,
      succs => place_402_succs,
      token => place_402_token,
      clk   => clk,
      reset => reset);

  place_403_preds(0) <= transition_399_symbol_out;
  place_403_succs(0) <= transition_400_symbol_out;
  place_403 : place
    generic map(marking => false)
    port map(
      preds => place_403_preds,
      succs => place_403_succs,
      token => place_403_token,
      clk   => clk,
      reset => reset);

  place_404_preds(0) <= transition_400_symbol_out;
  place_404_succs(0) <= transition_401_symbol_out;
  place_404 : place
    generic map(marking => false)
    port map(
      preds => place_404_preds,
      succs => place_404_succs,
      token => place_404_token,
      clk   => clk,
      reset => reset);

  place_410_preds(0) <= transition_406_symbol_out;
  place_410_succs(0) <= transition_407_symbol_out;
  place_410 : place
    generic map(marking => false)
    port map(
      preds => place_410_preds,
      succs => place_410_succs,
      token => place_410_token,
      clk   => clk,
      reset => reset);

  place_411_preds(0) <= transition_407_symbol_out;
  place_411_succs(0) <= transition_408_symbol_out;
  place_411 : place
    generic map(marking => false)
    port map(
      preds => place_411_preds,
      succs => place_411_succs,
      token => place_411_token,
      clk   => clk,
      reset => reset);

  place_412_preds(0) <= transition_408_symbol_out;
  place_412_succs(0) <= transition_409_symbol_out;
  place_412 : place
    generic map(marking => false)
    port map(
      preds => place_412_preds,
      succs => place_412_succs,
      token => place_412_token,
      clk   => clk,
      reset => reset);

  place_417_preds(0) <= transition_413_symbol_out;
  place_417_succs(0) <= transition_414_symbol_out;
  place_417 : place
    generic map(marking => false)
    port map(
      preds => place_417_preds,
      succs => place_417_succs,
      token => place_417_token,
      clk   => clk,
      reset => reset);

  place_418_preds(0) <= transition_414_symbol_out;
  place_418_succs(0) <= transition_415_symbol_out;
  place_418 : place
    generic map(marking => false)
    port map(
      preds => place_418_preds,
      succs => place_418_succs,
      token => place_418_token,
      clk   => clk,
      reset => reset);

  place_419_preds(0) <= transition_415_symbol_out;
  place_419_succs(0) <= transition_416_symbol_out;
  place_419 : place
    generic map(marking => false)
    port map(
      preds => place_419_preds,
      succs => place_419_succs,
      token => place_419_token,
      clk   => clk,
      reset => reset);

  place_425_preds(0) <= transition_421_symbol_out;
  place_425_succs(0) <= transition_422_symbol_out;
  place_425 : place
    generic map(marking => false)
    port map(
      preds => place_425_preds,
      succs => place_425_succs,
      token => place_425_token,
      clk   => clk,
      reset => reset);

  place_426_preds(0) <= transition_422_symbol_out;
  place_426_succs(0) <= transition_423_symbol_out;
  place_426 : place
    generic map(marking => false)
    port map(
      preds => place_426_preds,
      succs => place_426_succs,
      token => place_426_token,
      clk   => clk,
      reset => reset);

  place_427_preds(0) <= transition_423_symbol_out;
  place_427_succs(0) <= transition_424_symbol_out;
  place_427 : place
    generic map(marking => false)
    port map(
      preds => place_427_preds,
      succs => place_427_succs,
      token => place_427_token,
      clk   => clk,
      reset => reset);

  place_428_preds(0) <= transition_430_symbol_out;
  place_428_succs(0) <= transition_429_symbol_out;
  place_428 : place
    generic map(marking => false)
    port map(
      preds => place_428_preds,
      succs => place_428_succs,
      token => place_428_token,
      clk   => clk,
      reset => reset);

  place_432_preds(0) <= transition_434_symbol_out;
  place_432_succs(0) <= transition_433_symbol_out;
  place_432 : place
    generic map(marking => false)
    port map(
      preds => place_432_preds,
      succs => place_432_succs,
      token => place_432_token,
      clk   => clk,
      reset => reset);

  place_440_preds(0) <= transition_436_symbol_out;
  place_440_succs(0) <= transition_437_symbol_out;
  place_440 : place
    generic map(marking => false)
    port map(
      preds => place_440_preds,
      succs => place_440_succs,
      token => place_440_token,
      clk   => clk,
      reset => reset);

  place_441_preds(0) <= transition_437_symbol_out;
  place_441_succs(0) <= transition_438_symbol_out;
  place_441 : place
    generic map(marking => false)
    port map(
      preds => place_441_preds,
      succs => place_441_succs,
      token => place_441_token,
      clk   => clk,
      reset => reset);

  place_442_preds(0) <= transition_438_symbol_out;
  place_442_succs(0) <= transition_439_symbol_out;
  place_442 : place
    generic map(marking => false)
    port map(
      preds => place_442_preds,
      succs => place_442_succs,
      token => place_442_token,
      clk   => clk,
      reset => reset);

  place_449_preds(0) <= transition_445_symbol_out;
  place_449_succs(0) <= transition_446_symbol_out;
  place_449 : place
    generic map(marking => false)
    port map(
      preds => place_449_preds,
      succs => place_449_succs,
      token => place_449_token,
      clk   => clk,
      reset => reset);

  place_450_preds(0) <= transition_446_symbol_out;
  place_450_succs(0) <= transition_447_symbol_out;
  place_450 : place
    generic map(marking => false)
    port map(
      preds => place_450_preds,
      succs => place_450_succs,
      token => place_450_token,
      clk   => clk,
      reset => reset);

  place_451_preds(0) <= transition_447_symbol_out;
  place_451_succs(0) <= transition_448_symbol_out;
  place_451 : place
    generic map(marking => false)
    port map(
      preds => place_451_preds,
      succs => place_451_succs,
      token => place_451_token,
      clk   => clk,
      reset => reset);

  place_456_preds(0) <= transition_452_symbol_out;
  place_456_succs(0) <= transition_453_symbol_out;
  place_456 : place
    generic map(marking => false)
    port map(
      preds => place_456_preds,
      succs => place_456_succs,
      token => place_456_token,
      clk   => clk,
      reset => reset);

  place_457_preds(0) <= transition_453_symbol_out;
  place_457_succs(0) <= transition_454_symbol_out;
  place_457 : place
    generic map(marking => false)
    port map(
      preds => place_457_preds,
      succs => place_457_succs,
      token => place_457_token,
      clk   => clk,
      reset => reset);

  place_458_preds(0) <= transition_454_symbol_out;
  place_458_succs(0) <= transition_455_symbol_out;
  place_458 : place
    generic map(marking => false)
    port map(
      preds => place_458_preds,
      succs => place_458_succs,
      token => place_458_token,
      clk   => clk,
      reset => reset);

  place_463_preds(0) <= transition_459_symbol_out;
  place_463_succs(0) <= transition_460_symbol_out;
  place_463 : place
    generic map(marking => false)
    port map(
      preds => place_463_preds,
      succs => place_463_succs,
      token => place_463_token,
      clk   => clk,
      reset => reset);

  place_464_preds(0) <= transition_460_symbol_out;
  place_464_succs(0) <= transition_461_symbol_out;
  place_464 : place
    generic map(marking => false)
    port map(
      preds => place_464_preds,
      succs => place_464_succs,
      token => place_464_token,
      clk   => clk,
      reset => reset);

  place_465_preds(0) <= transition_461_symbol_out;
  place_465_succs(0) <= transition_462_symbol_out;
  place_465 : place
    generic map(marking => false)
    port map(
      preds => place_465_preds,
      succs => place_465_succs,
      token => place_465_token,
      clk   => clk,
      reset => reset);

  place_471_preds(0) <= transition_467_symbol_out;
  place_471_succs(0) <= transition_468_symbol_out;
  place_471 : place
    generic map(marking => false)
    port map(
      preds => place_471_preds,
      succs => place_471_succs,
      token => place_471_token,
      clk   => clk,
      reset => reset);

  place_472_preds(0) <= transition_468_symbol_out;
  place_472_succs(0) <= transition_469_symbol_out;
  place_472 : place
    generic map(marking => false)
    port map(
      preds => place_472_preds,
      succs => place_472_succs,
      token => place_472_token,
      clk   => clk,
      reset => reset);

  place_473_preds(0) <= transition_469_symbol_out;
  place_473_succs(0) <= transition_470_symbol_out;
  place_473 : place
    generic map(marking => false)
    port map(
      preds => place_473_preds,
      succs => place_473_succs,
      token => place_473_token,
      clk   => clk,
      reset => reset);

  place_478_preds(0) <= transition_474_symbol_out;
  place_478_succs(0) <= transition_475_symbol_out;
  place_478 : place
    generic map(marking => false)
    port map(
      preds => place_478_preds,
      succs => place_478_succs,
      token => place_478_token,
      clk   => clk,
      reset => reset);

  place_479_preds(0) <= transition_475_symbol_out;
  place_479_succs(0) <= transition_476_symbol_out;
  place_479 : place
    generic map(marking => false)
    port map(
      preds => place_479_preds,
      succs => place_479_succs,
      token => place_479_token,
      clk   => clk,
      reset => reset);

  place_480_preds(0) <= transition_476_symbol_out;
  place_480_succs(0) <= transition_477_symbol_out;
  place_480 : place
    generic map(marking => false)
    port map(
      preds => place_480_preds,
      succs => place_480_succs,
      token => place_480_token,
      clk   => clk,
      reset => reset);

  place_486_preds(0) <= transition_482_symbol_out;
  place_486_succs(0) <= transition_483_symbol_out;
  place_486 : place
    generic map(marking => false)
    port map(
      preds => place_486_preds,
      succs => place_486_succs,
      token => place_486_token,
      clk   => clk,
      reset => reset);

  place_487_preds(0) <= transition_483_symbol_out;
  place_487_succs(0) <= transition_484_symbol_out;
  place_487 : place
    generic map(marking => false)
    port map(
      preds => place_487_preds,
      succs => place_487_succs,
      token => place_487_token,
      clk   => clk,
      reset => reset);

  place_488_preds(0) <= transition_484_symbol_out;
  place_488_succs(0) <= transition_485_symbol_out;
  place_488 : place
    generic map(marking => false)
    port map(
      preds => place_488_preds,
      succs => place_488_succs,
      token => place_488_token,
      clk   => clk,
      reset => reset);

  place_489_preds(0) <= transition_491_symbol_out;
  place_489_succs(0) <= transition_490_symbol_out;
  place_489 : place
    generic map(marking => false)
    port map(
      preds => place_489_preds,
      succs => place_489_succs,
      token => place_489_token,
      clk   => clk,
      reset => reset);

  place_497_preds(0) <= transition_493_symbol_out;
  place_497_succs(0) <= transition_494_symbol_out;
  place_497 : place
    generic map(marking => false)
    port map(
      preds => place_497_preds,
      succs => place_497_succs,
      token => place_497_token,
      clk   => clk,
      reset => reset);

  place_498_preds(0) <= transition_494_symbol_out;
  place_498_succs(0) <= transition_495_symbol_out;
  place_498 : place
    generic map(marking => false)
    port map(
      preds => place_498_preds,
      succs => place_498_succs,
      token => place_498_token,
      clk   => clk,
      reset => reset);

  place_499_preds(0) <= transition_495_symbol_out;
  place_499_succs(0) <= transition_496_symbol_out;
  place_499 : place
    generic map(marking => false)
    port map(
      preds => place_499_preds,
      succs => place_499_succs,
      token => place_499_token,
      clk   => clk,
      reset => reset);

  place_505_preds(0) <= transition_501_symbol_out;
  place_505_succs(0) <= transition_502_symbol_out;
  place_505 : place
    generic map(marking => false)
    port map(
      preds => place_505_preds,
      succs => place_505_succs,
      token => place_505_token,
      clk   => clk,
      reset => reset);

  place_506_preds(0) <= transition_502_symbol_out;
  place_506_succs(0) <= transition_503_symbol_out;
  place_506 : place
    generic map(marking => false)
    port map(
      preds => place_506_preds,
      succs => place_506_succs,
      token => place_506_token,
      clk   => clk,
      reset => reset);

  place_507_preds(0) <= transition_503_symbol_out;
  place_507_succs(0) <= transition_504_symbol_out;
  place_507 : place
    generic map(marking => false)
    port map(
      preds => place_507_preds,
      succs => place_507_succs,
      token => place_507_token,
      clk   => clk,
      reset => reset);

  place_512_preds(0) <= transition_508_symbol_out;
  place_512_succs(0) <= transition_509_symbol_out;
  place_512 : place
    generic map(marking => false)
    port map(
      preds => place_512_preds,
      succs => place_512_succs,
      token => place_512_token,
      clk   => clk,
      reset => reset);

  place_513_preds(0) <= transition_509_symbol_out;
  place_513_succs(0) <= transition_510_symbol_out;
  place_513 : place
    generic map(marking => false)
    port map(
      preds => place_513_preds,
      succs => place_513_succs,
      token => place_513_token,
      clk   => clk,
      reset => reset);

  place_514_preds(0) <= transition_510_symbol_out;
  place_514_succs(0) <= transition_511_symbol_out;
  place_514 : place
    generic map(marking => false)
    port map(
      preds => place_514_preds,
      succs => place_514_succs,
      token => place_514_token,
      clk   => clk,
      reset => reset);

  place_519_preds(0) <= transition_515_symbol_out;
  place_519_succs(0) <= transition_516_symbol_out;
  place_519 : place
    generic map(marking => false)
    port map(
      preds => place_519_preds,
      succs => place_519_succs,
      token => place_519_token,
      clk   => clk,
      reset => reset);

  place_520_preds(0) <= transition_516_symbol_out;
  place_520_succs(0) <= transition_517_symbol_out;
  place_520 : place
    generic map(marking => false)
    port map(
      preds => place_520_preds,
      succs => place_520_succs,
      token => place_520_token,
      clk   => clk,
      reset => reset);

  place_521_preds(0) <= transition_517_symbol_out;
  place_521_succs(0) <= transition_518_symbol_out;
  place_521 : place
    generic map(marking => false)
    port map(
      preds => place_521_preds,
      succs => place_521_succs,
      token => place_521_token,
      clk   => clk,
      reset => reset);

  place_526_preds(0) <= transition_522_symbol_out;
  place_526_succs(0) <= transition_523_symbol_out;
  place_526 : place
    generic map(marking => false)
    port map(
      preds => place_526_preds,
      succs => place_526_succs,
      token => place_526_token,
      clk   => clk,
      reset => reset);

  place_527_preds(0) <= transition_523_symbol_out;
  place_527_succs(0) <= transition_524_symbol_out;
  place_527 : place
    generic map(marking => false)
    port map(
      preds => place_527_preds,
      succs => place_527_succs,
      token => place_527_token,
      clk   => clk,
      reset => reset);

  place_528_preds(0) <= transition_524_symbol_out;
  place_528_succs(0) <= transition_525_symbol_out;
  place_528 : place
    generic map(marking => false)
    port map(
      preds => place_528_preds,
      succs => place_528_succs,
      token => place_528_token,
      clk   => clk,
      reset => reset);

  place_534_preds(0) <= transition_530_symbol_out;
  place_534_succs(0) <= transition_531_symbol_out;
  place_534 : place
    generic map(marking => false)
    port map(
      preds => place_534_preds,
      succs => place_534_succs,
      token => place_534_token,
      clk   => clk,
      reset => reset);

  place_535_preds(0) <= transition_531_symbol_out;
  place_535_succs(0) <= transition_532_symbol_out;
  place_535 : place
    generic map(marking => false)
    port map(
      preds => place_535_preds,
      succs => place_535_succs,
      token => place_535_token,
      clk   => clk,
      reset => reset);

  place_536_preds(0) <= transition_532_symbol_out;
  place_536_succs(0) <= transition_533_symbol_out;
  place_536 : place
    generic map(marking => false)
    port map(
      preds => place_536_preds,
      succs => place_536_succs,
      token => place_536_token,
      clk   => clk,
      reset => reset);

  place_541_preds(0) <= transition_537_symbol_out;
  place_541_succs(0) <= transition_538_symbol_out;
  place_541 : place
    generic map(marking => false)
    port map(
      preds => place_541_preds,
      succs => place_541_succs,
      token => place_541_token,
      clk   => clk,
      reset => reset);

  place_542_preds(0) <= transition_538_symbol_out;
  place_542_succs(0) <= transition_539_symbol_out;
  place_542 : place
    generic map(marking => false)
    port map(
      preds => place_542_preds,
      succs => place_542_succs,
      token => place_542_token,
      clk   => clk,
      reset => reset);

  place_543_preds(0) <= transition_539_symbol_out;
  place_543_succs(0) <= transition_540_symbol_out;
  place_543 : place
    generic map(marking => false)
    port map(
      preds => place_543_preds,
      succs => place_543_succs,
      token => place_543_token,
      clk   => clk,
      reset => reset);

  place_549_preds(0) <= transition_545_symbol_out;
  place_549_succs(0) <= transition_546_symbol_out;
  place_549 : place
    generic map(marking => false)
    port map(
      preds => place_549_preds,
      succs => place_549_succs,
      token => place_549_token,
      clk   => clk,
      reset => reset);

  place_550_preds(0) <= transition_546_symbol_out;
  place_550_succs(0) <= transition_547_symbol_out;
  place_550 : place
    generic map(marking => false)
    port map(
      preds => place_550_preds,
      succs => place_550_succs,
      token => place_550_token,
      clk   => clk,
      reset => reset);

  place_551_preds(0) <= transition_547_symbol_out;
  place_551_succs(0) <= transition_548_symbol_out;
  place_551 : place
    generic map(marking => false)
    port map(
      preds => place_551_preds,
      succs => place_551_succs,
      token => place_551_token,
      clk   => clk,
      reset => reset);

  place_552_preds(0) <= transition_554_symbol_out;
  place_552_succs(0) <= transition_553_symbol_out;
  place_552 : place
    generic map(marking => false)
    port map(
      preds => place_552_preds,
      succs => place_552_succs,
      token => place_552_token,
      clk   => clk,
      reset => reset);

  place_560_preds(0) <= transition_556_symbol_out;
  place_560_succs(0) <= transition_557_symbol_out;
  place_560 : place
    generic map(marking => false)
    port map(
      preds => place_560_preds,
      succs => place_560_succs,
      token => place_560_token,
      clk   => clk,
      reset => reset);

  place_561_preds(0) <= transition_557_symbol_out;
  place_561_succs(0) <= transition_558_symbol_out;
  place_561 : place
    generic map(marking => false)
    port map(
      preds => place_561_preds,
      succs => place_561_succs,
      token => place_561_token,
      clk   => clk,
      reset => reset);

  place_562_preds(0) <= transition_558_symbol_out;
  place_562_succs(0) <= transition_559_symbol_out;
  place_562 : place
    generic map(marking => false)
    port map(
      preds => place_562_preds,
      succs => place_562_succs,
      token => place_562_token,
      clk   => clk,
      reset => reset);

  place_568_preds(0) <= transition_564_symbol_out;
  place_568_succs(0) <= transition_565_symbol_out;
  place_568 : place
    generic map(marking => false)
    port map(
      preds => place_568_preds,
      succs => place_568_succs,
      token => place_568_token,
      clk   => clk,
      reset => reset);

  place_569_preds(0) <= transition_565_symbol_out;
  place_569_succs(0) <= transition_566_symbol_out;
  place_569 : place
    generic map(marking => false)
    port map(
      preds => place_569_preds,
      succs => place_569_succs,
      token => place_569_token,
      clk   => clk,
      reset => reset);

  place_570_preds(0) <= transition_566_symbol_out;
  place_570_succs(0) <= transition_567_symbol_out;
  place_570 : place
    generic map(marking => false)
    port map(
      preds => place_570_preds,
      succs => place_570_succs,
      token => place_570_token,
      clk   => clk,
      reset => reset);

  place_575_preds(0) <= transition_571_symbol_out;
  place_575_succs(0) <= transition_572_symbol_out;
  place_575 : place
    generic map(marking => false)
    port map(
      preds => place_575_preds,
      succs => place_575_succs,
      token => place_575_token,
      clk   => clk,
      reset => reset);

  place_576_preds(0) <= transition_572_symbol_out;
  place_576_succs(0) <= transition_573_symbol_out;
  place_576 : place
    generic map(marking => false)
    port map(
      preds => place_576_preds,
      succs => place_576_succs,
      token => place_576_token,
      clk   => clk,
      reset => reset);

  place_577_preds(0) <= transition_573_symbol_out;
  place_577_succs(0) <= transition_574_symbol_out;
  place_577 : place
    generic map(marking => false)
    port map(
      preds => place_577_preds,
      succs => place_577_succs,
      token => place_577_token,
      clk   => clk,
      reset => reset);

  place_582_preds(0) <= transition_578_symbol_out;
  place_582_succs(0) <= transition_579_symbol_out;
  place_582 : place
    generic map(marking => false)
    port map(
      preds => place_582_preds,
      succs => place_582_succs,
      token => place_582_token,
      clk   => clk,
      reset => reset);

  place_583_preds(0) <= transition_579_symbol_out;
  place_583_succs(0) <= transition_580_symbol_out;
  place_583 : place
    generic map(marking => false)
    port map(
      preds => place_583_preds,
      succs => place_583_succs,
      token => place_583_token,
      clk   => clk,
      reset => reset);

  place_584_preds(0) <= transition_580_symbol_out;
  place_584_succs(0) <= transition_581_symbol_out;
  place_584 : place
    generic map(marking => false)
    port map(
      preds => place_584_preds,
      succs => place_584_succs,
      token => place_584_token,
      clk   => clk,
      reset => reset);

  place_589_preds(0) <= transition_585_symbol_out;
  place_589_succs(0) <= transition_586_symbol_out;
  place_589 : place
    generic map(marking => false)
    port map(
      preds => place_589_preds,
      succs => place_589_succs,
      token => place_589_token,
      clk   => clk,
      reset => reset);

  place_590_preds(0) <= transition_586_symbol_out;
  place_590_succs(0) <= transition_587_symbol_out;
  place_590 : place
    generic map(marking => false)
    port map(
      preds => place_590_preds,
      succs => place_590_succs,
      token => place_590_token,
      clk   => clk,
      reset => reset);

  place_591_preds(0) <= transition_587_symbol_out;
  place_591_succs(0) <= transition_588_symbol_out;
  place_591 : place
    generic map(marking => false)
    port map(
      preds => place_591_preds,
      succs => place_591_succs,
      token => place_591_token,
      clk   => clk,
      reset => reset);

  place_597_preds(0) <= transition_593_symbol_out;
  place_597_succs(0) <= transition_594_symbol_out;
  place_597 : place
    generic map(marking => false)
    port map(
      preds => place_597_preds,
      succs => place_597_succs,
      token => place_597_token,
      clk   => clk,
      reset => reset);

  place_598_preds(0) <= transition_594_symbol_out;
  place_598_succs(0) <= transition_595_symbol_out;
  place_598 : place
    generic map(marking => false)
    port map(
      preds => place_598_preds,
      succs => place_598_succs,
      token => place_598_token,
      clk   => clk,
      reset => reset);

  place_599_preds(0) <= transition_595_symbol_out;
  place_599_succs(0) <= transition_596_symbol_out;
  place_599 : place
    generic map(marking => false)
    port map(
      preds => place_599_preds,
      succs => place_599_succs,
      token => place_599_token,
      clk   => clk,
      reset => reset);

  place_604_preds(0) <= transition_600_symbol_out;
  place_604_succs(0) <= transition_601_symbol_out;
  place_604 : place
    generic map(marking => false)
    port map(
      preds => place_604_preds,
      succs => place_604_succs,
      token => place_604_token,
      clk   => clk,
      reset => reset);

  place_605_preds(0) <= transition_601_symbol_out;
  place_605_succs(0) <= transition_602_symbol_out;
  place_605 : place
    generic map(marking => false)
    port map(
      preds => place_605_preds,
      succs => place_605_succs,
      token => place_605_token,
      clk   => clk,
      reset => reset);

  place_606_preds(0) <= transition_602_symbol_out;
  place_606_succs(0) <= transition_603_symbol_out;
  place_606 : place
    generic map(marking => false)
    port map(
      preds => place_606_preds,
      succs => place_606_succs,
      token => place_606_token,
      clk   => clk,
      reset => reset);

  place_612_preds(0) <= transition_608_symbol_out;
  place_612_succs(0) <= transition_609_symbol_out;
  place_612 : place
    generic map(marking => false)
    port map(
      preds => place_612_preds,
      succs => place_612_succs,
      token => place_612_token,
      clk   => clk,
      reset => reset);

  place_613_preds(0) <= transition_609_symbol_out;
  place_613_succs(0) <= transition_610_symbol_out;
  place_613 : place
    generic map(marking => false)
    port map(
      preds => place_613_preds,
      succs => place_613_succs,
      token => place_613_token,
      clk   => clk,
      reset => reset);

  place_614_preds(0) <= transition_610_symbol_out;
  place_614_succs(0) <= transition_611_symbol_out;
  place_614 : place
    generic map(marking => false)
    port map(
      preds => place_614_preds,
      succs => place_614_succs,
      token => place_614_token,
      clk   => clk,
      reset => reset);

  place_615_preds(0) <= transition_617_symbol_out;
  place_615_succs(0) <= transition_616_symbol_out;
  place_615 : place
    generic map(marking => false)
    port map(
      preds => place_615_preds,
      succs => place_615_succs,
      token => place_615_token,
      clk   => clk,
      reset => reset);

  place_623_preds(0) <= transition_619_symbol_out;
  place_623_succs(0) <= transition_620_symbol_out;
  place_623 : place
    generic map(marking => false)
    port map(
      preds => place_623_preds,
      succs => place_623_succs,
      token => place_623_token,
      clk   => clk,
      reset => reset);

  place_624_preds(0) <= transition_620_symbol_out;
  place_624_succs(0) <= transition_621_symbol_out;
  place_624 : place
    generic map(marking => false)
    port map(
      preds => place_624_preds,
      succs => place_624_succs,
      token => place_624_token,
      clk   => clk,
      reset => reset);

  place_625_preds(0) <= transition_621_symbol_out;
  place_625_succs(0) <= transition_622_symbol_out;
  place_625 : place
    generic map(marking => false)
    port map(
      preds => place_625_preds,
      succs => place_625_succs,
      token => place_625_token,
      clk   => clk,
      reset => reset);

  place_631_preds(0) <= transition_627_symbol_out;
  place_631_succs(0) <= transition_628_symbol_out;
  place_631 : place
    generic map(marking => false)
    port map(
      preds => place_631_preds,
      succs => place_631_succs,
      token => place_631_token,
      clk   => clk,
      reset => reset);

  place_632_preds(0) <= transition_628_symbol_out;
  place_632_succs(0) <= transition_629_symbol_out;
  place_632 : place
    generic map(marking => false)
    port map(
      preds => place_632_preds,
      succs => place_632_succs,
      token => place_632_token,
      clk   => clk,
      reset => reset);

  place_633_preds(0) <= transition_629_symbol_out;
  place_633_succs(0) <= transition_630_symbol_out;
  place_633 : place
    generic map(marking => false)
    port map(
      preds => place_633_preds,
      succs => place_633_succs,
      token => place_633_token,
      clk   => clk,
      reset => reset);

  place_638_preds(0) <= transition_634_symbol_out;
  place_638_succs(0) <= transition_635_symbol_out;
  place_638 : place
    generic map(marking => false)
    port map(
      preds => place_638_preds,
      succs => place_638_succs,
      token => place_638_token,
      clk   => clk,
      reset => reset);

  place_639_preds(0) <= transition_635_symbol_out;
  place_639_succs(0) <= transition_636_symbol_out;
  place_639 : place
    generic map(marking => false)
    port map(
      preds => place_639_preds,
      succs => place_639_succs,
      token => place_639_token,
      clk   => clk,
      reset => reset);

  place_640_preds(0) <= transition_636_symbol_out;
  place_640_succs(0) <= transition_637_symbol_out;
  place_640 : place
    generic map(marking => false)
    port map(
      preds => place_640_preds,
      succs => place_640_succs,
      token => place_640_token,
      clk   => clk,
      reset => reset);

  place_645_preds(0) <= transition_641_symbol_out;
  place_645_succs(0) <= transition_642_symbol_out;
  place_645 : place
    generic map(marking => false)
    port map(
      preds => place_645_preds,
      succs => place_645_succs,
      token => place_645_token,
      clk   => clk,
      reset => reset);

  place_646_preds(0) <= transition_642_symbol_out;
  place_646_succs(0) <= transition_643_symbol_out;
  place_646 : place
    generic map(marking => false)
    port map(
      preds => place_646_preds,
      succs => place_646_succs,
      token => place_646_token,
      clk   => clk,
      reset => reset);

  place_647_preds(0) <= transition_643_symbol_out;
  place_647_succs(0) <= transition_644_symbol_out;
  place_647 : place
    generic map(marking => false)
    port map(
      preds => place_647_preds,
      succs => place_647_succs,
      token => place_647_token,
      clk   => clk,
      reset => reset);

  place_652_preds(0) <= transition_648_symbol_out;
  place_652_succs(0) <= transition_649_symbol_out;
  place_652 : place
    generic map(marking => false)
    port map(
      preds => place_652_preds,
      succs => place_652_succs,
      token => place_652_token,
      clk   => clk,
      reset => reset);

  place_653_preds(0) <= transition_649_symbol_out;
  place_653_succs(0) <= transition_650_symbol_out;
  place_653 : place
    generic map(marking => false)
    port map(
      preds => place_653_preds,
      succs => place_653_succs,
      token => place_653_token,
      clk   => clk,
      reset => reset);

  place_654_preds(0) <= transition_650_symbol_out;
  place_654_succs(0) <= transition_651_symbol_out;
  place_654 : place
    generic map(marking => false)
    port map(
      preds => place_654_preds,
      succs => place_654_succs,
      token => place_654_token,
      clk   => clk,
      reset => reset);

  place_660_preds(0) <= transition_656_symbol_out;
  place_660_succs(0) <= transition_657_symbol_out;
  place_660 : place
    generic map(marking => false)
    port map(
      preds => place_660_preds,
      succs => place_660_succs,
      token => place_660_token,
      clk   => clk,
      reset => reset);

  place_661_preds(0) <= transition_657_symbol_out;
  place_661_succs(0) <= transition_658_symbol_out;
  place_661 : place
    generic map(marking => false)
    port map(
      preds => place_661_preds,
      succs => place_661_succs,
      token => place_661_token,
      clk   => clk,
      reset => reset);

  place_662_preds(0) <= transition_658_symbol_out;
  place_662_succs(0) <= transition_659_symbol_out;
  place_662 : place
    generic map(marking => false)
    port map(
      preds => place_662_preds,
      succs => place_662_succs,
      token => place_662_token,
      clk   => clk,
      reset => reset);

  place_667_preds(0) <= transition_663_symbol_out;
  place_667_succs(0) <= transition_664_symbol_out;
  place_667 : place
    generic map(marking => false)
    port map(
      preds => place_667_preds,
      succs => place_667_succs,
      token => place_667_token,
      clk   => clk,
      reset => reset);

  place_668_preds(0) <= transition_664_symbol_out;
  place_668_succs(0) <= transition_665_symbol_out;
  place_668 : place
    generic map(marking => false)
    port map(
      preds => place_668_preds,
      succs => place_668_succs,
      token => place_668_token,
      clk   => clk,
      reset => reset);

  place_669_preds(0) <= transition_665_symbol_out;
  place_669_succs(0) <= transition_666_symbol_out;
  place_669 : place
    generic map(marking => false)
    port map(
      preds => place_669_preds,
      succs => place_669_succs,
      token => place_669_token,
      clk   => clk,
      reset => reset);

  place_675_preds(0) <= transition_671_symbol_out;
  place_675_succs(0) <= transition_672_symbol_out;
  place_675 : place
    generic map(marking => false)
    port map(
      preds => place_675_preds,
      succs => place_675_succs,
      token => place_675_token,
      clk   => clk,
      reset => reset);

  place_676_preds(0) <= transition_672_symbol_out;
  place_676_succs(0) <= transition_673_symbol_out;
  place_676 : place
    generic map(marking => false)
    port map(
      preds => place_676_preds,
      succs => place_676_succs,
      token => place_676_token,
      clk   => clk,
      reset => reset);

  place_677_preds(0) <= transition_673_symbol_out;
  place_677_succs(0) <= transition_674_symbol_out;
  place_677 : place
    generic map(marking => false)
    port map(
      preds => place_677_preds,
      succs => place_677_succs,
      token => place_677_token,
      clk   => clk,
      reset => reset);

  place_678_preds(0) <= transition_680_symbol_out;
  place_678_succs(0) <= transition_679_symbol_out;
  place_678 : place
    generic map(marking => false)
    port map(
      preds => place_678_preds,
      succs => place_678_succs,
      token => place_678_token,
      clk   => clk,
      reset => reset);

  place_687_preds(0) <= transition_683_symbol_out;
  place_687_succs(0) <= transition_684_symbol_out;
  place_687 : place
    generic map(marking => false)
    port map(
      preds => place_687_preds,
      succs => place_687_succs,
      token => place_687_token,
      clk   => clk,
      reset => reset);

  place_688_preds(0) <= transition_684_symbol_out;
  place_688_succs(0) <= transition_685_symbol_out;
  place_688 : place
    generic map(marking => false)
    port map(
      preds => place_688_preds,
      succs => place_688_succs,
      token => place_688_token,
      clk   => clk,
      reset => reset);

  place_689_preds(0) <= transition_685_symbol_out;
  place_689_succs(0) <= transition_686_symbol_out;
  place_689 : place
    generic map(marking => false)
    port map(
      preds => place_689_preds,
      succs => place_689_succs,
      token => place_689_token,
      clk   => clk,
      reset => reset);

  place_694_preds(0) <= transition_690_symbol_out;
  place_694_succs(0) <= transition_691_symbol_out;
  place_694 : place
    generic map(marking => false)
    port map(
      preds => place_694_preds,
      succs => place_694_succs,
      token => place_694_token,
      clk   => clk,
      reset => reset);

  place_695_preds(0) <= transition_691_symbol_out;
  place_695_succs(0) <= transition_692_symbol_out;
  place_695 : place
    generic map(marking => false)
    port map(
      preds => place_695_preds,
      succs => place_695_succs,
      token => place_695_token,
      clk   => clk,
      reset => reset);

  place_696_preds(0) <= transition_692_symbol_out;
  place_696_succs(0) <= transition_693_symbol_out;
  place_696 : place
    generic map(marking => false)
    port map(
      preds => place_696_preds,
      succs => place_696_succs,
      token => place_696_token,
      clk   => clk,
      reset => reset);

  place_701_preds(0) <= transition_697_symbol_out;
  place_701_succs(0) <= transition_698_symbol_out;
  place_701 : place
    generic map(marking => false)
    port map(
      preds => place_701_preds,
      succs => place_701_succs,
      token => place_701_token,
      clk   => clk,
      reset => reset);

  place_702_preds(0) <= transition_698_symbol_out;
  place_702_succs(0) <= transition_699_symbol_out;
  place_702 : place
    generic map(marking => false)
    port map(
      preds => place_702_preds,
      succs => place_702_succs,
      token => place_702_token,
      clk   => clk,
      reset => reset);

  place_703_preds(0) <= transition_699_symbol_out;
  place_703_succs(0) <= transition_700_symbol_out;
  place_703 : place
    generic map(marking => false)
    port map(
      preds => place_703_preds,
      succs => place_703_succs,
      token => place_703_token,
      clk   => clk,
      reset => reset);

  place_709_preds(0) <= transition_705_symbol_out;
  place_709_succs(0) <= transition_706_symbol_out;
  place_709 : place
    generic map(marking => false)
    port map(
      preds => place_709_preds,
      succs => place_709_succs,
      token => place_709_token,
      clk   => clk,
      reset => reset);

  place_710_preds(0) <= transition_706_symbol_out;
  place_710_succs(0) <= transition_707_symbol_out;
  place_710 : place
    generic map(marking => false)
    port map(
      preds => place_710_preds,
      succs => place_710_succs,
      token => place_710_token,
      clk   => clk,
      reset => reset);

  place_711_preds(0) <= transition_707_symbol_out;
  place_711_succs(0) <= transition_708_symbol_out;
  place_711 : place
    generic map(marking => false)
    port map(
      preds => place_711_preds,
      succs => place_711_succs,
      token => place_711_token,
      clk   => clk,
      reset => reset);

  place_716_preds(0) <= transition_712_symbol_out;
  place_716_succs(0) <= transition_713_symbol_out;
  place_716 : place
    generic map(marking => false)
    port map(
      preds => place_716_preds,
      succs => place_716_succs,
      token => place_716_token,
      clk   => clk,
      reset => reset);

  place_717_preds(0) <= transition_713_symbol_out;
  place_717_succs(0) <= transition_714_symbol_out;
  place_717 : place
    generic map(marking => false)
    port map(
      preds => place_717_preds,
      succs => place_717_succs,
      token => place_717_token,
      clk   => clk,
      reset => reset);

  place_718_preds(0) <= transition_714_symbol_out;
  place_718_succs(0) <= transition_715_symbol_out;
  place_718 : place
    generic map(marking => false)
    port map(
      preds => place_718_preds,
      succs => place_718_succs,
      token => place_718_token,
      clk   => clk,
      reset => reset);

  place_724_preds(0) <= transition_720_symbol_out;
  place_724_succs(0) <= transition_721_symbol_out;
  place_724 : place
    generic map(marking => false)
    port map(
      preds => place_724_preds,
      succs => place_724_succs,
      token => place_724_token,
      clk   => clk,
      reset => reset);

  place_725_preds(0) <= transition_721_symbol_out;
  place_725_succs(0) <= transition_722_symbol_out;
  place_725 : place
    generic map(marking => false)
    port map(
      preds => place_725_preds,
      succs => place_725_succs,
      token => place_725_token,
      clk   => clk,
      reset => reset);

  place_726_preds(0) <= transition_722_symbol_out;
  place_726_succs(0) <= transition_723_symbol_out;
  place_726 : place
    generic map(marking => false)
    port map(
      preds => place_726_preds,
      succs => place_726_succs,
      token => place_726_token,
      clk   => clk,
      reset => reset);

  place_727_preds(0) <= transition_729_symbol_out;
  place_727_succs(0) <= transition_728_symbol_out;
  place_727 : place
    generic map(marking => false)
    port map(
      preds => place_727_preds,
      succs => place_727_succs,
      token => place_727_token,
      clk   => clk,
      reset => reset);

  place_731_preds(0) <= transition_733_symbol_out;
  place_731_succs(0) <= transition_732_symbol_out;
  place_731 : place
    generic map(marking => false)
    port map(
      preds => place_731_preds,
      succs => place_731_succs,
      token => place_731_token,
      clk   => clk,
      reset => reset);

  place_738_preds(0) <= transition_734_symbol_out;
  place_738_succs(0) <= transition_735_symbol_out;
  place_738 : place
    generic map(marking => false)
    port map(
      preds => place_738_preds,
      succs => place_738_succs,
      token => place_738_token,
      clk   => clk,
      reset => reset);

  place_739_preds(0) <= transition_735_symbol_out;
  place_739_succs(0) <= transition_736_symbol_out;
  place_739 : place
    generic map(marking => false)
    port map(
      preds => place_739_preds,
      succs => place_739_succs,
      token => place_739_token,
      clk   => clk,
      reset => reset);

  place_740_preds(0) <= transition_736_symbol_out;
  place_740_succs(0) <= transition_737_symbol_out;
  place_740 : place
    generic map(marking => false)
    port map(
      preds => place_740_preds,
      succs => place_740_succs,
      token => place_740_token,
      clk   => clk,
      reset => reset);

  place_745_preds(0) <= transition_741_symbol_out;
  place_745_succs(0) <= transition_742_symbol_out;
  place_745 : place
    generic map(marking => false)
    port map(
      preds => place_745_preds,
      succs => place_745_succs,
      token => place_745_token,
      clk   => clk,
      reset => reset);

  place_746_preds(0) <= transition_742_symbol_out;
  place_746_succs(0) <= transition_743_symbol_out;
  place_746 : place
    generic map(marking => false)
    port map(
      preds => place_746_preds,
      succs => place_746_succs,
      token => place_746_token,
      clk   => clk,
      reset => reset);

  place_747_preds(0) <= transition_743_symbol_out;
  place_747_succs(0) <= transition_744_symbol_out;
  place_747 : place
    generic map(marking => false)
    port map(
      preds => place_747_preds,
      succs => place_747_succs,
      token => place_747_token,
      clk   => clk,
      reset => reset);

  place_752_preds(0) <= transition_748_symbol_out;
  place_752_succs(0) <= transition_749_symbol_out;
  place_752 : place
    generic map(marking => false)
    port map(
      preds => place_752_preds,
      succs => place_752_succs,
      token => place_752_token,
      clk   => clk,
      reset => reset);

  place_753_preds(0) <= transition_749_symbol_out;
  place_753_succs(0) <= transition_750_symbol_out;
  place_753 : place
    generic map(marking => false)
    port map(
      preds => place_753_preds,
      succs => place_753_succs,
      token => place_753_token,
      clk   => clk,
      reset => reset);

  place_754_preds(0) <= transition_750_symbol_out;
  place_754_succs(0) <= transition_751_symbol_out;
  place_754 : place
    generic map(marking => false)
    port map(
      preds => place_754_preds,
      succs => place_754_succs,
      token => place_754_token,
      clk   => clk,
      reset => reset);

  place_760_preds(0) <= transition_756_symbol_out;
  place_760_succs(0) <= transition_757_symbol_out;
  place_760 : place
    generic map(marking => false)
    port map(
      preds => place_760_preds,
      succs => place_760_succs,
      token => place_760_token,
      clk   => clk,
      reset => reset);

  place_761_preds(0) <= transition_757_symbol_out;
  place_761_succs(0) <= transition_758_symbol_out;
  place_761 : place
    generic map(marking => false)
    port map(
      preds => place_761_preds,
      succs => place_761_succs,
      token => place_761_token,
      clk   => clk,
      reset => reset);

  place_762_preds(0) <= transition_758_symbol_out;
  place_762_succs(0) <= transition_759_symbol_out;
  place_762 : place
    generic map(marking => false)
    port map(
      preds => place_762_preds,
      succs => place_762_succs,
      token => place_762_token,
      clk   => clk,
      reset => reset);

  place_767_preds(0) <= transition_763_symbol_out;
  place_767_succs(0) <= transition_764_symbol_out;
  place_767 : place
    generic map(marking => false)
    port map(
      preds => place_767_preds,
      succs => place_767_succs,
      token => place_767_token,
      clk   => clk,
      reset => reset);

  place_768_preds(0) <= transition_764_symbol_out;
  place_768_succs(0) <= transition_765_symbol_out;
  place_768 : place
    generic map(marking => false)
    port map(
      preds => place_768_preds,
      succs => place_768_succs,
      token => place_768_token,
      clk   => clk,
      reset => reset);

  place_769_preds(0) <= transition_765_symbol_out;
  place_769_succs(0) <= transition_766_symbol_out;
  place_769 : place
    generic map(marking => false)
    port map(
      preds => place_769_preds,
      succs => place_769_succs,
      token => place_769_token,
      clk   => clk,
      reset => reset);

  place_775_preds(0) <= transition_771_symbol_out;
  place_775_succs(0) <= transition_772_symbol_out;
  place_775 : place
    generic map(marking => false)
    port map(
      preds => place_775_preds,
      succs => place_775_succs,
      token => place_775_token,
      clk   => clk,
      reset => reset);

  place_776_preds(0) <= transition_772_symbol_out;
  place_776_succs(0) <= transition_773_symbol_out;
  place_776 : place
    generic map(marking => false)
    port map(
      preds => place_776_preds,
      succs => place_776_succs,
      token => place_776_token,
      clk   => clk,
      reset => reset);

  place_777_preds(0) <= transition_773_symbol_out;
  place_777_succs(0) <= transition_774_symbol_out;
  place_777 : place
    generic map(marking => false)
    port map(
      preds => place_777_preds,
      succs => place_777_succs,
      token => place_777_token,
      clk   => clk,
      reset => reset);

  place_778_preds(0) <= transition_780_symbol_out;
  place_778_succs(0) <= transition_779_symbol_out;
  place_778 : place
    generic map(marking => false)
    port map(
      preds => place_778_preds,
      succs => place_778_succs,
      token => place_778_token,
      clk   => clk,
      reset => reset);

  place_782_preds(0) <= transition_784_symbol_out;
  place_782_succs(0) <= transition_783_symbol_out;
  place_782 : place
    generic map(marking => false)
    port map(
      preds => place_782_preds,
      succs => place_782_succs,
      token => place_782_token,
      clk   => clk,
      reset => reset);

  place_789_preds(0) <= transition_785_symbol_out;
  place_789_succs(0) <= transition_786_symbol_out;
  place_789 : place
    generic map(marking => false)
    port map(
      preds => place_789_preds,
      succs => place_789_succs,
      token => place_789_token,
      clk   => clk,
      reset => reset);

  place_790_preds(0) <= transition_786_symbol_out;
  place_790_succs(0) <= transition_787_symbol_out;
  place_790 : place
    generic map(marking => false)
    port map(
      preds => place_790_preds,
      succs => place_790_succs,
      token => place_790_token,
      clk   => clk,
      reset => reset);

  place_791_preds(0) <= transition_787_symbol_out;
  place_791_succs(0) <= transition_788_symbol_out;
  place_791 : place
    generic map(marking => false)
    port map(
      preds => place_791_preds,
      succs => place_791_succs,
      token => place_791_token,
      clk   => clk,
      reset => reset);

  place_797_preds(0) <= transition_793_symbol_out;
  place_797_succs(0) <= transition_794_symbol_out;
  place_797 : place
    generic map(marking => false)
    port map(
      preds => place_797_preds,
      succs => place_797_succs,
      token => place_797_token,
      clk   => clk,
      reset => reset);

  place_798_preds(0) <= transition_794_symbol_out;
  place_798_succs(0) <= transition_795_symbol_out;
  place_798 : place
    generic map(marking => false)
    port map(
      preds => place_798_preds,
      succs => place_798_succs,
      token => place_798_token,
      clk   => clk,
      reset => reset);

  place_799_preds(0) <= transition_795_symbol_out;
  place_799_succs(0) <= transition_796_symbol_out;
  place_799 : place
    generic map(marking => false)
    port map(
      preds => place_799_preds,
      succs => place_799_succs,
      token => place_799_token,
      clk   => clk,
      reset => reset);

  place_804_preds(0) <= transition_800_symbol_out;
  place_804_succs(0) <= transition_801_symbol_out;
  place_804 : place
    generic map(marking => false)
    port map(
      preds => place_804_preds,
      succs => place_804_succs,
      token => place_804_token,
      clk   => clk,
      reset => reset);

  place_805_preds(0) <= transition_801_symbol_out;
  place_805_succs(0) <= transition_802_symbol_out;
  place_805 : place
    generic map(marking => false)
    port map(
      preds => place_805_preds,
      succs => place_805_succs,
      token => place_805_token,
      clk   => clk,
      reset => reset);

  place_806_preds(0) <= transition_802_symbol_out;
  place_806_succs(0) <= transition_803_symbol_out;
  place_806 : place
    generic map(marking => false)
    port map(
      preds => place_806_preds,
      succs => place_806_succs,
      token => place_806_token,
      clk   => clk,
      reset => reset);

  place_811_preds(0) <= transition_807_symbol_out;
  place_811_succs(0) <= transition_808_symbol_out;
  place_811 : place
    generic map(marking => false)
    port map(
      preds => place_811_preds,
      succs => place_811_succs,
      token => place_811_token,
      clk   => clk,
      reset => reset);

  place_812_preds(0) <= transition_808_symbol_out;
  place_812_succs(0) <= transition_809_symbol_out;
  place_812 : place
    generic map(marking => false)
    port map(
      preds => place_812_preds,
      succs => place_812_succs,
      token => place_812_token,
      clk   => clk,
      reset => reset);

  place_813_preds(0) <= transition_809_symbol_out;
  place_813_succs(0) <= transition_810_symbol_out;
  place_813 : place
    generic map(marking => false)
    port map(
      preds => place_813_preds,
      succs => place_813_succs,
      token => place_813_token,
      clk   => clk,
      reset => reset);

  place_818_preds(0) <= transition_814_symbol_out;
  place_818_succs(0) <= transition_815_symbol_out;
  place_818 : place
    generic map(marking => false)
    port map(
      preds => place_818_preds,
      succs => place_818_succs,
      token => place_818_token,
      clk   => clk,
      reset => reset);

  place_819_preds(0) <= transition_815_symbol_out;
  place_819_succs(0) <= transition_816_symbol_out;
  place_819 : place
    generic map(marking => false)
    port map(
      preds => place_819_preds,
      succs => place_819_succs,
      token => place_819_token,
      clk   => clk,
      reset => reset);

  place_820_preds(0) <= transition_816_symbol_out;
  place_820_succs(0) <= transition_817_symbol_out;
  place_820 : place
    generic map(marking => false)
    port map(
      preds => place_820_preds,
      succs => place_820_succs,
      token => place_820_token,
      clk   => clk,
      reset => reset);

  place_826_preds(0) <= transition_822_symbol_out;
  place_826_succs(0) <= transition_823_symbol_out;
  place_826 : place
    generic map(marking => false)
    port map(
      preds => place_826_preds,
      succs => place_826_succs,
      token => place_826_token,
      clk   => clk,
      reset => reset);

  place_827_preds(0) <= transition_823_symbol_out;
  place_827_succs(0) <= transition_824_symbol_out;
  place_827 : place
    generic map(marking => false)
    port map(
      preds => place_827_preds,
      succs => place_827_succs,
      token => place_827_token,
      clk   => clk,
      reset => reset);

  place_828_preds(0) <= transition_824_symbol_out;
  place_828_succs(0) <= transition_825_symbol_out;
  place_828 : place
    generic map(marking => false)
    port map(
      preds => place_828_preds,
      succs => place_828_succs,
      token => place_828_token,
      clk   => clk,
      reset => reset);

  place_833_preds(0) <= transition_829_symbol_out;
  place_833_succs(0) <= transition_830_symbol_out;
  place_833 : place
    generic map(marking => false)
    port map(
      preds => place_833_preds,
      succs => place_833_succs,
      token => place_833_token,
      clk   => clk,
      reset => reset);

  place_834_preds(0) <= transition_830_symbol_out;
  place_834_succs(0) <= transition_831_symbol_out;
  place_834 : place
    generic map(marking => false)
    port map(
      preds => place_834_preds,
      succs => place_834_succs,
      token => place_834_token,
      clk   => clk,
      reset => reset);

  place_835_preds(0) <= transition_831_symbol_out;
  place_835_succs(0) <= transition_832_symbol_out;
  place_835 : place
    generic map(marking => false)
    port map(
      preds => place_835_preds,
      succs => place_835_succs,
      token => place_835_token,
      clk   => clk,
      reset => reset);

  place_841_preds(0) <= transition_837_symbol_out;
  place_841_succs(0) <= transition_838_symbol_out;
  place_841 : place
    generic map(marking => false)
    port map(
      preds => place_841_preds,
      succs => place_841_succs,
      token => place_841_token,
      clk   => clk,
      reset => reset);

  place_842_preds(0) <= transition_838_symbol_out;
  place_842_succs(0) <= transition_839_symbol_out;
  place_842 : place
    generic map(marking => false)
    port map(
      preds => place_842_preds,
      succs => place_842_succs,
      token => place_842_token,
      clk   => clk,
      reset => reset);

  place_843_preds(0) <= transition_839_symbol_out;
  place_843_succs(0) <= transition_840_symbol_out;
  place_843 : place
    generic map(marking => false)
    port map(
      preds => place_843_preds,
      succs => place_843_succs,
      token => place_843_token,
      clk   => clk,
      reset => reset);

  place_844_preds(0) <= transition_846_symbol_out;
  place_844_succs(0) <= transition_845_symbol_out;
  place_844 : place
    generic map(marking => false)
    port map(
      preds => place_844_preds,
      succs => place_844_succs,
      token => place_844_token,
      clk   => clk,
      reset => reset);

  place_853_preds(0) <= transition_849_symbol_out;
  place_853_succs(0) <= transition_850_symbol_out;
  place_853 : place
    generic map(marking => false)
    port map(
      preds => place_853_preds,
      succs => place_853_succs,
      token => place_853_token,
      clk   => clk,
      reset => reset);

  place_854_preds(0) <= transition_850_symbol_out;
  place_854_succs(0) <= transition_851_symbol_out;
  place_854 : place
    generic map(marking => false)
    port map(
      preds => place_854_preds,
      succs => place_854_succs,
      token => place_854_token,
      clk   => clk,
      reset => reset);

  place_855_preds(0) <= transition_851_symbol_out;
  place_855_succs(0) <= transition_852_symbol_out;
  place_855 : place
    generic map(marking => false)
    port map(
      preds => place_855_preds,
      succs => place_855_succs,
      token => place_855_token,
      clk   => clk,
      reset => reset);

  place_860_preds(0) <= transition_856_symbol_out;
  place_860_succs(0) <= transition_857_symbol_out;
  place_860 : place
    generic map(marking => false)
    port map(
      preds => place_860_preds,
      succs => place_860_succs,
      token => place_860_token,
      clk   => clk,
      reset => reset);

  place_861_preds(0) <= transition_857_symbol_out;
  place_861_succs(0) <= transition_858_symbol_out;
  place_861 : place
    generic map(marking => false)
    port map(
      preds => place_861_preds,
      succs => place_861_succs,
      token => place_861_token,
      clk   => clk,
      reset => reset);

  place_862_preds(0) <= transition_858_symbol_out;
  place_862_succs(0) <= transition_859_symbol_out;
  place_862 : place
    generic map(marking => false)
    port map(
      preds => place_862_preds,
      succs => place_862_succs,
      token => place_862_token,
      clk   => clk,
      reset => reset);

  place_867_preds(0) <= transition_863_symbol_out;
  place_867_succs(0) <= transition_864_symbol_out;
  place_867 : place
    generic map(marking => false)
    port map(
      preds => place_867_preds,
      succs => place_867_succs,
      token => place_867_token,
      clk   => clk,
      reset => reset);

  place_868_preds(0) <= transition_864_symbol_out;
  place_868_succs(0) <= transition_865_symbol_out;
  place_868 : place
    generic map(marking => false)
    port map(
      preds => place_868_preds,
      succs => place_868_succs,
      token => place_868_token,
      clk   => clk,
      reset => reset);

  place_869_preds(0) <= transition_865_symbol_out;
  place_869_succs(0) <= transition_866_symbol_out;
  place_869 : place
    generic map(marking => false)
    port map(
      preds => place_869_preds,
      succs => place_869_succs,
      token => place_869_token,
      clk   => clk,
      reset => reset);

  place_875_preds(0) <= transition_871_symbol_out;
  place_875_succs(0) <= transition_872_symbol_out;
  place_875 : place
    generic map(marking => false)
    port map(
      preds => place_875_preds,
      succs => place_875_succs,
      token => place_875_token,
      clk   => clk,
      reset => reset);

  place_876_preds(0) <= transition_872_symbol_out;
  place_876_succs(0) <= transition_873_symbol_out;
  place_876 : place
    generic map(marking => false)
    port map(
      preds => place_876_preds,
      succs => place_876_succs,
      token => place_876_token,
      clk   => clk,
      reset => reset);

  place_877_preds(0) <= transition_873_symbol_out;
  place_877_succs(0) <= transition_874_symbol_out;
  place_877 : place
    generic map(marking => false)
    port map(
      preds => place_877_preds,
      succs => place_877_succs,
      token => place_877_token,
      clk   => clk,
      reset => reset);

  place_882_preds(0) <= transition_878_symbol_out;
  place_882_succs(0) <= transition_879_symbol_out;
  place_882 : place
    generic map(marking => false)
    port map(
      preds => place_882_preds,
      succs => place_882_succs,
      token => place_882_token,
      clk   => clk,
      reset => reset);

  place_883_preds(0) <= transition_879_symbol_out;
  place_883_succs(0) <= transition_880_symbol_out;
  place_883 : place
    generic map(marking => false)
    port map(
      preds => place_883_preds,
      succs => place_883_succs,
      token => place_883_token,
      clk   => clk,
      reset => reset);

  place_884_preds(0) <= transition_880_symbol_out;
  place_884_succs(0) <= transition_881_symbol_out;
  place_884 : place
    generic map(marking => false)
    port map(
      preds => place_884_preds,
      succs => place_884_succs,
      token => place_884_token,
      clk   => clk,
      reset => reset);

  place_890_preds(0) <= transition_886_symbol_out;
  place_890_succs(0) <= transition_887_symbol_out;
  place_890 : place
    generic map(marking => false)
    port map(
      preds => place_890_preds,
      succs => place_890_succs,
      token => place_890_token,
      clk   => clk,
      reset => reset);

  place_891_preds(0) <= transition_887_symbol_out;
  place_891_succs(0) <= transition_888_symbol_out;
  place_891 : place
    generic map(marking => false)
    port map(
      preds => place_891_preds,
      succs => place_891_succs,
      token => place_891_token,
      clk   => clk,
      reset => reset);

  place_892_preds(0) <= transition_888_symbol_out;
  place_892_succs(0) <= transition_889_symbol_out;
  place_892 : place
    generic map(marking => false)
    port map(
      preds => place_892_preds,
      succs => place_892_succs,
      token => place_892_token,
      clk   => clk,
      reset => reset);

  place_893_preds(0) <= transition_895_symbol_out;
  place_893_succs(0) <= transition_894_symbol_out;
  place_893 : place
    generic map(marking => false)
    port map(
      preds => place_893_preds,
      succs => place_893_succs,
      token => place_893_token,
      clk   => clk,
      reset => reset);

  place_897_preds(0) <= transition_899_symbol_out;
  place_897_succs(0) <= transition_898_symbol_out;
  place_897 : place
    generic map(marking => false)
    port map(
      preds => place_897_preds,
      succs => place_897_succs,
      token => place_897_token,
      clk   => clk,
      reset => reset);

  place_904_preds(0) <= transition_900_symbol_out;
  place_904_succs(0) <= transition_901_symbol_out;
  place_904 : place
    generic map(marking => false)
    port map(
      preds => place_904_preds,
      succs => place_904_succs,
      token => place_904_token,
      clk   => clk,
      reset => reset);

  place_905_preds(0) <= transition_901_symbol_out;
  place_905_succs(0) <= transition_902_symbol_out;
  place_905 : place
    generic map(marking => false)
    port map(
      preds => place_905_preds,
      succs => place_905_succs,
      token => place_905_token,
      clk   => clk,
      reset => reset);

  place_906_preds(0) <= transition_902_symbol_out;
  place_906_succs(0) <= transition_903_symbol_out;
  place_906 : place
    generic map(marking => false)
    port map(
      preds => place_906_preds,
      succs => place_906_succs,
      token => place_906_token,
      clk   => clk,
      reset => reset);

  place_911_preds(0) <= transition_907_symbol_out;
  place_911_succs(0) <= transition_908_symbol_out;
  place_911 : place
    generic map(marking => false)
    port map(
      preds => place_911_preds,
      succs => place_911_succs,
      token => place_911_token,
      clk   => clk,
      reset => reset);

  place_912_preds(0) <= transition_908_symbol_out;
  place_912_succs(0) <= transition_909_symbol_out;
  place_912 : place
    generic map(marking => false)
    port map(
      preds => place_912_preds,
      succs => place_912_succs,
      token => place_912_token,
      clk   => clk,
      reset => reset);

  place_913_preds(0) <= transition_909_symbol_out;
  place_913_succs(0) <= transition_910_symbol_out;
  place_913 : place
    generic map(marking => false)
    port map(
      preds => place_913_preds,
      succs => place_913_succs,
      token => place_913_token,
      clk   => clk,
      reset => reset);

  place_918_preds(0) <= transition_914_symbol_out;
  place_918_succs(0) <= transition_915_symbol_out;
  place_918 : place
    generic map(marking => false)
    port map(
      preds => place_918_preds,
      succs => place_918_succs,
      token => place_918_token,
      clk   => clk,
      reset => reset);

  place_919_preds(0) <= transition_915_symbol_out;
  place_919_succs(0) <= transition_916_symbol_out;
  place_919 : place
    generic map(marking => false)
    port map(
      preds => place_919_preds,
      succs => place_919_succs,
      token => place_919_token,
      clk   => clk,
      reset => reset);

  place_920_preds(0) <= transition_916_symbol_out;
  place_920_succs(0) <= transition_917_symbol_out;
  place_920 : place
    generic map(marking => false)
    port map(
      preds => place_920_preds,
      succs => place_920_succs,
      token => place_920_token,
      clk   => clk,
      reset => reset);

  place_926_preds(0) <= transition_922_symbol_out;
  place_926_succs(0) <= transition_923_symbol_out;
  place_926 : place
    generic map(marking => false)
    port map(
      preds => place_926_preds,
      succs => place_926_succs,
      token => place_926_token,
      clk   => clk,
      reset => reset);

  place_927_preds(0) <= transition_923_symbol_out;
  place_927_succs(0) <= transition_924_symbol_out;
  place_927 : place
    generic map(marking => false)
    port map(
      preds => place_927_preds,
      succs => place_927_succs,
      token => place_927_token,
      clk   => clk,
      reset => reset);

  place_928_preds(0) <= transition_924_symbol_out;
  place_928_succs(0) <= transition_925_symbol_out;
  place_928 : place
    generic map(marking => false)
    port map(
      preds => place_928_preds,
      succs => place_928_succs,
      token => place_928_token,
      clk   => clk,
      reset => reset);

  place_933_preds(0) <= transition_929_symbol_out;
  place_933_succs(0) <= transition_930_symbol_out;
  place_933 : place
    generic map(marking => false)
    port map(
      preds => place_933_preds,
      succs => place_933_succs,
      token => place_933_token,
      clk   => clk,
      reset => reset);

  place_934_preds(0) <= transition_930_symbol_out;
  place_934_succs(0) <= transition_931_symbol_out;
  place_934 : place
    generic map(marking => false)
    port map(
      preds => place_934_preds,
      succs => place_934_succs,
      token => place_934_token,
      clk   => clk,
      reset => reset);

  place_935_preds(0) <= transition_931_symbol_out;
  place_935_succs(0) <= transition_932_symbol_out;
  place_935 : place
    generic map(marking => false)
    port map(
      preds => place_935_preds,
      succs => place_935_succs,
      token => place_935_token,
      clk   => clk,
      reset => reset);

  place_941_preds(0) <= transition_937_symbol_out;
  place_941_succs(0) <= transition_938_symbol_out;
  place_941 : place
    generic map(marking => false)
    port map(
      preds => place_941_preds,
      succs => place_941_succs,
      token => place_941_token,
      clk   => clk,
      reset => reset);

  place_942_preds(0) <= transition_938_symbol_out;
  place_942_succs(0) <= transition_939_symbol_out;
  place_942 : place
    generic map(marking => false)
    port map(
      preds => place_942_preds,
      succs => place_942_succs,
      token => place_942_token,
      clk   => clk,
      reset => reset);

  place_943_preds(0) <= transition_939_symbol_out;
  place_943_succs(0) <= transition_940_symbol_out;
  place_943 : place
    generic map(marking => false)
    port map(
      preds => place_943_preds,
      succs => place_943_succs,
      token => place_943_token,
      clk   => clk,
      reset => reset);

  place_944_preds(0) <= transition_946_symbol_out;
  place_944_succs(0) <= transition_945_symbol_out;
  place_944 : place
    generic map(marking => false)
    port map(
      preds => place_944_preds,
      succs => place_944_succs,
      token => place_944_token,
      clk   => clk,
      reset => reset);

  place_948_preds(0) <= transition_950_symbol_out;
  place_948_succs(0) <= transition_949_symbol_out;
  place_948 : place
    generic map(marking => false)
    port map(
      preds => place_948_preds,
      succs => place_948_succs,
      token => place_948_token,
      clk   => clk,
      reset => reset);

  place_955_preds(0) <= transition_951_symbol_out;
  place_955_succs(0) <= transition_952_symbol_out;
  place_955 : place
    generic map(marking => false)
    port map(
      preds => place_955_preds,
      succs => place_955_succs,
      token => place_955_token,
      clk   => clk,
      reset => reset);

  place_956_preds(0) <= transition_952_symbol_out;
  place_956_succs(0) <= transition_953_symbol_out;
  place_956 : place
    generic map(marking => false)
    port map(
      preds => place_956_preds,
      succs => place_956_succs,
      token => place_956_token,
      clk   => clk,
      reset => reset);

  place_957_preds(0) <= transition_953_symbol_out;
  place_957_succs(0) <= transition_954_symbol_out;
  place_957 : place
    generic map(marking => false)
    port map(
      preds => place_957_preds,
      succs => place_957_succs,
      token => place_957_token,
      clk   => clk,
      reset => reset);

  place_963_preds(0) <= transition_959_symbol_out;
  place_963_succs(0) <= transition_960_symbol_out;
  place_963 : place
    generic map(marking => false)
    port map(
      preds => place_963_preds,
      succs => place_963_succs,
      token => place_963_token,
      clk   => clk,
      reset => reset);

  place_964_preds(0) <= transition_960_symbol_out;
  place_964_succs(0) <= transition_961_symbol_out;
  place_964 : place
    generic map(marking => false)
    port map(
      preds => place_964_preds,
      succs => place_964_succs,
      token => place_964_token,
      clk   => clk,
      reset => reset);

  place_965_preds(0) <= transition_961_symbol_out;
  place_965_succs(0) <= transition_962_symbol_out;
  place_965 : place
    generic map(marking => false)
    port map(
      preds => place_965_preds,
      succs => place_965_succs,
      token => place_965_token,
      clk   => clk,
      reset => reset);

  place_970_preds(0) <= transition_966_symbol_out;
  place_970_succs(0) <= transition_967_symbol_out;
  place_970 : place
    generic map(marking => false)
    port map(
      preds => place_970_preds,
      succs => place_970_succs,
      token => place_970_token,
      clk   => clk,
      reset => reset);

  place_971_preds(0) <= transition_967_symbol_out;
  place_971_succs(0) <= transition_968_symbol_out;
  place_971 : place
    generic map(marking => false)
    port map(
      preds => place_971_preds,
      succs => place_971_succs,
      token => place_971_token,
      clk   => clk,
      reset => reset);

  place_972_preds(0) <= transition_968_symbol_out;
  place_972_succs(0) <= transition_969_symbol_out;
  place_972 : place
    generic map(marking => false)
    port map(
      preds => place_972_preds,
      succs => place_972_succs,
      token => place_972_token,
      clk   => clk,
      reset => reset);

  place_977_preds(0) <= transition_973_symbol_out;
  place_977_succs(0) <= transition_974_symbol_out;
  place_977 : place
    generic map(marking => false)
    port map(
      preds => place_977_preds,
      succs => place_977_succs,
      token => place_977_token,
      clk   => clk,
      reset => reset);

  place_978_preds(0) <= transition_974_symbol_out;
  place_978_succs(0) <= transition_975_symbol_out;
  place_978 : place
    generic map(marking => false)
    port map(
      preds => place_978_preds,
      succs => place_978_succs,
      token => place_978_token,
      clk   => clk,
      reset => reset);

  place_979_preds(0) <= transition_975_symbol_out;
  place_979_succs(0) <= transition_976_symbol_out;
  place_979 : place
    generic map(marking => false)
    port map(
      preds => place_979_preds,
      succs => place_979_succs,
      token => place_979_token,
      clk   => clk,
      reset => reset);

  place_984_preds(0) <= transition_980_symbol_out;
  place_984_succs(0) <= transition_981_symbol_out;
  place_984 : place
    generic map(marking => false)
    port map(
      preds => place_984_preds,
      succs => place_984_succs,
      token => place_984_token,
      clk   => clk,
      reset => reset);

  place_985_preds(0) <= transition_981_symbol_out;
  place_985_succs(0) <= transition_982_symbol_out;
  place_985 : place
    generic map(marking => false)
    port map(
      preds => place_985_preds,
      succs => place_985_succs,
      token => place_985_token,
      clk   => clk,
      reset => reset);

  place_986_preds(0) <= transition_982_symbol_out;
  place_986_succs(0) <= transition_983_symbol_out;
  place_986 : place
    generic map(marking => false)
    port map(
      preds => place_986_preds,
      succs => place_986_succs,
      token => place_986_token,
      clk   => clk,
      reset => reset);

  place_992_preds(0) <= transition_988_symbol_out;
  place_992_succs(0) <= transition_989_symbol_out;
  place_992 : place
    generic map(marking => false)
    port map(
      preds => place_992_preds,
      succs => place_992_succs,
      token => place_992_token,
      clk   => clk,
      reset => reset);

  place_993_preds(0) <= transition_989_symbol_out;
  place_993_succs(0) <= transition_990_symbol_out;
  place_993 : place
    generic map(marking => false)
    port map(
      preds => place_993_preds,
      succs => place_993_succs,
      token => place_993_token,
      clk   => clk,
      reset => reset);

  place_994_preds(0) <= transition_990_symbol_out;
  place_994_succs(0) <= transition_991_symbol_out;
  place_994 : place
    generic map(marking => false)
    port map(
      preds => place_994_preds,
      succs => place_994_succs,
      token => place_994_token,
      clk   => clk,
      reset => reset);

  place_999_preds(0) <= transition_995_symbol_out;
  place_999_succs(0) <= transition_996_symbol_out;
  place_999 : place
    generic map(marking => false)
    port map(
      preds => place_999_preds,
      succs => place_999_succs,
      token => place_999_token,
      clk   => clk,
      reset => reset);

  place_1000_preds(0) <= transition_996_symbol_out;
  place_1000_succs(0) <= transition_997_symbol_out;
  place_1000 : place
    generic map(marking => false)
    port map(
      preds => place_1000_preds,
      succs => place_1000_succs,
      token => place_1000_token,
      clk   => clk,
      reset => reset);

  place_1001_preds(0) <= transition_997_symbol_out;
  place_1001_succs(0) <= transition_998_symbol_out;
  place_1001 : place
    generic map(marking => false)
    port map(
      preds => place_1001_preds,
      succs => place_1001_succs,
      token => place_1001_token,
      clk   => clk,
      reset => reset);

  place_1007_preds(0) <= transition_1003_symbol_out;
  place_1007_succs(0) <= transition_1004_symbol_out;
  place_1007 : place
    generic map(marking => false)
    port map(
      preds => place_1007_preds,
      succs => place_1007_succs,
      token => place_1007_token,
      clk   => clk,
      reset => reset);

  place_1008_preds(0) <= transition_1004_symbol_out;
  place_1008_succs(0) <= transition_1005_symbol_out;
  place_1008 : place
    generic map(marking => false)
    port map(
      preds => place_1008_preds,
      succs => place_1008_succs,
      token => place_1008_token,
      clk   => clk,
      reset => reset);

  place_1009_preds(0) <= transition_1005_symbol_out;
  place_1009_succs(0) <= transition_1006_symbol_out;
  place_1009 : place
    generic map(marking => false)
    port map(
      preds => place_1009_preds,
      succs => place_1009_succs,
      token => place_1009_token,
      clk   => clk,
      reset => reset);

  place_1010_preds(0) <= transition_1012_symbol_out;
  place_1010_succs(0) <= transition_1011_symbol_out;
  place_1010 : place
    generic map(marking => false)
    port map(
      preds => place_1010_preds,
      succs => place_1010_succs,
      token => place_1010_token,
      clk   => clk,
      reset => reset);

  place_1019_preds(0) <= transition_1015_symbol_out;
  place_1019_succs(0) <= transition_1016_symbol_out;
  place_1019 : place
    generic map(marking => false)
    port map(
      preds => place_1019_preds,
      succs => place_1019_succs,
      token => place_1019_token,
      clk   => clk,
      reset => reset);

  place_1020_preds(0) <= transition_1016_symbol_out;
  place_1020_succs(0) <= transition_1017_symbol_out;
  place_1020 : place
    generic map(marking => false)
    port map(
      preds => place_1020_preds,
      succs => place_1020_succs,
      token => place_1020_token,
      clk   => clk,
      reset => reset);

  place_1021_preds(0) <= transition_1017_symbol_out;
  place_1021_succs(0) <= transition_1018_symbol_out;
  place_1021 : place
    generic map(marking => false)
    port map(
      preds => place_1021_preds,
      succs => place_1021_succs,
      token => place_1021_token,
      clk   => clk,
      reset => reset);

  place_1026_preds(0) <= transition_1022_symbol_out;
  place_1026_succs(0) <= transition_1023_symbol_out;
  place_1026 : place
    generic map(marking => false)
    port map(
      preds => place_1026_preds,
      succs => place_1026_succs,
      token => place_1026_token,
      clk   => clk,
      reset => reset);

  place_1027_preds(0) <= transition_1023_symbol_out;
  place_1027_succs(0) <= transition_1024_symbol_out;
  place_1027 : place
    generic map(marking => false)
    port map(
      preds => place_1027_preds,
      succs => place_1027_succs,
      token => place_1027_token,
      clk   => clk,
      reset => reset);

  place_1028_preds(0) <= transition_1024_symbol_out;
  place_1028_succs(0) <= transition_1025_symbol_out;
  place_1028 : place
    generic map(marking => false)
    port map(
      preds => place_1028_preds,
      succs => place_1028_succs,
      token => place_1028_token,
      clk   => clk,
      reset => reset);

  place_1033_preds(0) <= transition_1029_symbol_out;
  place_1033_succs(0) <= transition_1030_symbol_out;
  place_1033 : place
    generic map(marking => false)
    port map(
      preds => place_1033_preds,
      succs => place_1033_succs,
      token => place_1033_token,
      clk   => clk,
      reset => reset);

  place_1034_preds(0) <= transition_1030_symbol_out;
  place_1034_succs(0) <= transition_1031_symbol_out;
  place_1034 : place
    generic map(marking => false)
    port map(
      preds => place_1034_preds,
      succs => place_1034_succs,
      token => place_1034_token,
      clk   => clk,
      reset => reset);

  place_1035_preds(0) <= transition_1031_symbol_out;
  place_1035_succs(0) <= transition_1032_symbol_out;
  place_1035 : place
    generic map(marking => false)
    port map(
      preds => place_1035_preds,
      succs => place_1035_succs,
      token => place_1035_token,
      clk   => clk,
      reset => reset);

  place_1041_preds(0) <= transition_1037_symbol_out;
  place_1041_succs(0) <= transition_1038_symbol_out;
  place_1041 : place
    generic map(marking => false)
    port map(
      preds => place_1041_preds,
      succs => place_1041_succs,
      token => place_1041_token,
      clk   => clk,
      reset => reset);

  place_1042_preds(0) <= transition_1038_symbol_out;
  place_1042_succs(0) <= transition_1039_symbol_out;
  place_1042 : place
    generic map(marking => false)
    port map(
      preds => place_1042_preds,
      succs => place_1042_succs,
      token => place_1042_token,
      clk   => clk,
      reset => reset);

  place_1043_preds(0) <= transition_1039_symbol_out;
  place_1043_succs(0) <= transition_1040_symbol_out;
  place_1043 : place
    generic map(marking => false)
    port map(
      preds => place_1043_preds,
      succs => place_1043_succs,
      token => place_1043_token,
      clk   => clk,
      reset => reset);

  place_1048_preds(0) <= transition_1044_symbol_out;
  place_1048_succs(0) <= transition_1045_symbol_out;
  place_1048 : place
    generic map(marking => false)
    port map(
      preds => place_1048_preds,
      succs => place_1048_succs,
      token => place_1048_token,
      clk   => clk,
      reset => reset);

  place_1049_preds(0) <= transition_1045_symbol_out;
  place_1049_succs(0) <= transition_1046_symbol_out;
  place_1049 : place
    generic map(marking => false)
    port map(
      preds => place_1049_preds,
      succs => place_1049_succs,
      token => place_1049_token,
      clk   => clk,
      reset => reset);

  place_1050_preds(0) <= transition_1046_symbol_out;
  place_1050_succs(0) <= transition_1047_symbol_out;
  place_1050 : place
    generic map(marking => false)
    port map(
      preds => place_1050_preds,
      succs => place_1050_succs,
      token => place_1050_token,
      clk   => clk,
      reset => reset);

  place_1056_preds(0) <= transition_1052_symbol_out;
  place_1056_succs(0) <= transition_1053_symbol_out;
  place_1056 : place
    generic map(marking => false)
    port map(
      preds => place_1056_preds,
      succs => place_1056_succs,
      token => place_1056_token,
      clk   => clk,
      reset => reset);

  place_1057_preds(0) <= transition_1053_symbol_out;
  place_1057_succs(0) <= transition_1054_symbol_out;
  place_1057 : place
    generic map(marking => false)
    port map(
      preds => place_1057_preds,
      succs => place_1057_succs,
      token => place_1057_token,
      clk   => clk,
      reset => reset);

  place_1058_preds(0) <= transition_1054_symbol_out;
  place_1058_succs(0) <= transition_1055_symbol_out;
  place_1058 : place
    generic map(marking => false)
    port map(
      preds => place_1058_preds,
      succs => place_1058_succs,
      token => place_1058_token,
      clk   => clk,
      reset => reset);

  place_1059_preds(0) <= transition_1061_symbol_out;
  place_1059_succs(0) <= transition_1060_symbol_out;
  place_1059 : place
    generic map(marking => false)
    port map(
      preds => place_1059_preds,
      succs => place_1059_succs,
      token => place_1059_token,
      clk   => clk,
      reset => reset);

  place_1063_preds(0) <= transition_1065_symbol_out;
  place_1063_succs(0) <= transition_1064_symbol_out;
  place_1063 : place
    generic map(marking => false)
    port map(
      preds => place_1063_preds,
      succs => place_1063_succs,
      token => place_1063_token,
      clk   => clk,
      reset => reset);

  place_1070_preds(0) <= transition_1066_symbol_out;
  place_1070_succs(0) <= transition_1067_symbol_out;
  place_1070 : place
    generic map(marking => false)
    port map(
      preds => place_1070_preds,
      succs => place_1070_succs,
      token => place_1070_token,
      clk   => clk,
      reset => reset);

  place_1071_preds(0) <= transition_1067_symbol_out;
  place_1071_succs(0) <= transition_1068_symbol_out;
  place_1071 : place
    generic map(marking => false)
    port map(
      preds => place_1071_preds,
      succs => place_1071_succs,
      token => place_1071_token,
      clk   => clk,
      reset => reset);

  place_1072_preds(0) <= transition_1068_symbol_out;
  place_1072_succs(0) <= transition_1069_symbol_out;
  place_1072 : place
    generic map(marking => false)
    port map(
      preds => place_1072_preds,
      succs => place_1072_succs,
      token => place_1072_token,
      clk   => clk,
      reset => reset);

  place_1077_preds(0) <= transition_1073_symbol_out;
  place_1077_succs(0) <= transition_1074_symbol_out;
  place_1077 : place
    generic map(marking => false)
    port map(
      preds => place_1077_preds,
      succs => place_1077_succs,
      token => place_1077_token,
      clk   => clk,
      reset => reset);

  place_1078_preds(0) <= transition_1074_symbol_out;
  place_1078_succs(0) <= transition_1075_symbol_out;
  place_1078 : place
    generic map(marking => false)
    port map(
      preds => place_1078_preds,
      succs => place_1078_succs,
      token => place_1078_token,
      clk   => clk,
      reset => reset);

  place_1079_preds(0) <= transition_1075_symbol_out;
  place_1079_succs(0) <= transition_1076_symbol_out;
  place_1079 : place
    generic map(marking => false)
    port map(
      preds => place_1079_preds,
      succs => place_1079_succs,
      token => place_1079_token,
      clk   => clk,
      reset => reset);

  place_1084_preds(0) <= transition_1080_symbol_out;
  place_1084_succs(0) <= transition_1081_symbol_out;
  place_1084 : place
    generic map(marking => false)
    port map(
      preds => place_1084_preds,
      succs => place_1084_succs,
      token => place_1084_token,
      clk   => clk,
      reset => reset);

  place_1085_preds(0) <= transition_1081_symbol_out;
  place_1085_succs(0) <= transition_1082_symbol_out;
  place_1085 : place
    generic map(marking => false)
    port map(
      preds => place_1085_preds,
      succs => place_1085_succs,
      token => place_1085_token,
      clk   => clk,
      reset => reset);

  place_1086_preds(0) <= transition_1082_symbol_out;
  place_1086_succs(0) <= transition_1083_symbol_out;
  place_1086 : place
    generic map(marking => false)
    port map(
      preds => place_1086_preds,
      succs => place_1086_succs,
      token => place_1086_token,
      clk   => clk,
      reset => reset);

  place_1092_preds(0) <= transition_1088_symbol_out;
  place_1092_succs(0) <= transition_1089_symbol_out;
  place_1092 : place
    generic map(marking => false)
    port map(
      preds => place_1092_preds,
      succs => place_1092_succs,
      token => place_1092_token,
      clk   => clk,
      reset => reset);

  place_1093_preds(0) <= transition_1089_symbol_out;
  place_1093_succs(0) <= transition_1090_symbol_out;
  place_1093 : place
    generic map(marking => false)
    port map(
      preds => place_1093_preds,
      succs => place_1093_succs,
      token => place_1093_token,
      clk   => clk,
      reset => reset);

  place_1094_preds(0) <= transition_1090_symbol_out;
  place_1094_succs(0) <= transition_1091_symbol_out;
  place_1094 : place
    generic map(marking => false)
    port map(
      preds => place_1094_preds,
      succs => place_1094_succs,
      token => place_1094_token,
      clk   => clk,
      reset => reset);

  place_1099_preds(0) <= transition_1095_symbol_out;
  place_1099_succs(0) <= transition_1096_symbol_out;
  place_1099 : place
    generic map(marking => false)
    port map(
      preds => place_1099_preds,
      succs => place_1099_succs,
      token => place_1099_token,
      clk   => clk,
      reset => reset);

  place_1100_preds(0) <= transition_1096_symbol_out;
  place_1100_succs(0) <= transition_1097_symbol_out;
  place_1100 : place
    generic map(marking => false)
    port map(
      preds => place_1100_preds,
      succs => place_1100_succs,
      token => place_1100_token,
      clk   => clk,
      reset => reset);

  place_1101_preds(0) <= transition_1097_symbol_out;
  place_1101_succs(0) <= transition_1098_symbol_out;
  place_1101 : place
    generic map(marking => false)
    port map(
      preds => place_1101_preds,
      succs => place_1101_succs,
      token => place_1101_token,
      clk   => clk,
      reset => reset);

  place_1107_preds(0) <= transition_1103_symbol_out;
  place_1107_succs(0) <= transition_1104_symbol_out;
  place_1107 : place
    generic map(marking => false)
    port map(
      preds => place_1107_preds,
      succs => place_1107_succs,
      token => place_1107_token,
      clk   => clk,
      reset => reset);

  place_1108_preds(0) <= transition_1104_symbol_out;
  place_1108_succs(0) <= transition_1105_symbol_out;
  place_1108 : place
    generic map(marking => false)
    port map(
      preds => place_1108_preds,
      succs => place_1108_succs,
      token => place_1108_token,
      clk   => clk,
      reset => reset);

  place_1109_preds(0) <= transition_1105_symbol_out;
  place_1109_succs(0) <= transition_1106_symbol_out;
  place_1109 : place
    generic map(marking => false)
    port map(
      preds => place_1109_preds,
      succs => place_1109_succs,
      token => place_1109_token,
      clk   => clk,
      reset => reset);

  place_1110_preds(0) <= transition_1112_symbol_out;
  place_1110_succs(0) <= transition_1111_symbol_out;
  place_1110 : place
    generic map(marking => false)
    port map(
      preds => place_1110_preds,
      succs => place_1110_succs,
      token => place_1110_token,
      clk   => clk,
      reset => reset);

  place_1114_preds(0) <= transition_1116_symbol_out;
  place_1114_succs(0) <= transition_1115_symbol_out;
  place_1114 : place
    generic map(marking => false)
    port map(
      preds => place_1114_preds,
      succs => place_1114_succs,
      token => place_1114_token,
      clk   => clk,
      reset => reset);

  place_1121_preds(0) <= transition_1117_symbol_out;
  place_1121_succs(0) <= transition_1118_symbol_out;
  place_1121 : place
    generic map(marking => false)
    port map(
      preds => place_1121_preds,
      succs => place_1121_succs,
      token => place_1121_token,
      clk   => clk,
      reset => reset);

  place_1122_preds(0) <= transition_1118_symbol_out;
  place_1122_succs(0) <= transition_1119_symbol_out;
  place_1122 : place
    generic map(marking => false)
    port map(
      preds => place_1122_preds,
      succs => place_1122_succs,
      token => place_1122_token,
      clk   => clk,
      reset => reset);

  place_1123_preds(0) <= transition_1119_symbol_out;
  place_1123_succs(0) <= transition_1120_symbol_out;
  place_1123 : place
    generic map(marking => false)
    port map(
      preds => place_1123_preds,
      succs => place_1123_succs,
      token => place_1123_token,
      clk   => clk,
      reset => reset);

  place_1129_preds(0) <= transition_1125_symbol_out;
  place_1129_succs(0) <= transition_1126_symbol_out;
  place_1129 : place
    generic map(marking => false)
    port map(
      preds => place_1129_preds,
      succs => place_1129_succs,
      token => place_1129_token,
      clk   => clk,
      reset => reset);

  place_1130_preds(0) <= transition_1126_symbol_out;
  place_1130_succs(0) <= transition_1127_symbol_out;
  place_1130 : place
    generic map(marking => false)
    port map(
      preds => place_1130_preds,
      succs => place_1130_succs,
      token => place_1130_token,
      clk   => clk,
      reset => reset);

  place_1131_preds(0) <= transition_1127_symbol_out;
  place_1131_succs(0) <= transition_1128_symbol_out;
  place_1131 : place
    generic map(marking => false)
    port map(
      preds => place_1131_preds,
      succs => place_1131_succs,
      token => place_1131_token,
      clk   => clk,
      reset => reset);

  place_1136_preds(0) <= transition_1132_symbol_out;
  place_1136_succs(0) <= transition_1133_symbol_out;
  place_1136 : place
    generic map(marking => false)
    port map(
      preds => place_1136_preds,
      succs => place_1136_succs,
      token => place_1136_token,
      clk   => clk,
      reset => reset);

  place_1137_preds(0) <= transition_1133_symbol_out;
  place_1137_succs(0) <= transition_1134_symbol_out;
  place_1137 : place
    generic map(marking => false)
    port map(
      preds => place_1137_preds,
      succs => place_1137_succs,
      token => place_1137_token,
      clk   => clk,
      reset => reset);

  place_1138_preds(0) <= transition_1134_symbol_out;
  place_1138_succs(0) <= transition_1135_symbol_out;
  place_1138 : place
    generic map(marking => false)
    port map(
      preds => place_1138_preds,
      succs => place_1138_succs,
      token => place_1138_token,
      clk   => clk,
      reset => reset);

  place_1143_preds(0) <= transition_1139_symbol_out;
  place_1143_succs(0) <= transition_1140_symbol_out;
  place_1143 : place
    generic map(marking => false)
    port map(
      preds => place_1143_preds,
      succs => place_1143_succs,
      token => place_1143_token,
      clk   => clk,
      reset => reset);

  place_1144_preds(0) <= transition_1140_symbol_out;
  place_1144_succs(0) <= transition_1141_symbol_out;
  place_1144 : place
    generic map(marking => false)
    port map(
      preds => place_1144_preds,
      succs => place_1144_succs,
      token => place_1144_token,
      clk   => clk,
      reset => reset);

  place_1145_preds(0) <= transition_1141_symbol_out;
  place_1145_succs(0) <= transition_1142_symbol_out;
  place_1145 : place
    generic map(marking => false)
    port map(
      preds => place_1145_preds,
      succs => place_1145_succs,
      token => place_1145_token,
      clk   => clk,
      reset => reset);

  place_1150_preds(0) <= transition_1146_symbol_out;
  place_1150_succs(0) <= transition_1147_symbol_out;
  place_1150 : place
    generic map(marking => false)
    port map(
      preds => place_1150_preds,
      succs => place_1150_succs,
      token => place_1150_token,
      clk   => clk,
      reset => reset);

  place_1151_preds(0) <= transition_1147_symbol_out;
  place_1151_succs(0) <= transition_1148_symbol_out;
  place_1151 : place
    generic map(marking => false)
    port map(
      preds => place_1151_preds,
      succs => place_1151_succs,
      token => place_1151_token,
      clk   => clk,
      reset => reset);

  place_1152_preds(0) <= transition_1148_symbol_out;
  place_1152_succs(0) <= transition_1149_symbol_out;
  place_1152 : place
    generic map(marking => false)
    port map(
      preds => place_1152_preds,
      succs => place_1152_succs,
      token => place_1152_token,
      clk   => clk,
      reset => reset);

  place_1158_preds(0) <= transition_1154_symbol_out;
  place_1158_succs(0) <= transition_1155_symbol_out;
  place_1158 : place
    generic map(marking => false)
    port map(
      preds => place_1158_preds,
      succs => place_1158_succs,
      token => place_1158_token,
      clk   => clk,
      reset => reset);

  place_1159_preds(0) <= transition_1155_symbol_out;
  place_1159_succs(0) <= transition_1156_symbol_out;
  place_1159 : place
    generic map(marking => false)
    port map(
      preds => place_1159_preds,
      succs => place_1159_succs,
      token => place_1159_token,
      clk   => clk,
      reset => reset);

  place_1160_preds(0) <= transition_1156_symbol_out;
  place_1160_succs(0) <= transition_1157_symbol_out;
  place_1160 : place
    generic map(marking => false)
    port map(
      preds => place_1160_preds,
      succs => place_1160_succs,
      token => place_1160_token,
      clk   => clk,
      reset => reset);

  place_1165_preds(0) <= transition_1161_symbol_out;
  place_1165_succs(0) <= transition_1162_symbol_out;
  place_1165 : place
    generic map(marking => false)
    port map(
      preds => place_1165_preds,
      succs => place_1165_succs,
      token => place_1165_token,
      clk   => clk,
      reset => reset);

  place_1166_preds(0) <= transition_1162_symbol_out;
  place_1166_succs(0) <= transition_1163_symbol_out;
  place_1166 : place
    generic map(marking => false)
    port map(
      preds => place_1166_preds,
      succs => place_1166_succs,
      token => place_1166_token,
      clk   => clk,
      reset => reset);

  place_1167_preds(0) <= transition_1163_symbol_out;
  place_1167_succs(0) <= transition_1164_symbol_out;
  place_1167 : place
    generic map(marking => false)
    port map(
      preds => place_1167_preds,
      succs => place_1167_succs,
      token => place_1167_token,
      clk   => clk,
      reset => reset);

  place_1173_preds(0) <= transition_1169_symbol_out;
  place_1173_succs(0) <= transition_1170_symbol_out;
  place_1173 : place
    generic map(marking => false)
    port map(
      preds => place_1173_preds,
      succs => place_1173_succs,
      token => place_1173_token,
      clk   => clk,
      reset => reset);

  place_1174_preds(0) <= transition_1170_symbol_out;
  place_1174_succs(0) <= transition_1171_symbol_out;
  place_1174 : place
    generic map(marking => false)
    port map(
      preds => place_1174_preds,
      succs => place_1174_succs,
      token => place_1174_token,
      clk   => clk,
      reset => reset);

  place_1175_preds(0) <= transition_1171_symbol_out;
  place_1175_succs(0) <= transition_1172_symbol_out;
  place_1175 : place
    generic map(marking => false)
    port map(
      preds => place_1175_preds,
      succs => place_1175_succs,
      token => place_1175_token,
      clk   => clk,
      reset => reset);

  place_1176_preds(0) <= transition_1178_symbol_out;
  place_1176_succs(0) <= transition_1177_symbol_out;
  place_1176 : place
    generic map(marking => false)
    port map(
      preds => place_1176_preds,
      succs => place_1176_succs,
      token => place_1176_token,
      clk   => clk,
      reset => reset);

  place_1184_preds(0) <= transition_1180_symbol_out;
  place_1184_succs(0) <= transition_1181_symbol_out;
  place_1184 : place
    generic map(marking => false)
    port map(
      preds => place_1184_preds,
      succs => place_1184_succs,
      token => place_1184_token,
      clk   => clk,
      reset => reset);

  place_1185_preds(0) <= transition_1181_symbol_out;
  place_1185_succs(0) <= transition_1182_symbol_out;
  place_1185 : place
    generic map(marking => false)
    port map(
      preds => place_1185_preds,
      succs => place_1185_succs,
      token => place_1185_token,
      clk   => clk,
      reset => reset);

  place_1186_preds(0) <= transition_1182_symbol_out;
  place_1186_succs(0) <= transition_1183_symbol_out;
  place_1186 : place
    generic map(marking => false)
    port map(
      preds => place_1186_preds,
      succs => place_1186_succs,
      token => place_1186_token,
      clk   => clk,
      reset => reset);

  place_1192_preds(0) <= transition_1188_symbol_out;
  place_1192_succs(0) <= transition_1189_symbol_out;
  place_1192 : place
    generic map(marking => false)
    port map(
      preds => place_1192_preds,
      succs => place_1192_succs,
      token => place_1192_token,
      clk   => clk,
      reset => reset);

  place_1193_preds(0) <= transition_1189_symbol_out;
  place_1193_succs(0) <= transition_1190_symbol_out;
  place_1193 : place
    generic map(marking => false)
    port map(
      preds => place_1193_preds,
      succs => place_1193_succs,
      token => place_1193_token,
      clk   => clk,
      reset => reset);

  place_1194_preds(0) <= transition_1190_symbol_out;
  place_1194_succs(0) <= transition_1191_symbol_out;
  place_1194 : place
    generic map(marking => false)
    port map(
      preds => place_1194_preds,
      succs => place_1194_succs,
      token => place_1194_token,
      clk   => clk,
      reset => reset);

  place_1200_preds(0) <= transition_1196_symbol_out;
  place_1200_succs(0) <= transition_1197_symbol_out;
  place_1200 : place
    generic map(marking => false)
    port map(
      preds => place_1200_preds,
      succs => place_1200_succs,
      token => place_1200_token,
      clk   => clk,
      reset => reset);

  place_1201_preds(0) <= transition_1197_symbol_out;
  place_1201_succs(0) <= transition_1198_symbol_out;
  place_1201 : place
    generic map(marking => false)
    port map(
      preds => place_1201_preds,
      succs => place_1201_succs,
      token => place_1201_token,
      clk   => clk,
      reset => reset);

  place_1202_preds(0) <= transition_1198_symbol_out;
  place_1202_succs(0) <= transition_1199_symbol_out;
  place_1202 : place
    generic map(marking => false)
    port map(
      preds => place_1202_preds,
      succs => place_1202_succs,
      token => place_1202_token,
      clk   => clk,
      reset => reset);

  place_1203_preds(0) <= transition_1205_symbol_out;
  place_1203_succs(0) <= transition_1204_symbol_out;
  place_1203 : place
    generic map(marking => false)
    port map(
      preds => place_1203_preds,
      succs => place_1203_succs,
      token => place_1203_token,
      clk   => clk,
      reset => reset);

  place_1206_preds(0) <= transition_1_symbol_out;
  place_1206_succs(0) <= transition_7_symbol_out;
  place_1206 : place
    generic map(marking => false)
    port map(
      preds => place_1206_preds,
      succs => place_1206_succs,
      token => place_1206_token,
      clk   => clk,
      reset => reset);

  place_1207_preds(0) <= transition_157_symbol_out;
  place_1207_succs(0) <= transition_150_symbol_out;
  place_1207 : place
    generic map(marking => false)
    port map(
      preds => place_1207_preds,
      succs => place_1207_succs,
      token => place_1207_token,
      clk   => clk,
      reset => reset);

  place_1208_preds(0) <= transition_153_symbol_out;
  place_1208_succs(0) <= transition_158_symbol_out;
  place_1208 : place
    generic map(marking => false)
    port map(
      preds => place_1208_preds,
      succs => place_1208_succs,
      token => place_1208_token,
      clk   => clk,
      reset => reset);

  place_1209_preds(0) <= transition_161_symbol_out;
  place_1209_succs(0) <= transition_168_symbol_out;
  place_1209 : place
    generic map(marking => false)
    port map(
      preds => place_1209_preds,
      succs => place_1209_succs,
      token => place_1209_token,
      clk   => clk,
      reset => reset);

  place_1210_preds(0) <= transition_168_symbol_out;
  place_1210_succs(0) <= transition_167_symbol_out;
  place_1210 : place
    generic map(marking => false)
    port map(
      preds => place_1210_preds,
      succs => place_1210_succs,
      token => place_1210_token,
      clk   => clk,
      reset => reset);

  place_1211_preds(0) <= transition_166_symbol_out;
  place_1211_succs(0) <= transition_169_symbol_out;
  place_1211 : place
    generic map(marking => false)
    port map(
      preds => place_1211_preds,
      succs => place_1211_succs,
      token => place_1211_token,
      clk   => clk,
      reset => reset);

  place_1212_preds(0) <= transition_120_symbol_out;
  place_1212_succs(0) <= transition_168_symbol_out;
  place_1212 : place
    generic map(marking => false)
    port map(
      preds => place_1212_preds,
      succs => place_1212_succs,
      token => place_1212_token,
      clk   => clk,
      reset => reset);

  place_1213_preds(0) <= transition_173_symbol_out;
  place_1213_succs(0) <= transition_191_symbol_out;
  place_1213 : place
    generic map(marking => false)
    port map(
      preds => place_1213_preds,
      succs => place_1213_succs,
      token => place_1213_token,
      clk   => clk,
      reset => reset);

  place_1214_preds(0) <= transition_3_symbol_out;
  place_1214_succs(0) <= transition_170_symbol_out;
  place_1214 : place
    generic map(marking => false)
    port map(
      preds => place_1214_preds,
      succs => place_1214_succs,
      token => place_1214_token,
      clk   => clk,
      reset => reset);

  place_1215_preds(0) <= transition_180_symbol_out;
  place_1215_succs(0) <= transition_191_symbol_out;
  place_1215 : place
    generic map(marking => false)
    port map(
      preds => place_1215_preds,
      succs => place_1215_succs,
      token => place_1215_token,
      clk   => clk,
      reset => reset);

  place_1216_preds(0) <= transition_3_symbol_out;
  place_1216_succs(0) <= transition_177_symbol_out;
  place_1216 : place
    generic map(marking => false)
    port map(
      preds => place_1216_preds,
      succs => place_1216_succs,
      token => place_1216_token,
      clk   => clk,
      reset => reset);

  place_1217_preds(0) <= transition_191_symbol_out;
  place_1217_succs(0) <= transition_184_symbol_out;
  place_1217 : place
    generic map(marking => false)
    port map(
      preds => place_1217_preds,
      succs => place_1217_succs,
      token => place_1217_token,
      clk   => clk,
      reset => reset);

  place_1218_preds(0) <= transition_187_symbol_out;
  place_1218_succs(0) <= transition_206_symbol_out;
  place_1218 : place
    generic map(marking => false)
    port map(
      preds => place_1218_preds,
      succs => place_1218_succs,
      token => place_1218_token,
      clk   => clk,
      reset => reset);

  place_1219_preds(0) <= transition_195_symbol_out;
  place_1219_succs(0) <= transition_206_symbol_out;
  place_1219 : place
    generic map(marking => false)
    port map(
      preds => place_1219_preds,
      succs => place_1219_succs,
      token => place_1219_token,
      clk   => clk,
      reset => reset);

  place_1220_preds(0) <= transition_3_symbol_out;
  place_1220_succs(0) <= transition_15_symbol_out;
  place_1220 : place
    generic map(marking => false)
    port map(
      preds => place_1220_preds,
      succs => place_1220_succs,
      token => place_1220_token,
      clk   => clk,
      reset => reset);

  place_1221_preds(0) <= transition_3_symbol_out;
  place_1221_succs(0) <= transition_192_symbol_out;
  place_1221 : place
    generic map(marking => false)
    port map(
      preds => place_1221_preds,
      succs => place_1221_succs,
      token => place_1221_token,
      clk   => clk,
      reset => reset);

  place_1222_preds(0) <= transition_206_symbol_out;
  place_1222_succs(0) <= transition_199_symbol_out;
  place_1222 : place
    generic map(marking => false)
    port map(
      preds => place_1222_preds,
      succs => place_1222_succs,
      token => place_1222_token,
      clk   => clk,
      reset => reset);

  place_1223_preds(0) <= transition_202_symbol_out;
  place_1223_succs(0) <= transition_207_symbol_out;
  place_1223 : place
    generic map(marking => false)
    port map(
      preds => place_1223_preds,
      succs => place_1223_succs,
      token => place_1223_token,
      clk   => clk,
      reset => reset);

  place_1224_preds(0) <= transition_210_symbol_out;
  place_1224_succs(0) <= transition_217_symbol_out;
  place_1224 : place
    generic map(marking => false)
    port map(
      preds => place_1224_preds,
      succs => place_1224_succs,
      token => place_1224_token,
      clk   => clk,
      reset => reset);

  place_1225_preds(0) <= transition_29_symbol_out;
  place_1225_succs(0) <= transition_22_symbol_out;
  place_1225 : place
    generic map(marking => false)
    port map(
      preds => place_1225_preds,
      succs => place_1225_succs,
      token => place_1225_token,
      clk   => clk,
      reset => reset);

  place_1226_preds(0) <= transition_217_symbol_out;
  place_1226_succs(0) <= transition_216_symbol_out;
  place_1226 : place
    generic map(marking => false)
    port map(
      preds => place_1226_preds,
      succs => place_1226_succs,
      token => place_1226_token,
      clk   => clk,
      reset => reset);

  place_1227_preds(0) <= transition_215_symbol_out;
  place_1227_succs(0) <= transition_220_symbol_out;
  place_1227 : place
    generic map(marking => false)
    port map(
      preds => place_1227_preds,
      succs => place_1227_succs,
      token => place_1227_token,
      clk   => clk,
      reset => reset);

  place_1228_preds(0) <= transition_219_symbol_out;
  place_1228_succs(0) <= transition_221_symbol_out;
  place_1228 : place
    generic map(marking => false)
    port map(
      preds => place_1228_preds,
      succs => place_1228_succs,
      token => place_1228_token,
      clk   => clk,
      reset => reset);

  place_1229_preds(0) <= transition_169_symbol_out;
  place_1229_succs(0) <= transition_217_symbol_out;
  place_1229 : place
    generic map(marking => false)
    port map(
      preds => place_1229_preds,
      succs => place_1229_succs,
      token => place_1229_token,
      clk   => clk,
      reset => reset);

  place_1230_preds(0) <= transition_225_symbol_out;
  place_1230_succs(0) <= transition_243_symbol_out;
  place_1230 : place
    generic map(marking => false)
    port map(
      preds => place_1230_preds,
      succs => place_1230_succs,
      token => place_1230_token,
      clk   => clk,
      reset => reset);

  place_1231_preds(0) <= transition_25_symbol_out;
  place_1231_succs(0) <= transition_44_symbol_out;
  place_1231 : place
    generic map(marking => false)
    port map(
      preds => place_1231_preds,
      succs => place_1231_succs,
      token => place_1231_token,
      clk   => clk,
      reset => reset);

  place_1232_preds(0) <= transition_3_symbol_out;
  place_1232_succs(0) <= transition_222_symbol_out;
  place_1232 : place
    generic map(marking => false)
    port map(
      preds => place_1232_preds,
      succs => place_1232_succs,
      token => place_1232_token,
      clk   => clk,
      reset => reset);

  place_1233_preds(0) <= transition_232_symbol_out;
  place_1233_succs(0) <= transition_243_symbol_out;
  place_1233 : place
    generic map(marking => false)
    port map(
      preds => place_1233_preds,
      succs => place_1233_succs,
      token => place_1233_token,
      clk   => clk,
      reset => reset);

  place_1234_preds(0) <= transition_3_symbol_out;
  place_1234_succs(0) <= transition_229_symbol_out;
  place_1234 : place
    generic map(marking => false)
    port map(
      preds => place_1234_preds,
      succs => place_1234_succs,
      token => place_1234_token,
      clk   => clk,
      reset => reset);

  place_1235_preds(0) <= transition_243_symbol_out;
  place_1235_succs(0) <= transition_236_symbol_out;
  place_1235 : place
    generic map(marking => false)
    port map(
      preds => place_1235_preds,
      succs => place_1235_succs,
      token => place_1235_token,
      clk   => clk,
      reset => reset);

  place_1236_preds(0) <= transition_239_symbol_out;
  place_1236_succs(0) <= transition_258_symbol_out;
  place_1236 : place
    generic map(marking => false)
    port map(
      preds => place_1236_preds,
      succs => place_1236_succs,
      token => place_1236_token,
      clk   => clk,
      reset => reset);

  place_1237_preds(0) <= transition_247_symbol_out;
  place_1237_succs(0) <= transition_258_symbol_out;
  place_1237 : place
    generic map(marking => false)
    port map(
      preds => place_1237_preds,
      succs => place_1237_succs,
      token => place_1237_token,
      clk   => clk,
      reset => reset);

  place_1238_preds(0) <= transition_3_symbol_out;
  place_1238_succs(0) <= transition_244_symbol_out;
  place_1238 : place
    generic map(marking => false)
    port map(
      preds => place_1238_preds,
      succs => place_1238_succs,
      token => place_1238_token,
      clk   => clk,
      reset => reset);

  place_1239_preds(0) <= transition_258_symbol_out;
  place_1239_succs(0) <= transition_251_symbol_out;
  place_1239 : place
    generic map(marking => false)
    port map(
      preds => place_1239_preds,
      succs => place_1239_succs,
      token => place_1239_token,
      clk   => clk,
      reset => reset);

  place_1240_preds(0) <= transition_254_symbol_out;
  place_1240_succs(0) <= transition_259_symbol_out;
  place_1240 : place
    generic map(marking => false)
    port map(
      preds => place_1240_preds,
      succs => place_1240_succs,
      token => place_1240_token,
      clk   => clk,
      reset => reset);

  place_1241_preds(0) <= transition_262_symbol_out;
  place_1241_succs(0) <= transition_269_symbol_out;
  place_1241 : place
    generic map(marking => false)
    port map(
      preds => place_1241_preds,
      succs => place_1241_succs,
      token => place_1241_token,
      clk   => clk,
      reset => reset);

  place_1242_preds(0) <= transition_269_symbol_out;
  place_1242_succs(0) <= transition_268_symbol_out;
  place_1242 : place
    generic map(marking => false)
    port map(
      preds => place_1242_preds,
      succs => place_1242_succs,
      token => place_1242_token,
      clk   => clk,
      reset => reset);

  place_1243_preds(0) <= transition_267_symbol_out;
  place_1243_succs(0) <= transition_272_symbol_out;
  place_1243 : place
    generic map(marking => false)
    port map(
      preds => place_1243_preds,
      succs => place_1243_succs,
      token => place_1243_token,
      clk   => clk,
      reset => reset);

  place_1244_preds(0) <= transition_271_symbol_out;
  place_1244_succs(0) <= transition_273_symbol_out;
  place_1244 : place
    generic map(marking => false)
    port map(
      preds => place_1244_preds,
      succs => place_1244_succs,
      token => place_1244_token,
      clk   => clk,
      reset => reset);

  place_1245_preds(0) <= transition_169_symbol_out;
  place_1245_succs(0) <= transition_269_symbol_out;
  place_1245 : place
    generic map(marking => false)
    port map(
      preds => place_1245_preds,
      succs => place_1245_succs,
      token => place_1245_token,
      clk   => clk,
      reset => reset);

  place_1246_preds(0) <= transition_281_symbol_out;
  place_1246_succs(0) <= transition_274_symbol_out;
  place_1246 : place
    generic map(marking => false)
    port map(
      preds => place_1246_preds,
      succs => place_1246_succs,
      token => place_1246_token,
      clk   => clk,
      reset => reset);

  place_1247_preds(0) <= transition_277_symbol_out;
  place_1247_succs(0) <= transition_282_symbol_out;
  place_1247 : place
    generic map(marking => false)
    port map(
      preds => place_1247_preds,
      succs => place_1247_succs,
      token => place_1247_token,
      clk   => clk,
      reset => reset);

  place_1248_preds(0) <= transition_221_symbol_out;
  place_1248_succs(0) <= transition_281_symbol_out;
  place_1248 : place
    generic map(marking => false)
    port map(
      preds => place_1248_preds,
      succs => place_1248_succs,
      token => place_1248_token,
      clk   => clk,
      reset => reset);

  place_1249_preds(0) <= transition_273_symbol_out;
  place_1249_succs(0) <= transition_281_symbol_out;
  place_1249 : place
    generic map(marking => false)
    port map(
      preds => place_1249_preds,
      succs => place_1249_succs,
      token => place_1249_token,
      clk   => clk,
      reset => reset);

  place_1250_preds(0) <= transition_286_symbol_out;
  place_1250_succs(0) <= transition_304_symbol_out;
  place_1250 : place
    generic map(marking => false)
    port map(
      preds => place_1250_preds,
      succs => place_1250_succs,
      token => place_1250_token,
      clk   => clk,
      reset => reset);

  place_1251_preds(0) <= transition_3_symbol_out;
  place_1251_succs(0) <= transition_283_symbol_out;
  place_1251 : place
    generic map(marking => false)
    port map(
      preds => place_1251_preds,
      succs => place_1251_succs,
      token => place_1251_token,
      clk   => clk,
      reset => reset);

  place_1252_preds(0) <= transition_293_symbol_out;
  place_1252_succs(0) <= transition_304_symbol_out;
  place_1252 : place
    generic map(marking => false)
    port map(
      preds => place_1252_preds,
      succs => place_1252_succs,
      token => place_1252_token,
      clk   => clk,
      reset => reset);

  place_1253_preds(0) <= transition_3_symbol_out;
  place_1253_succs(0) <= transition_290_symbol_out;
  place_1253 : place
    generic map(marking => false)
    port map(
      preds => place_1253_preds,
      succs => place_1253_succs,
      token => place_1253_token,
      clk   => clk,
      reset => reset);

  place_1254_preds(0) <= transition_304_symbol_out;
  place_1254_succs(0) <= transition_297_symbol_out;
  place_1254 : place
    generic map(marking => false)
    port map(
      preds => place_1254_preds,
      succs => place_1254_succs,
      token => place_1254_token,
      clk   => clk,
      reset => reset);

  place_1255_preds(0) <= transition_300_symbol_out;
  place_1255_succs(0) <= transition_319_symbol_out;
  place_1255 : place
    generic map(marking => false)
    port map(
      preds => place_1255_preds,
      succs => place_1255_succs,
      token => place_1255_token,
      clk   => clk,
      reset => reset);

  place_1256_preds(0) <= transition_6_symbol_out;
  place_1256_succs(0) <= transition_3_symbol_out;
  place_1256 : place
    generic map(marking => false)
    port map(
      preds => place_1256_preds,
      succs => place_1256_succs,
      token => place_1256_token,
      clk   => clk,
      reset => reset);

  place_1257_preds(0) <= transition_33_symbol_out;
  place_1257_succs(0) <= transition_44_symbol_out;
  place_1257 : place
    generic map(marking => false)
    port map(
      preds => place_1257_preds,
      succs => place_1257_succs,
      token => place_1257_token,
      clk   => clk,
      reset => reset);

  place_1258_preds(0) <= transition_308_symbol_out;
  place_1258_succs(0) <= transition_319_symbol_out;
  place_1258 : place
    generic map(marking => false)
    port map(
      preds => place_1258_preds,
      succs => place_1258_succs,
      token => place_1258_token,
      clk   => clk,
      reset => reset);

  place_1259_preds(0) <= transition_3_symbol_out;
  place_1259_succs(0) <= transition_305_symbol_out;
  place_1259 : place
    generic map(marking => false)
    port map(
      preds => place_1259_preds,
      succs => place_1259_succs,
      token => place_1259_token,
      clk   => clk,
      reset => reset);

  place_1260_preds(0) <= transition_319_symbol_out;
  place_1260_succs(0) <= transition_312_symbol_out;
  place_1260 : place
    generic map(marking => false)
    port map(
      preds => place_1260_preds,
      succs => place_1260_succs,
      token => place_1260_token,
      clk   => clk,
      reset => reset);

  place_1261_preds(0) <= transition_315_symbol_out;
  place_1261_succs(0) <= transition_320_symbol_out;
  place_1261 : place
    generic map(marking => false)
    port map(
      preds => place_1261_preds,
      succs => place_1261_succs,
      token => place_1261_token,
      clk   => clk,
      reset => reset);

  place_1262_preds(0) <= transition_323_symbol_out;
  place_1262_succs(0) <= transition_330_symbol_out;
  place_1262 : place
    generic map(marking => false)
    port map(
      preds => place_1262_preds,
      succs => place_1262_succs,
      token => place_1262_token,
      clk   => clk,
      reset => reset);

  place_1263_preds(0) <= transition_330_symbol_out;
  place_1263_succs(0) <= transition_329_symbol_out;
  place_1263 : place
    generic map(marking => false)
    port map(
      preds => place_1263_preds,
      succs => place_1263_succs,
      token => place_1263_token,
      clk   => clk,
      reset => reset);

  place_1264_preds(0) <= transition_328_symbol_out;
  place_1264_succs(0) <= transition_331_symbol_out;
  place_1264 : place
    generic map(marking => false)
    port map(
      preds => place_1264_preds,
      succs => place_1264_succs,
      token => place_1264_token,
      clk   => clk,
      reset => reset);

  place_1265_preds(0) <= transition_282_symbol_out;
  place_1265_succs(0) <= transition_330_symbol_out;
  place_1265 : place
    generic map(marking => false)
    port map(
      preds => place_1265_preds,
      succs => place_1265_succs,
      token => place_1265_token,
      clk   => clk,
      reset => reset);

  place_1266_preds(0) <= transition_335_symbol_out;
  place_1266_succs(0) <= transition_353_symbol_out;
  place_1266 : place
    generic map(marking => false)
    port map(
      preds => place_1266_preds,
      succs => place_1266_succs,
      token => place_1266_token,
      clk   => clk,
      reset => reset);

  place_1267_preds(0) <= transition_3_symbol_out;
  place_1267_succs(0) <= transition_332_symbol_out;
  place_1267 : place
    generic map(marking => false)
    port map(
      preds => place_1267_preds,
      succs => place_1267_succs,
      token => place_1267_token,
      clk   => clk,
      reset => reset);

  place_1268_preds(0) <= transition_342_symbol_out;
  place_1268_succs(0) <= transition_353_symbol_out;
  place_1268 : place
    generic map(marking => false)
    port map(
      preds => place_1268_preds,
      succs => place_1268_succs,
      token => place_1268_token,
      clk   => clk,
      reset => reset);

  place_1269_preds(0) <= transition_3_symbol_out;
  place_1269_succs(0) <= transition_339_symbol_out;
  place_1269 : place
    generic map(marking => false)
    port map(
      preds => place_1269_preds,
      succs => place_1269_succs,
      token => place_1269_token,
      clk   => clk,
      reset => reset);

  place_1270_preds(0) <= transition_353_symbol_out;
  place_1270_succs(0) <= transition_346_symbol_out;
  place_1270 : place
    generic map(marking => false)
    port map(
      preds => place_1270_preds,
      succs => place_1270_succs,
      token => place_1270_token,
      clk   => clk,
      reset => reset);

  place_1271_preds(0) <= transition_349_symbol_out;
  place_1271_succs(0) <= transition_368_symbol_out;
  place_1271 : place
    generic map(marking => false)
    port map(
      preds => place_1271_preds,
      succs => place_1271_succs,
      token => place_1271_token,
      clk   => clk,
      reset => reset);

  place_1272_preds(0) <= transition_3_symbol_out;
  place_1272_succs(0) <= transition_30_symbol_out;
  place_1272 : place
    generic map(marking => false)
    port map(
      preds => place_1272_preds,
      succs => place_1272_succs,
      token => place_1272_token,
      clk   => clk,
      reset => reset);

  place_1273_preds(0) <= transition_357_symbol_out;
  place_1273_succs(0) <= transition_368_symbol_out;
  place_1273 : place
    generic map(marking => false)
    port map(
      preds => place_1273_preds,
      succs => place_1273_succs,
      token => place_1273_token,
      clk   => clk,
      reset => reset);

  place_1274_preds(0) <= transition_3_symbol_out;
  place_1274_succs(0) <= transition_354_symbol_out;
  place_1274 : place
    generic map(marking => false)
    port map(
      preds => place_1274_preds,
      succs => place_1274_succs,
      token => place_1274_token,
      clk   => clk,
      reset => reset);

  place_1275_preds(0) <= transition_368_symbol_out;
  place_1275_succs(0) <= transition_361_symbol_out;
  place_1275 : place
    generic map(marking => false)
    port map(
      preds => place_1275_preds,
      succs => place_1275_succs,
      token => place_1275_token,
      clk   => clk,
      reset => reset);

  place_1276_preds(0) <= transition_364_symbol_out;
  place_1276_succs(0) <= transition_369_symbol_out;
  place_1276 : place
    generic map(marking => false)
    port map(
      preds => place_1276_preds,
      succs => place_1276_succs,
      token => place_1276_token,
      clk   => clk,
      reset => reset);

  place_1277_preds(0) <= transition_44_symbol_out;
  place_1277_succs(0) <= transition_37_symbol_out;
  place_1277 : place
    generic map(marking => false)
    port map(
      preds => place_1277_preds,
      succs => place_1277_succs,
      token => place_1277_token,
      clk   => clk,
      reset => reset);

  place_1278_preds(0) <= transition_372_symbol_out;
  place_1278_succs(0) <= transition_379_symbol_out;
  place_1278 : place
    generic map(marking => false)
    port map(
      preds => place_1278_preds,
      succs => place_1278_succs,
      token => place_1278_token,
      clk   => clk,
      reset => reset);

  place_1279_preds(0) <= transition_379_symbol_out;
  place_1279_succs(0) <= transition_378_symbol_out;
  place_1279 : place
    generic map(marking => false)
    port map(
      preds => place_1279_preds,
      succs => place_1279_succs,
      token => place_1279_token,
      clk   => clk,
      reset => reset);

  place_1280_preds(0) <= transition_377_symbol_out;
  place_1280_succs(0) <= transition_382_symbol_out;
  place_1280 : place
    generic map(marking => false)
    port map(
      preds => place_1280_preds,
      succs => place_1280_succs,
      token => place_1280_token,
      clk   => clk,
      reset => reset);

  place_1281_preds(0) <= transition_381_symbol_out;
  place_1281_succs(0) <= transition_383_symbol_out;
  place_1281 : place
    generic map(marking => false)
    port map(
      preds => place_1281_preds,
      succs => place_1281_succs,
      token => place_1281_token,
      clk   => clk,
      reset => reset);

  place_1282_preds(0) <= transition_40_symbol_out;
  place_1282_succs(0) <= transition_45_symbol_out;
  place_1282 : place
    generic map(marking => false)
    port map(
      preds => place_1282_preds,
      succs => place_1282_succs,
      token => place_1282_token,
      clk   => clk,
      reset => reset);

  place_1283_preds(0) <= transition_331_symbol_out;
  place_1283_succs(0) <= transition_379_symbol_out;
  place_1283 : place
    generic map(marking => false)
    port map(
      preds => place_1283_preds,
      succs => place_1283_succs,
      token => place_1283_token,
      clk   => clk,
      reset => reset);

  place_1284_preds(0) <= transition_387_symbol_out;
  place_1284_succs(0) <= transition_405_symbol_out;
  place_1284 : place
    generic map(marking => false)
    port map(
      preds => place_1284_preds,
      succs => place_1284_succs,
      token => place_1284_token,
      clk   => clk,
      reset => reset);

  place_1285_preds(0) <= transition_3_symbol_out;
  place_1285_succs(0) <= transition_384_symbol_out;
  place_1285 : place
    generic map(marking => false)
    port map(
      preds => place_1285_preds,
      succs => place_1285_succs,
      token => place_1285_token,
      clk   => clk,
      reset => reset);

  place_1286_preds(0) <= transition_394_symbol_out;
  place_1286_succs(0) <= transition_405_symbol_out;
  place_1286 : place
    generic map(marking => false)
    port map(
      preds => place_1286_preds,
      succs => place_1286_succs,
      token => place_1286_token,
      clk   => clk,
      reset => reset);

  place_1287_preds(0) <= transition_3_symbol_out;
  place_1287_succs(0) <= transition_391_symbol_out;
  place_1287 : place
    generic map(marking => false)
    port map(
      preds => place_1287_preds,
      succs => place_1287_succs,
      token => place_1287_token,
      clk   => clk,
      reset => reset);

  place_1288_preds(0) <= transition_405_symbol_out;
  place_1288_succs(0) <= transition_398_symbol_out;
  place_1288 : place
    generic map(marking => false)
    port map(
      preds => place_1288_preds,
      succs => place_1288_succs,
      token => place_1288_token,
      clk   => clk,
      reset => reset);

  place_1289_preds(0) <= transition_401_symbol_out;
  place_1289_succs(0) <= transition_420_symbol_out;
  place_1289 : place
    generic map(marking => false)
    port map(
      preds => place_1289_preds,
      succs => place_1289_succs,
      token => place_1289_token,
      clk   => clk,
      reset => reset);

  place_1290_preds(0) <= transition_409_symbol_out;
  place_1290_succs(0) <= transition_420_symbol_out;
  place_1290 : place
    generic map(marking => false)
    port map(
      preds => place_1290_preds,
      succs => place_1290_succs,
      token => place_1290_token,
      clk   => clk,
      reset => reset);

  place_1291_preds(0) <= transition_3_symbol_out;
  place_1291_succs(0) <= transition_406_symbol_out;
  place_1291 : place
    generic map(marking => false)
    port map(
      preds => place_1291_preds,
      succs => place_1291_succs,
      token => place_1291_token,
      clk   => clk,
      reset => reset);

  place_1292_preds(0) <= transition_420_symbol_out;
  place_1292_succs(0) <= transition_413_symbol_out;
  place_1292 : place
    generic map(marking => false)
    port map(
      preds => place_1292_preds,
      succs => place_1292_succs,
      token => place_1292_token,
      clk   => clk,
      reset => reset);

  place_1293_preds(0) <= transition_416_symbol_out;
  place_1293_succs(0) <= transition_421_symbol_out;
  place_1293 : place
    generic map(marking => false)
    port map(
      preds => place_1293_preds,
      succs => place_1293_succs,
      token => place_1293_token,
      clk   => clk,
      reset => reset);

  place_1294_preds(0) <= transition_424_symbol_out;
  place_1294_succs(0) <= transition_431_symbol_out;
  place_1294 : place
    generic map(marking => false)
    port map(
      preds => place_1294_preds,
      succs => place_1294_succs,
      token => place_1294_token,
      clk   => clk,
      reset => reset);

  place_1295_preds(0) <= transition_431_symbol_out;
  place_1295_succs(0) <= transition_430_symbol_out;
  place_1295 : place
    generic map(marking => false)
    port map(
      preds => place_1295_preds,
      succs => place_1295_succs,
      token => place_1295_token,
      clk   => clk,
      reset => reset);

  place_1296_preds(0) <= transition_429_symbol_out;
  place_1296_succs(0) <= transition_434_symbol_out;
  place_1296 : place
    generic map(marking => false)
    port map(
      preds => place_1296_preds,
      succs => place_1296_succs,
      token => place_1296_token,
      clk   => clk,
      reset => reset);

  place_1297_preds(0) <= transition_433_symbol_out;
  place_1297_succs(0) <= transition_435_symbol_out;
  place_1297 : place
    generic map(marking => false)
    port map(
      preds => place_1297_preds,
      succs => place_1297_succs,
      token => place_1297_token,
      clk   => clk,
      reset => reset);

  place_1298_preds(0) <= transition_331_symbol_out;
  place_1298_succs(0) <= transition_431_symbol_out;
  place_1298 : place
    generic map(marking => false)
    port map(
      preds => place_1298_preds,
      succs => place_1298_succs,
      token => place_1298_token,
      clk   => clk,
      reset => reset);

  place_1299_preds(0) <= transition_443_symbol_out;
  place_1299_succs(0) <= transition_436_symbol_out;
  place_1299 : place
    generic map(marking => false)
    port map(
      preds => place_1299_preds,
      succs => place_1299_succs,
      token => place_1299_token,
      clk   => clk,
      reset => reset);

  place_1300_preds(0) <= transition_439_symbol_out;
  place_1300_succs(0) <= transition_444_symbol_out;
  place_1300 : place
    generic map(marking => false)
    port map(
      preds => place_1300_preds,
      succs => place_1300_succs,
      token => place_1300_token,
      clk   => clk,
      reset => reset);

  place_1301_preds(0) <= transition_383_symbol_out;
  place_1301_succs(0) <= transition_443_symbol_out;
  place_1301 : place
    generic map(marking => false)
    port map(
      preds => place_1301_preds,
      succs => place_1301_succs,
      token => place_1301_token,
      clk   => clk,
      reset => reset);

  place_1302_preds(0) <= transition_435_symbol_out;
  place_1302_succs(0) <= transition_443_symbol_out;
  place_1302 : place
    generic map(marking => false)
    port map(
      preds => place_1302_preds,
      succs => place_1302_succs,
      token => place_1302_token,
      clk   => clk,
      reset => reset);

  place_1303_preds(0) <= transition_448_symbol_out;
  place_1303_succs(0) <= transition_466_symbol_out;
  place_1303 : place
    generic map(marking => false)
    port map(
      preds => place_1303_preds,
      succs => place_1303_succs,
      token => place_1303_token,
      clk   => clk,
      reset => reset);

  place_1304_preds(0) <= transition_3_symbol_out;
  place_1304_succs(0) <= transition_445_symbol_out;
  place_1304 : place
    generic map(marking => false)
    port map(
      preds => place_1304_preds,
      succs => place_1304_succs,
      token => place_1304_token,
      clk   => clk,
      reset => reset);

  place_1305_preds(0) <= transition_455_symbol_out;
  place_1305_succs(0) <= transition_466_symbol_out;
  place_1305 : place
    generic map(marking => false)
    port map(
      preds => place_1305_preds,
      succs => place_1305_succs,
      token => place_1305_token,
      clk   => clk,
      reset => reset);

  place_1306_preds(0) <= transition_3_symbol_out;
  place_1306_succs(0) <= transition_452_symbol_out;
  place_1306 : place
    generic map(marking => false)
    port map(
      preds => place_1306_preds,
      succs => place_1306_succs,
      token => place_1306_token,
      clk   => clk,
      reset => reset);

  place_1307_preds(0) <= transition_466_symbol_out;
  place_1307_succs(0) <= transition_459_symbol_out;
  place_1307 : place
    generic map(marking => false)
    port map(
      preds => place_1307_preds,
      succs => place_1307_succs,
      token => place_1307_token,
      clk   => clk,
      reset => reset);

  place_1308_preds(0) <= transition_48_symbol_out;
  place_1308_succs(0) <= transition_55_symbol_out;
  place_1308 : place
    generic map(marking => false)
    port map(
      preds => place_1308_preds,
      succs => place_1308_succs,
      token => place_1308_token,
      clk   => clk,
      reset => reset);

  place_1309_preds(0) <= transition_462_symbol_out;
  place_1309_succs(0) <= transition_481_symbol_out;
  place_1309 : place
    generic map(marking => false)
    port map(
      preds => place_1309_preds,
      succs => place_1309_succs,
      token => place_1309_token,
      clk   => clk,
      reset => reset);

  place_1310_preds(0) <= transition_470_symbol_out;
  place_1310_succs(0) <= transition_481_symbol_out;
  place_1310 : place
    generic map(marking => false)
    port map(
      preds => place_1310_preds,
      succs => place_1310_succs,
      token => place_1310_token,
      clk   => clk,
      reset => reset);

  place_1311_preds(0) <= transition_3_symbol_out;
  place_1311_succs(0) <= transition_467_symbol_out;
  place_1311 : place
    generic map(marking => false)
    port map(
      preds => place_1311_preds,
      succs => place_1311_succs,
      token => place_1311_token,
      clk   => clk,
      reset => reset);

  place_1312_preds(0) <= transition_481_symbol_out;
  place_1312_succs(0) <= transition_474_symbol_out;
  place_1312 : place
    generic map(marking => false)
    port map(
      preds => place_1312_preds,
      succs => place_1312_succs,
      token => place_1312_token,
      clk   => clk,
      reset => reset);

  place_1313_preds(0) <= transition_477_symbol_out;
  place_1313_succs(0) <= transition_482_symbol_out;
  place_1313 : place
    generic map(marking => false)
    port map(
      preds => place_1313_preds,
      succs => place_1313_succs,
      token => place_1313_token,
      clk   => clk,
      reset => reset);

  place_1314_preds(0) <= transition_485_symbol_out;
  place_1314_succs(0) <= transition_492_symbol_out;
  place_1314 : place
    generic map(marking => false)
    port map(
      preds => place_1314_preds,
      succs => place_1314_succs,
      token => place_1314_token,
      clk   => clk,
      reset => reset);

  place_1315_preds(0) <= transition_492_symbol_out;
  place_1315_succs(0) <= transition_491_symbol_out;
  place_1315 : place
    generic map(marking => false)
    port map(
      preds => place_1315_preds,
      succs => place_1315_succs,
      token => place_1315_token,
      clk   => clk,
      reset => reset);

  place_1316_preds(0) <= transition_490_symbol_out;
  place_1316_succs(0) <= transition_555_symbol_out;
  place_1316 : place
    generic map(marking => false)
    port map(
      preds => place_1316_preds,
      succs => place_1316_succs,
      token => place_1316_token,
      clk   => clk,
      reset => reset);

  place_1317_preds(0) <= transition_444_symbol_out;
  place_1317_succs(0) <= transition_492_symbol_out;
  place_1317 : place
    generic map(marking => false)
    port map(
      preds => place_1317_preds,
      succs => place_1317_succs,
      token => place_1317_token,
      clk   => clk,
      reset => reset);

  place_1318_preds(0) <= transition_500_symbol_out;
  place_1318_succs(0) <= transition_493_symbol_out;
  place_1318 : place
    generic map(marking => false)
    port map(
      preds => place_1318_preds,
      succs => place_1318_succs,
      token => place_1318_token,
      clk   => clk,
      reset => reset);

  place_1319_preds(0) <= transition_496_symbol_out;
  place_1319_succs(0) <= transition_501_symbol_out;
  place_1319 : place
    generic map(marking => false)
    port map(
      preds => place_1319_preds,
      succs => place_1319_succs,
      token => place_1319_token,
      clk   => clk,
      reset => reset);

  place_1320_preds(0) <= transition_59_symbol_out;
  place_1320_succs(0) <= transition_500_symbol_out;
  place_1320 : place
    generic map(marking => false)
    port map(
      preds => place_1320_preds,
      succs => place_1320_succs,
      token => place_1320_token,
      clk   => clk,
      reset => reset);

  place_1321_preds(0) <= transition_111_symbol_out;
  place_1321_succs(0) <= transition_500_symbol_out;
  place_1321 : place
    generic map(marking => false)
    port map(
      preds => place_1321_preds,
      succs => place_1321_succs,
      token => place_1321_token,
      clk   => clk,
      reset => reset);

  place_1322_preds(0) <= transition_504_symbol_out;
  place_1322_succs(0) <= transition_555_symbol_out;
  place_1322 : place
    generic map(marking => false)
    port map(
      preds => place_1322_preds,
      succs => place_1322_succs,
      token => place_1322_token,
      clk   => clk,
      reset => reset);

  place_1323_preds(0) <= transition_55_symbol_out;
  place_1323_succs(0) <= transition_54_symbol_out;
  place_1323 : place
    generic map(marking => false)
    port map(
      preds => place_1323_preds,
      succs => place_1323_succs,
      token => place_1323_token,
      clk   => clk,
      reset => reset);

  place_1324_preds(0) <= transition_511_symbol_out;
  place_1324_succs(0) <= transition_529_symbol_out;
  place_1324 : place
    generic map(marking => false)
    port map(
      preds => place_1324_preds,
      succs => place_1324_succs,
      token => place_1324_token,
      clk   => clk,
      reset => reset);

  place_1325_preds(0) <= transition_3_symbol_out;
  place_1325_succs(0) <= transition_508_symbol_out;
  place_1325 : place
    generic map(marking => false)
    port map(
      preds => place_1325_preds,
      succs => place_1325_succs,
      token => place_1325_token,
      clk   => clk,
      reset => reset);

  place_1326_preds(0) <= transition_518_symbol_out;
  place_1326_succs(0) <= transition_529_symbol_out;
  place_1326 : place
    generic map(marking => false)
    port map(
      preds => place_1326_preds,
      succs => place_1326_succs,
      token => place_1326_token,
      clk   => clk,
      reset => reset);

  place_1327_preds(0) <= transition_3_symbol_out;
  place_1327_succs(0) <= transition_515_symbol_out;
  place_1327 : place
    generic map(marking => false)
    port map(
      preds => place_1327_preds,
      succs => place_1327_succs,
      token => place_1327_token,
      clk   => clk,
      reset => reset);

  place_1328_preds(0) <= transition_529_symbol_out;
  place_1328_succs(0) <= transition_522_symbol_out;
  place_1328 : place
    generic map(marking => false)
    port map(
      preds => place_1328_preds,
      succs => place_1328_succs,
      token => place_1328_token,
      clk   => clk,
      reset => reset);

  place_1329_preds(0) <= transition_53_symbol_out;
  place_1329_succs(0) <= transition_58_symbol_out;
  place_1329 : place
    generic map(marking => false)
    port map(
      preds => place_1329_preds,
      succs => place_1329_succs,
      token => place_1329_token,
      clk   => clk,
      reset => reset);

  place_1330_preds(0) <= transition_525_symbol_out;
  place_1330_succs(0) <= transition_544_symbol_out;
  place_1330 : place
    generic map(marking => false)
    port map(
      preds => place_1330_preds,
      succs => place_1330_succs,
      token => place_1330_token,
      clk   => clk,
      reset => reset);

  place_1331_preds(0) <= transition_533_symbol_out;
  place_1331_succs(0) <= transition_544_symbol_out;
  place_1331 : place
    generic map(marking => false)
    port map(
      preds => place_1331_preds,
      succs => place_1331_succs,
      token => place_1331_token,
      clk   => clk,
      reset => reset);

  place_1332_preds(0) <= transition_3_symbol_out;
  place_1332_succs(0) <= transition_530_symbol_out;
  place_1332 : place
    generic map(marking => false)
    port map(
      preds => place_1332_preds,
      succs => place_1332_succs,
      token => place_1332_token,
      clk   => clk,
      reset => reset);

  place_1333_preds(0) <= transition_544_symbol_out;
  place_1333_succs(0) <= transition_537_symbol_out;
  place_1333 : place
    generic map(marking => false)
    port map(
      preds => place_1333_preds,
      succs => place_1333_succs,
      token => place_1333_token,
      clk   => clk,
      reset => reset);

  place_1334_preds(0) <= transition_540_symbol_out;
  place_1334_succs(0) <= transition_545_symbol_out;
  place_1334 : place
    generic map(marking => false)
    port map(
      preds => place_1334_preds,
      succs => place_1334_succs,
      token => place_1334_token,
      clk   => clk,
      reset => reset);

  place_1335_preds(0) <= transition_548_symbol_out;
  place_1335_succs(0) <= transition_555_symbol_out;
  place_1335 : place
    generic map(marking => false)
    port map(
      preds => place_1335_preds,
      succs => place_1335_succs,
      token => place_1335_token,
      clk   => clk,
      reset => reset);

  place_1336_preds(0) <= transition_555_symbol_out;
  place_1336_succs(0) <= transition_554_symbol_out;
  place_1336 : place
    generic map(marking => false)
    port map(
      preds => place_1336_preds,
      succs => place_1336_succs,
      token => place_1336_token,
      clk   => clk,
      reset => reset);

  place_1337_preds(0) <= transition_553_symbol_out;
  place_1337_succs(0) <= transition_618_symbol_out;
  place_1337 : place
    generic map(marking => false)
    port map(
      preds => place_1337_preds,
      succs => place_1337_succs,
      token => place_1337_token,
      clk   => clk,
      reset => reset);

  place_1338_preds(0) <= transition_57_symbol_out;
  place_1338_succs(0) <= transition_59_symbol_out;
  place_1338 : place
    generic map(marking => false)
    port map(
      preds => place_1338_preds,
      succs => place_1338_succs,
      token => place_1338_token,
      clk   => clk,
      reset => reset);

  place_1339_preds(0) <= transition_563_symbol_out;
  place_1339_succs(0) <= transition_556_symbol_out;
  place_1339 : place
    generic map(marking => false)
    port map(
      preds => place_1339_preds,
      succs => place_1339_succs,
      token => place_1339_token,
      clk   => clk,
      reset => reset);

  place_1340_preds(0) <= transition_559_symbol_out;
  place_1340_succs(0) <= transition_564_symbol_out;
  place_1340 : place
    generic map(marking => false)
    port map(
      preds => place_1340_preds,
      succs => place_1340_succs,
      token => place_1340_token,
      clk   => clk,
      reset => reset);

  place_1341_preds(0) <= transition_221_symbol_out;
  place_1341_succs(0) <= transition_563_symbol_out;
  place_1341 : place
    generic map(marking => false)
    port map(
      preds => place_1341_preds,
      succs => place_1341_succs,
      token => place_1341_token,
      clk   => clk,
      reset => reset);

  place_1342_preds(0) <= transition_273_symbol_out;
  place_1342_succs(0) <= transition_563_symbol_out;
  place_1342 : place
    generic map(marking => false)
    port map(
      preds => place_1342_preds,
      succs => place_1342_succs,
      token => place_1342_token,
      clk   => clk,
      reset => reset);

  place_1343_preds(0) <= transition_567_symbol_out;
  place_1343_succs(0) <= transition_618_symbol_out;
  place_1343 : place
    generic map(marking => false)
    port map(
      preds => place_1343_preds,
      succs => place_1343_succs,
      token => place_1343_token,
      clk   => clk,
      reset => reset);

  place_1344_preds(0) <= transition_574_symbol_out;
  place_1344_succs(0) <= transition_592_symbol_out;
  place_1344 : place
    generic map(marking => false)
    port map(
      preds => place_1344_preds,
      succs => place_1344_succs,
      token => place_1344_token,
      clk   => clk,
      reset => reset);

  place_1345_preds(0) <= transition_3_symbol_out;
  place_1345_succs(0) <= transition_571_symbol_out;
  place_1345 : place
    generic map(marking => false)
    port map(
      preds => place_1345_preds,
      succs => place_1345_succs,
      token => place_1345_token,
      clk   => clk,
      reset => reset);

  place_1346_preds(0) <= transition_581_symbol_out;
  place_1346_succs(0) <= transition_592_symbol_out;
  place_1346 : place
    generic map(marking => false)
    port map(
      preds => place_1346_preds,
      succs => place_1346_succs,
      token => place_1346_token,
      clk   => clk,
      reset => reset);

  place_1347_preds(0) <= transition_3_symbol_out;
  place_1347_succs(0) <= transition_578_symbol_out;
  place_1347 : place
    generic map(marking => false)
    port map(
      preds => place_1347_preds,
      succs => place_1347_succs,
      token => place_1347_token,
      clk   => clk,
      reset => reset);

  place_1348_preds(0) <= transition_592_symbol_out;
  place_1348_succs(0) <= transition_585_symbol_out;
  place_1348 : place
    generic map(marking => false)
    port map(
      preds => place_1348_preds,
      succs => place_1348_succs,
      token => place_1348_token,
      clk   => clk,
      reset => reset);

  place_1349_preds(0) <= transition_588_symbol_out;
  place_1349_succs(0) <= transition_607_symbol_out;
  place_1349 : place
    generic map(marking => false)
    port map(
      preds => place_1349_preds,
      succs => place_1349_succs,
      token => place_1349_token,
      clk   => clk,
      reset => reset);

  place_1350_preds(0) <= transition_596_symbol_out;
  place_1350_succs(0) <= transition_607_symbol_out;
  place_1350 : place
    generic map(marking => false)
    port map(
      preds => place_1350_preds,
      succs => place_1350_succs,
      token => place_1350_token,
      clk   => clk,
      reset => reset);

  place_1351_preds(0) <= transition_3_symbol_out;
  place_1351_succs(0) <= transition_593_symbol_out;
  place_1351 : place
    generic map(marking => false)
    port map(
      preds => place_1351_preds,
      succs => place_1351_succs,
      token => place_1351_token,
      clk   => clk,
      reset => reset);

  place_1352_preds(0) <= transition_607_symbol_out;
  place_1352_succs(0) <= transition_600_symbol_out;
  place_1352 : place
    generic map(marking => false)
    port map(
      preds => place_1352_preds,
      succs => place_1352_succs,
      token => place_1352_token,
      clk   => clk,
      reset => reset);

  place_1353_preds(0) <= transition_603_symbol_out;
  place_1353_succs(0) <= transition_608_symbol_out;
  place_1353 : place
    generic map(marking => false)
    port map(
      preds => place_1353_preds,
      succs => place_1353_succs,
      token => place_1353_token,
      clk   => clk,
      reset => reset);

  place_1354_preds(0) <= transition_611_symbol_out;
  place_1354_succs(0) <= transition_618_symbol_out;
  place_1354 : place
    generic map(marking => false)
    port map(
      preds => place_1354_preds,
      succs => place_1354_succs,
      token => place_1354_token,
      clk   => clk,
      reset => reset);

  place_1355_preds(0) <= transition_618_symbol_out;
  place_1355_succs(0) <= transition_617_symbol_out;
  place_1355 : place
    generic map(marking => false)
    port map(
      preds => place_1355_preds,
      succs => place_1355_succs,
      token => place_1355_token,
      clk   => clk,
      reset => reset);

  place_1356_preds(0) <= transition_616_symbol_out;
  place_1356_succs(0) <= transition_681_symbol_out;
  place_1356 : place
    generic map(marking => false)
    port map(
      preds => place_1356_preds,
      succs => place_1356_succs,
      token => place_1356_token,
      clk   => clk,
      reset => reset);

  place_1357_preds(0) <= transition_11_symbol_out;
  place_1357_succs(0) <= transition_29_symbol_out;
  place_1357 : place
    generic map(marking => false)
    port map(
      preds => place_1357_preds,
      succs => place_1357_succs,
      token => place_1357_token,
      clk   => clk,
      reset => reset);

  place_1358_preds(0) <= transition_3_symbol_out;
  place_1358_succs(0) <= transition_55_symbol_out;
  place_1358 : place
    generic map(marking => false)
    port map(
      preds => place_1358_preds,
      succs => place_1358_succs,
      token => place_1358_token,
      clk   => clk,
      reset => reset);

  place_1359_preds(0) <= transition_626_symbol_out;
  place_1359_succs(0) <= transition_619_symbol_out;
  place_1359 : place
    generic map(marking => false)
    port map(
      preds => place_1359_preds,
      succs => place_1359_succs,
      token => place_1359_token,
      clk   => clk,
      reset => reset);

  place_1360_preds(0) <= transition_622_symbol_out;
  place_1360_succs(0) <= transition_627_symbol_out;
  place_1360 : place
    generic map(marking => false)
    port map(
      preds => place_1360_preds,
      succs => place_1360_succs,
      token => place_1360_token,
      clk   => clk,
      reset => reset);

  place_1361_preds(0) <= transition_383_symbol_out;
  place_1361_succs(0) <= transition_626_symbol_out;
  place_1361 : place
    generic map(marking => false)
    port map(
      preds => place_1361_preds,
      succs => place_1361_succs,
      token => place_1361_token,
      clk   => clk,
      reset => reset);

  place_1362_preds(0) <= transition_435_symbol_out;
  place_1362_succs(0) <= transition_626_symbol_out;
  place_1362 : place
    generic map(marking => false)
    port map(
      preds => place_1362_preds,
      succs => place_1362_succs,
      token => place_1362_token,
      clk   => clk,
      reset => reset);

  place_1363_preds(0) <= transition_630_symbol_out;
  place_1363_succs(0) <= transition_681_symbol_out;
  place_1363 : place
    generic map(marking => false)
    port map(
      preds => place_1363_preds,
      succs => place_1363_succs,
      token => place_1363_token,
      clk   => clk,
      reset => reset);

  place_1364_preds(0) <= transition_637_symbol_out;
  place_1364_succs(0) <= transition_655_symbol_out;
  place_1364 : place
    generic map(marking => false)
    port map(
      preds => place_1364_preds,
      succs => place_1364_succs,
      token => place_1364_token,
      clk   => clk,
      reset => reset);

  place_1365_preds(0) <= transition_3_symbol_out;
  place_1365_succs(0) <= transition_634_symbol_out;
  place_1365 : place
    generic map(marking => false)
    port map(
      preds => place_1365_preds,
      succs => place_1365_succs,
      token => place_1365_token,
      clk   => clk,
      reset => reset);

  place_1366_preds(0) <= transition_644_symbol_out;
  place_1366_succs(0) <= transition_655_symbol_out;
  place_1366 : place
    generic map(marking => false)
    port map(
      preds => place_1366_preds,
      succs => place_1366_succs,
      token => place_1366_token,
      clk   => clk,
      reset => reset);

  place_1367_preds(0) <= transition_3_symbol_out;
  place_1367_succs(0) <= transition_641_symbol_out;
  place_1367 : place
    generic map(marking => false)
    port map(
      preds => place_1367_preds,
      succs => place_1367_succs,
      token => place_1367_token,
      clk   => clk,
      reset => reset);

  place_1368_preds(0) <= transition_655_symbol_out;
  place_1368_succs(0) <= transition_648_symbol_out;
  place_1368 : place
    generic map(marking => false)
    port map(
      preds => place_1368_preds,
      succs => place_1368_succs,
      token => place_1368_token,
      clk   => clk,
      reset => reset);

  place_1369_preds(0) <= transition_63_symbol_out;
  place_1369_succs(0) <= transition_81_symbol_out;
  place_1369 : place
    generic map(marking => false)
    port map(
      preds => place_1369_preds,
      succs => place_1369_succs,
      token => place_1369_token,
      clk   => clk,
      reset => reset);

  place_1370_preds(0) <= transition_651_symbol_out;
  place_1370_succs(0) <= transition_670_symbol_out;
  place_1370 : place
    generic map(marking => false)
    port map(
      preds => place_1370_preds,
      succs => place_1370_succs,
      token => place_1370_token,
      clk   => clk,
      reset => reset);

  place_1371_preds(0) <= transition_659_symbol_out;
  place_1371_succs(0) <= transition_670_symbol_out;
  place_1371 : place
    generic map(marking => false)
    port map(
      preds => place_1371_preds,
      succs => place_1371_succs,
      token => place_1371_token,
      clk   => clk,
      reset => reset);

  place_1372_preds(0) <= transition_3_symbol_out;
  place_1372_succs(0) <= transition_656_symbol_out;
  place_1372 : place
    generic map(marking => false)
    port map(
      preds => place_1372_preds,
      succs => place_1372_succs,
      token => place_1372_token,
      clk   => clk,
      reset => reset);

  place_1373_preds(0) <= transition_670_symbol_out;
  place_1373_succs(0) <= transition_663_symbol_out;
  place_1373 : place
    generic map(marking => false)
    port map(
      preds => place_1373_preds,
      succs => place_1373_succs,
      token => place_1373_token,
      clk   => clk,
      reset => reset);

  place_1374_preds(0) <= transition_666_symbol_out;
  place_1374_succs(0) <= transition_671_symbol_out;
  place_1374 : place
    generic map(marking => false)
    port map(
      preds => place_1374_preds,
      succs => place_1374_succs,
      token => place_1374_token,
      clk   => clk,
      reset => reset);

  place_1375_preds(0) <= transition_674_symbol_out;
  place_1375_succs(0) <= transition_681_symbol_out;
  place_1375 : place
    generic map(marking => false)
    port map(
      preds => place_1375_preds,
      succs => place_1375_succs,
      token => place_1375_token,
      clk   => clk,
      reset => reset);

  place_1376_preds(0) <= transition_681_symbol_out;
  place_1376_succs(0) <= transition_680_symbol_out;
  place_1376 : place
    generic map(marking => false)
    port map(
      preds => place_1376_preds,
      succs => place_1376_succs,
      token => place_1376_token,
      clk   => clk,
      reset => reset);

  place_1377_preds(0) <= transition_679_symbol_out;
  place_1377_succs(0) <= transition_682_symbol_out;
  place_1377 : place
    generic map(marking => false)
    port map(
      preds => place_1377_preds,
      succs => place_1377_succs,
      token => place_1377_token,
      clk   => clk,
      reset => reset);

  place_1378_preds(0) <= transition_686_symbol_out;
  place_1378_succs(0) <= transition_704_symbol_out;
  place_1378 : place
    generic map(marking => false)
    port map(
      preds => place_1378_preds,
      succs => place_1378_succs,
      token => place_1378_token,
      clk   => clk,
      reset => reset);

  place_1379_preds(0) <= transition_3_symbol_out;
  place_1379_succs(0) <= transition_683_symbol_out;
  place_1379 : place
    generic map(marking => false)
    port map(
      preds => place_1379_preds,
      succs => place_1379_succs,
      token => place_1379_token,
      clk   => clk,
      reset => reset);

  place_1380_preds(0) <= transition_693_symbol_out;
  place_1380_succs(0) <= transition_704_symbol_out;
  place_1380 : place
    generic map(marking => false)
    port map(
      preds => place_1380_preds,
      succs => place_1380_succs,
      token => place_1380_token,
      clk   => clk,
      reset => reset);

  place_1381_preds(0) <= transition_3_symbol_out;
  place_1381_succs(0) <= transition_690_symbol_out;
  place_1381 : place
    generic map(marking => false)
    port map(
      preds => place_1381_preds,
      succs => place_1381_succs,
      token => place_1381_token,
      clk   => clk,
      reset => reset);

  place_1382_preds(0) <= transition_3_symbol_out;
  place_1382_succs(0) <= transition_60_symbol_out;
  place_1382 : place
    generic map(marking => false)
    port map(
      preds => place_1382_preds,
      succs => place_1382_succs,
      token => place_1382_token,
      clk   => clk,
      reset => reset);

  place_1383_preds(0) <= transition_704_symbol_out;
  place_1383_succs(0) <= transition_697_symbol_out;
  place_1383 : place
    generic map(marking => false)
    port map(
      preds => place_1383_preds,
      succs => place_1383_succs,
      token => place_1383_token,
      clk   => clk,
      reset => reset);

  place_1384_preds(0) <= transition_700_symbol_out;
  place_1384_succs(0) <= transition_719_symbol_out;
  place_1384 : place
    generic map(marking => false)
    port map(
      preds => place_1384_preds,
      succs => place_1384_succs,
      token => place_1384_token,
      clk   => clk,
      reset => reset);

  place_1385_preds(0) <= transition_708_symbol_out;
  place_1385_succs(0) <= transition_719_symbol_out;
  place_1385 : place
    generic map(marking => false)
    port map(
      preds => place_1385_preds,
      succs => place_1385_succs,
      token => place_1385_token,
      clk   => clk,
      reset => reset);

  place_1386_preds(0) <= transition_3_symbol_out;
  place_1386_succs(0) <= transition_705_symbol_out;
  place_1386 : place
    generic map(marking => false)
    port map(
      preds => place_1386_preds,
      succs => place_1386_succs,
      token => place_1386_token,
      clk   => clk,
      reset => reset);

  place_1387_preds(0) <= transition_719_symbol_out;
  place_1387_succs(0) <= transition_712_symbol_out;
  place_1387 : place
    generic map(marking => false)
    port map(
      preds => place_1387_preds,
      succs => place_1387_succs,
      token => place_1387_token,
      clk   => clk,
      reset => reset);

  place_1388_preds(0) <= transition_715_symbol_out;
  place_1388_succs(0) <= transition_720_symbol_out;
  place_1388 : place
    generic map(marking => false)
    port map(
      preds => place_1388_preds,
      succs => place_1388_succs,
      token => place_1388_token,
      clk   => clk,
      reset => reset);

  place_1389_preds(0) <= transition_723_symbol_out;
  place_1389_succs(0) <= transition_730_symbol_out;
  place_1389 : place
    generic map(marking => false)
    port map(
      preds => place_1389_preds,
      succs => place_1389_succs,
      token => place_1389_token,
      clk   => clk,
      reset => reset);

  place_1390_preds(0) <= transition_730_symbol_out;
  place_1390_succs(0) <= transition_729_symbol_out;
  place_1390 : place
    generic map(marking => false)
    port map(
      preds => place_1390_preds,
      succs => place_1390_succs,
      token => place_1390_token,
      clk   => clk,
      reset => reset);

  place_1391_preds(0) <= transition_70_symbol_out;
  place_1391_succs(0) <= transition_81_symbol_out;
  place_1391 : place
    generic map(marking => false)
    port map(
      preds => place_1391_preds,
      succs => place_1391_succs,
      token => place_1391_token,
      clk   => clk,
      reset => reset);

  place_1392_preds(0) <= transition_728_symbol_out;
  place_1392_succs(0) <= transition_733_symbol_out;
  place_1392 : place
    generic map(marking => false)
    port map(
      preds => place_1392_preds,
      succs => place_1392_succs,
      token => place_1392_token,
      clk   => clk,
      reset => reset);

  place_1393_preds(0) <= transition_732_symbol_out;
  place_1393_succs(0) <= transition_792_symbol_out;
  place_1393 : place
    generic map(marking => false)
    port map(
      preds => place_1393_preds,
      succs => place_1393_succs,
      token => place_1393_token,
      clk   => clk,
      reset => reset);

  place_1394_preds(0) <= transition_682_symbol_out;
  place_1394_succs(0) <= transition_730_symbol_out;
  place_1394 : place
    generic map(marking => false)
    port map(
      preds => place_1394_preds,
      succs => place_1394_succs,
      token => place_1394_token,
      clk   => clk,
      reset => reset);

  place_1395_preds(0) <= transition_737_symbol_out;
  place_1395_succs(0) <= transition_755_symbol_out;
  place_1395 : place
    generic map(marking => false)
    port map(
      preds => place_1395_preds,
      succs => place_1395_succs,
      token => place_1395_token,
      clk   => clk,
      reset => reset);

  place_1396_preds(0) <= transition_3_symbol_out;
  place_1396_succs(0) <= transition_734_symbol_out;
  place_1396 : place
    generic map(marking => false)
    port map(
      preds => place_1396_preds,
      succs => place_1396_succs,
      token => place_1396_token,
      clk   => clk,
      reset => reset);

  place_1397_preds(0) <= transition_744_symbol_out;
  place_1397_succs(0) <= transition_755_symbol_out;
  place_1397 : place
    generic map(marking => false)
    port map(
      preds => place_1397_preds,
      succs => place_1397_succs,
      token => place_1397_token,
      clk   => clk,
      reset => reset);

  place_1398_preds(0) <= transition_3_symbol_out;
  place_1398_succs(0) <= transition_741_symbol_out;
  place_1398 : place
    generic map(marking => false)
    port map(
      preds => place_1398_preds,
      succs => place_1398_succs,
      token => place_1398_token,
      clk   => clk,
      reset => reset);

  place_1399_preds(0) <= transition_755_symbol_out;
  place_1399_succs(0) <= transition_748_symbol_out;
  place_1399 : place
    generic map(marking => false)
    port map(
      preds => place_1399_preds,
      succs => place_1399_succs,
      token => place_1399_token,
      clk   => clk,
      reset => reset);

  place_1400_preds(0) <= transition_751_symbol_out;
  place_1400_succs(0) <= transition_770_symbol_out;
  place_1400 : place
    generic map(marking => false)
    port map(
      preds => place_1400_preds,
      succs => place_1400_succs,
      token => place_1400_token,
      clk   => clk,
      reset => reset);

  place_1401_preds(0) <= transition_3_symbol_out;
  place_1401_succs(0) <= transition_67_symbol_out;
  place_1401 : place
    generic map(marking => false)
    port map(
      preds => place_1401_preds,
      succs => place_1401_succs,
      token => place_1401_token,
      clk   => clk,
      reset => reset);

  place_1402_preds(0) <= transition_759_symbol_out;
  place_1402_succs(0) <= transition_770_symbol_out;
  place_1402 : place
    generic map(marking => false)
    port map(
      preds => place_1402_preds,
      succs => place_1402_succs,
      token => place_1402_token,
      clk   => clk,
      reset => reset);

  place_1403_preds(0) <= transition_3_symbol_out;
  place_1403_succs(0) <= transition_756_symbol_out;
  place_1403 : place
    generic map(marking => false)
    port map(
      preds => place_1403_preds,
      succs => place_1403_succs,
      token => place_1403_token,
      clk   => clk,
      reset => reset);

  place_1404_preds(0) <= transition_770_symbol_out;
  place_1404_succs(0) <= transition_763_symbol_out;
  place_1404 : place
    generic map(marking => false)
    port map(
      preds => place_1404_preds,
      succs => place_1404_succs,
      token => place_1404_token,
      clk   => clk,
      reset => reset);

  place_1405_preds(0) <= transition_766_symbol_out;
  place_1405_succs(0) <= transition_771_symbol_out;
  place_1405 : place
    generic map(marking => false)
    port map(
      preds => place_1405_preds,
      succs => place_1405_succs,
      token => place_1405_token,
      clk   => clk,
      reset => reset);

  place_1406_preds(0) <= transition_81_symbol_out;
  place_1406_succs(0) <= transition_74_symbol_out;
  place_1406 : place
    generic map(marking => false)
    port map(
      preds => place_1406_preds,
      succs => place_1406_succs,
      token => place_1406_token,
      clk   => clk,
      reset => reset);

  place_1407_preds(0) <= transition_774_symbol_out;
  place_1407_succs(0) <= transition_781_symbol_out;
  place_1407 : place
    generic map(marking => false)
    port map(
      preds => place_1407_preds,
      succs => place_1407_succs,
      token => place_1407_token,
      clk   => clk,
      reset => reset);

  place_1408_preds(0) <= transition_781_symbol_out;
  place_1408_succs(0) <= transition_780_symbol_out;
  place_1408 : place
    generic map(marking => false)
    port map(
      preds => place_1408_preds,
      succs => place_1408_succs,
      token => place_1408_token,
      clk   => clk,
      reset => reset);

  place_1409_preds(0) <= transition_779_symbol_out;
  place_1409_succs(0) <= transition_784_symbol_out;
  place_1409 : place
    generic map(marking => false)
    port map(
      preds => place_1409_preds,
      succs => place_1409_succs,
      token => place_1409_token,
      clk   => clk,
      reset => reset);

  place_1410_preds(0) <= transition_783_symbol_out;
  place_1410_succs(0) <= transition_792_symbol_out;
  place_1410 : place
    generic map(marking => false)
    port map(
      preds => place_1410_preds,
      succs => place_1410_succs,
      token => place_1410_token,
      clk   => clk,
      reset => reset);

  place_1411_preds(0) <= transition_77_symbol_out;
  place_1411_succs(0) <= transition_96_symbol_out;
  place_1411 : place
    generic map(marking => false)
    port map(
      preds => place_1411_preds,
      succs => place_1411_succs,
      token => place_1411_token,
      clk   => clk,
      reset => reset);

  place_1412_preds(0) <= transition_682_symbol_out;
  place_1412_succs(0) <= transition_781_symbol_out;
  place_1412 : place
    generic map(marking => false)
    port map(
      preds => place_1412_preds,
      succs => place_1412_succs,
      token => place_1412_token,
      clk   => clk,
      reset => reset);

  place_1413_preds(0) <= transition_792_symbol_out;
  place_1413_succs(0) <= transition_785_symbol_out;
  place_1413 : place
    generic map(marking => false)
    port map(
      preds => place_1413_preds,
      succs => place_1413_succs,
      token => place_1413_token,
      clk   => clk,
      reset => reset);

  place_1414_preds(0) <= transition_788_symbol_out;
  place_1414_succs(0) <= transition_793_symbol_out;
  place_1414 : place
    generic map(marking => false)
    port map(
      preds => place_1414_preds,
      succs => place_1414_succs,
      token => place_1414_token,
      clk   => clk,
      reset => reset);

  place_1415_preds(0) <= transition_796_symbol_out;
  place_1415_succs(0) <= transition_847_symbol_out;
  place_1415 : place
    generic map(marking => false)
    port map(
      preds => place_1415_preds,
      succs => place_1415_succs,
      token => place_1415_token,
      clk   => clk,
      reset => reset);

  place_1416_preds(0) <= transition_803_symbol_out;
  place_1416_succs(0) <= transition_821_symbol_out;
  place_1416 : place
    generic map(marking => false)
    port map(
      preds => place_1416_preds,
      succs => place_1416_succs,
      token => place_1416_token,
      clk   => clk,
      reset => reset);

  place_1417_preds(0) <= transition_3_symbol_out;
  place_1417_succs(0) <= transition_800_symbol_out;
  place_1417 : place
    generic map(marking => false)
    port map(
      preds => place_1417_preds,
      succs => place_1417_succs,
      token => place_1417_token,
      clk   => clk,
      reset => reset);

  place_1418_preds(0) <= transition_810_symbol_out;
  place_1418_succs(0) <= transition_821_symbol_out;
  place_1418 : place
    generic map(marking => false)
    port map(
      preds => place_1418_preds,
      succs => place_1418_succs,
      token => place_1418_token,
      clk   => clk,
      reset => reset);

  place_1419_preds(0) <= transition_3_symbol_out;
  place_1419_succs(0) <= transition_807_symbol_out;
  place_1419 : place
    generic map(marking => false)
    port map(
      preds => place_1419_preds,
      succs => place_1419_succs,
      token => place_1419_token,
      clk   => clk,
      reset => reset);

  place_1420_preds(0) <= transition_821_symbol_out;
  place_1420_succs(0) <= transition_814_symbol_out;
  place_1420 : place
    generic map(marking => false)
    port map(
      preds => place_1420_preds,
      succs => place_1420_succs,
      token => place_1420_token,
      clk   => clk,
      reset => reset);

  place_1421_preds(0) <= transition_817_symbol_out;
  place_1421_succs(0) <= transition_836_symbol_out;
  place_1421 : place
    generic map(marking => false)
    port map(
      preds => place_1421_preds,
      succs => place_1421_succs,
      token => place_1421_token,
      clk   => clk,
      reset => reset);

  place_1422_preds(0) <= transition_825_symbol_out;
  place_1422_succs(0) <= transition_836_symbol_out;
  place_1422 : place
    generic map(marking => false)
    port map(
      preds => place_1422_preds,
      succs => place_1422_succs,
      token => place_1422_token,
      clk   => clk,
      reset => reset);

  place_1423_preds(0) <= transition_3_symbol_out;
  place_1423_succs(0) <= transition_822_symbol_out;
  place_1423 : place
    generic map(marking => false)
    port map(
      preds => place_1423_preds,
      succs => place_1423_succs,
      token => place_1423_token,
      clk   => clk,
      reset => reset);

  place_1424_preds(0) <= transition_836_symbol_out;
  place_1424_succs(0) <= transition_829_symbol_out;
  place_1424 : place
    generic map(marking => false)
    port map(
      preds => place_1424_preds,
      succs => place_1424_succs,
      token => place_1424_token,
      clk   => clk,
      reset => reset);

  place_1425_preds(0) <= transition_832_symbol_out;
  place_1425_succs(0) <= transition_837_symbol_out;
  place_1425 : place
    generic map(marking => false)
    port map(
      preds => place_1425_preds,
      succs => place_1425_succs,
      token => place_1425_token,
      clk   => clk,
      reset => reset);

  place_1426_preds(0) <= transition_840_symbol_out;
  place_1426_succs(0) <= transition_847_symbol_out;
  place_1426 : place
    generic map(marking => false)
    port map(
      preds => place_1426_preds,
      succs => place_1426_succs,
      token => place_1426_token,
      clk   => clk,
      reset => reset);

  place_1427_preds(0) <= transition_847_symbol_out;
  place_1427_succs(0) <= transition_846_symbol_out;
  place_1427 : place
    generic map(marking => false)
    port map(
      preds => place_1427_preds,
      succs => place_1427_succs,
      token => place_1427_token,
      clk   => clk,
      reset => reset);

  place_1428_preds(0) <= transition_845_symbol_out;
  place_1428_succs(0) <= transition_848_symbol_out;
  place_1428 : place
    generic map(marking => false)
    port map(
      preds => place_1428_preds,
      succs => place_1428_succs,
      token => place_1428_token,
      clk   => clk,
      reset => reset);

  place_1429_preds(0) <= transition_852_symbol_out;
  place_1429_succs(0) <= transition_870_symbol_out;
  place_1429 : place
    generic map(marking => false)
    port map(
      preds => place_1429_preds,
      succs => place_1429_succs,
      token => place_1429_token,
      clk   => clk,
      reset => reset);

  place_1430_preds(0) <= transition_3_symbol_out;
  place_1430_succs(0) <= transition_849_symbol_out;
  place_1430 : place
    generic map(marking => false)
    port map(
      preds => place_1430_preds,
      succs => place_1430_succs,
      token => place_1430_token,
      clk   => clk,
      reset => reset);

  place_1431_preds(0) <= transition_859_symbol_out;
  place_1431_succs(0) <= transition_870_symbol_out;
  place_1431 : place
    generic map(marking => false)
    port map(
      preds => place_1431_preds,
      succs => place_1431_succs,
      token => place_1431_token,
      clk   => clk,
      reset => reset);

  place_1432_preds(0) <= transition_3_symbol_out;
  place_1432_succs(0) <= transition_856_symbol_out;
  place_1432 : place
    generic map(marking => false)
    port map(
      preds => place_1432_preds,
      succs => place_1432_succs,
      token => place_1432_token,
      clk   => clk,
      reset => reset);

  place_1433_preds(0) <= transition_870_symbol_out;
  place_1433_succs(0) <= transition_863_symbol_out;
  place_1433 : place
    generic map(marking => false)
    port map(
      preds => place_1433_preds,
      succs => place_1433_succs,
      token => place_1433_token,
      clk   => clk,
      reset => reset);

  place_1434_preds(0) <= transition_866_symbol_out;
  place_1434_succs(0) <= transition_885_symbol_out;
  place_1434 : place
    generic map(marking => false)
    port map(
      preds => place_1434_preds,
      succs => place_1434_succs,
      token => place_1434_token,
      clk   => clk,
      reset => reset);

  place_1435_preds(0) <= transition_85_symbol_out;
  place_1435_succs(0) <= transition_96_symbol_out;
  place_1435 : place
    generic map(marking => false)
    port map(
      preds => place_1435_preds,
      succs => place_1435_succs,
      token => place_1435_token,
      clk   => clk,
      reset => reset);

  place_1436_preds(0) <= transition_874_symbol_out;
  place_1436_succs(0) <= transition_885_symbol_out;
  place_1436 : place
    generic map(marking => false)
    port map(
      preds => place_1436_preds,
      succs => place_1436_succs,
      token => place_1436_token,
      clk   => clk,
      reset => reset);

  place_1437_preds(0) <= transition_3_symbol_out;
  place_1437_succs(0) <= transition_871_symbol_out;
  place_1437 : place
    generic map(marking => false)
    port map(
      preds => place_1437_preds,
      succs => place_1437_succs,
      token => place_1437_token,
      clk   => clk,
      reset => reset);

  place_1438_preds(0) <= transition_885_symbol_out;
  place_1438_succs(0) <= transition_878_symbol_out;
  place_1438 : place
    generic map(marking => false)
    port map(
      preds => place_1438_preds,
      succs => place_1438_succs,
      token => place_1438_token,
      clk   => clk,
      reset => reset);

  place_1439_preds(0) <= transition_881_symbol_out;
  place_1439_succs(0) <= transition_886_symbol_out;
  place_1439 : place
    generic map(marking => false)
    port map(
      preds => place_1439_preds,
      succs => place_1439_succs,
      token => place_1439_token,
      clk   => clk,
      reset => reset);

  place_1440_preds(0) <= transition_889_symbol_out;
  place_1440_succs(0) <= transition_896_symbol_out;
  place_1440 : place
    generic map(marking => false)
    port map(
      preds => place_1440_preds,
      succs => place_1440_succs,
      token => place_1440_token,
      clk   => clk,
      reset => reset);

  place_1441_preds(0) <= transition_896_symbol_out;
  place_1441_succs(0) <= transition_895_symbol_out;
  place_1441 : place
    generic map(marking => false)
    port map(
      preds => place_1441_preds,
      succs => place_1441_succs,
      token => place_1441_token,
      clk   => clk,
      reset => reset);

  place_1442_preds(0) <= transition_894_symbol_out;
  place_1442_succs(0) <= transition_899_symbol_out;
  place_1442 : place
    generic map(marking => false)
    port map(
      preds => place_1442_preds,
      succs => place_1442_succs,
      token => place_1442_token,
      clk   => clk,
      reset => reset);

  place_1443_preds(0) <= transition_898_symbol_out;
  place_1443_succs(0) <= transition_958_symbol_out;
  place_1443 : place
    generic map(marking => false)
    port map(
      preds => place_1443_preds,
      succs => place_1443_succs,
      token => place_1443_token,
      clk   => clk,
      reset => reset);

  place_1444_preds(0) <= transition_3_symbol_out;
  place_1444_succs(0) <= transition_82_symbol_out;
  place_1444 : place
    generic map(marking => false)
    port map(
      preds => place_1444_preds,
      succs => place_1444_succs,
      token => place_1444_token,
      clk   => clk,
      reset => reset);

  place_1445_preds(0) <= transition_848_symbol_out;
  place_1445_succs(0) <= transition_896_symbol_out;
  place_1445 : place
    generic map(marking => false)
    port map(
      preds => place_1445_preds,
      succs => place_1445_succs,
      token => place_1445_token,
      clk   => clk,
      reset => reset);

  place_1446_preds(0) <= transition_903_symbol_out;
  place_1446_succs(0) <= transition_921_symbol_out;
  place_1446 : place
    generic map(marking => false)
    port map(
      preds => place_1446_preds,
      succs => place_1446_succs,
      token => place_1446_token,
      clk   => clk,
      reset => reset);

  place_1447_preds(0) <= transition_3_symbol_out;
  place_1447_succs(0) <= transition_900_symbol_out;
  place_1447 : place
    generic map(marking => false)
    port map(
      preds => place_1447_preds,
      succs => place_1447_succs,
      token => place_1447_token,
      clk   => clk,
      reset => reset);

  place_1448_preds(0) <= transition_910_symbol_out;
  place_1448_succs(0) <= transition_921_symbol_out;
  place_1448 : place
    generic map(marking => false)
    port map(
      preds => place_1448_preds,
      succs => place_1448_succs,
      token => place_1448_token,
      clk   => clk,
      reset => reset);

  place_1449_preds(0) <= transition_96_symbol_out;
  place_1449_succs(0) <= transition_89_symbol_out;
  place_1449 : place
    generic map(marking => false)
    port map(
      preds => place_1449_preds,
      succs => place_1449_succs,
      token => place_1449_token,
      clk   => clk,
      reset => reset);

  place_1450_preds(0) <= transition_3_symbol_out;
  place_1450_succs(0) <= transition_907_symbol_out;
  place_1450 : place
    generic map(marking => false)
    port map(
      preds => place_1450_preds,
      succs => place_1450_succs,
      token => place_1450_token,
      clk   => clk,
      reset => reset);

  place_1451_preds(0) <= transition_921_symbol_out;
  place_1451_succs(0) <= transition_914_symbol_out;
  place_1451 : place
    generic map(marking => false)
    port map(
      preds => place_1451_preds,
      succs => place_1451_succs,
      token => place_1451_token,
      clk   => clk,
      reset => reset);

  place_1452_preds(0) <= transition_917_symbol_out;
  place_1452_succs(0) <= transition_936_symbol_out;
  place_1452 : place
    generic map(marking => false)
    port map(
      preds => place_1452_preds,
      succs => place_1452_succs,
      token => place_1452_token,
      clk   => clk,
      reset => reset);

  place_1453_preds(0) <= transition_925_symbol_out;
  place_1453_succs(0) <= transition_936_symbol_out;
  place_1453 : place
    generic map(marking => false)
    port map(
      preds => place_1453_preds,
      succs => place_1453_succs,
      token => place_1453_token,
      clk   => clk,
      reset => reset);

  place_1454_preds(0) <= transition_92_symbol_out;
  place_1454_succs(0) <= transition_97_symbol_out;
  place_1454 : place
    generic map(marking => false)
    port map(
      preds => place_1454_preds,
      succs => place_1454_succs,
      token => place_1454_token,
      clk   => clk,
      reset => reset);

  place_1455_preds(0) <= transition_3_symbol_out;
  place_1455_succs(0) <= transition_922_symbol_out;
  place_1455 : place
    generic map(marking => false)
    port map(
      preds => place_1455_preds,
      succs => place_1455_succs,
      token => place_1455_token,
      clk   => clk,
      reset => reset);

  place_1456_preds(0) <= transition_936_symbol_out;
  place_1456_succs(0) <= transition_929_symbol_out;
  place_1456 : place
    generic map(marking => false)
    port map(
      preds => place_1456_preds,
      succs => place_1456_succs,
      token => place_1456_token,
      clk   => clk,
      reset => reset);

  place_1457_preds(0) <= transition_932_symbol_out;
  place_1457_succs(0) <= transition_937_symbol_out;
  place_1457 : place
    generic map(marking => false)
    port map(
      preds => place_1457_preds,
      succs => place_1457_succs,
      token => place_1457_token,
      clk   => clk,
      reset => reset);

  place_1458_preds(0) <= transition_940_symbol_out;
  place_1458_succs(0) <= transition_947_symbol_out;
  place_1458 : place
    generic map(marking => false)
    port map(
      preds => place_1458_preds,
      succs => place_1458_succs,
      token => place_1458_token,
      clk   => clk,
      reset => reset);

  place_1459_preds(0) <= transition_947_symbol_out;
  place_1459_succs(0) <= transition_946_symbol_out;
  place_1459 : place
    generic map(marking => false)
    port map(
      preds => place_1459_preds,
      succs => place_1459_succs,
      token => place_1459_token,
      clk   => clk,
      reset => reset);

  place_1460_preds(0) <= transition_945_symbol_out;
  place_1460_succs(0) <= transition_950_symbol_out;
  place_1460 : place
    generic map(marking => false)
    port map(
      preds => place_1460_preds,
      succs => place_1460_succs,
      token => place_1460_token,
      clk   => clk,
      reset => reset);

  place_1461_preds(0) <= transition_949_symbol_out;
  place_1461_succs(0) <= transition_958_symbol_out;
  place_1461 : place
    generic map(marking => false)
    port map(
      preds => place_1461_preds,
      succs => place_1461_succs,
      token => place_1461_token,
      clk   => clk,
      reset => reset);

  place_1462_preds(0) <= transition_848_symbol_out;
  place_1462_succs(0) <= transition_947_symbol_out;
  place_1462 : place
    generic map(marking => false)
    port map(
      preds => place_1462_preds,
      succs => place_1462_succs,
      token => place_1462_token,
      clk   => clk,
      reset => reset);

  place_1463_preds(0) <= transition_958_symbol_out;
  place_1463_succs(0) <= transition_951_symbol_out;
  place_1463 : place
    generic map(marking => false)
    port map(
      preds => place_1463_preds,
      succs => place_1463_succs,
      token => place_1463_token,
      clk   => clk,
      reset => reset);

  place_1464_preds(0) <= transition_954_symbol_out;
  place_1464_succs(0) <= transition_959_symbol_out;
  place_1464 : place
    generic map(marking => false)
    port map(
      preds => place_1464_preds,
      succs => place_1464_succs,
      token => place_1464_token,
      clk   => clk,
      reset => reset);

  place_1465_preds(0) <= transition_962_symbol_out;
  place_1465_succs(0) <= transition_1013_symbol_out;
  place_1465 : place
    generic map(marking => false)
    port map(
      preds => place_1465_preds,
      succs => place_1465_succs,
      token => place_1465_token,
      clk   => clk,
      reset => reset);

  place_1466_preds(0) <= transition_969_symbol_out;
  place_1466_succs(0) <= transition_987_symbol_out;
  place_1466 : place
    generic map(marking => false)
    port map(
      preds => place_1466_preds,
      succs => place_1466_succs,
      token => place_1466_token,
      clk   => clk,
      reset => reset);

  place_1467_preds(0) <= transition_3_symbol_out;
  place_1467_succs(0) <= transition_966_symbol_out;
  place_1467 : place
    generic map(marking => false)
    port map(
      preds => place_1467_preds,
      succs => place_1467_succs,
      token => place_1467_token,
      clk   => clk,
      reset => reset);

  place_1468_preds(0) <= transition_976_symbol_out;
  place_1468_succs(0) <= transition_987_symbol_out;
  place_1468 : place
    generic map(marking => false)
    port map(
      preds => place_1468_preds,
      succs => place_1468_succs,
      token => place_1468_token,
      clk   => clk,
      reset => reset);

  place_1469_preds(0) <= transition_3_symbol_out;
  place_1469_succs(0) <= transition_973_symbol_out;
  place_1469 : place
    generic map(marking => false)
    port map(
      preds => place_1469_preds,
      succs => place_1469_succs,
      token => place_1469_token,
      clk   => clk,
      reset => reset);

  place_1470_preds(0) <= transition_987_symbol_out;
  place_1470_succs(0) <= transition_980_symbol_out;
  place_1470 : place
    generic map(marking => false)
    port map(
      preds => place_1470_preds,
      succs => place_1470_succs,
      token => place_1470_token,
      clk   => clk,
      reset => reset);

  place_1471_preds(0) <= transition_983_symbol_out;
  place_1471_succs(0) <= transition_1002_symbol_out;
  place_1471 : place
    generic map(marking => false)
    port map(
      preds => place_1471_preds,
      succs => place_1471_succs,
      token => place_1471_token,
      clk   => clk,
      reset => reset);

  place_1472_preds(0) <= transition_991_symbol_out;
  place_1472_succs(0) <= transition_1002_symbol_out;
  place_1472 : place
    generic map(marking => false)
    port map(
      preds => place_1472_preds,
      succs => place_1472_succs,
      token => place_1472_token,
      clk   => clk,
      reset => reset);

  place_1473_preds(0) <= transition_3_symbol_out;
  place_1473_succs(0) <= transition_988_symbol_out;
  place_1473 : place
    generic map(marking => false)
    port map(
      preds => place_1473_preds,
      succs => place_1473_succs,
      token => place_1473_token,
      clk   => clk,
      reset => reset);

  place_1474_preds(0) <= transition_1002_symbol_out;
  place_1474_succs(0) <= transition_995_symbol_out;
  place_1474 : place
    generic map(marking => false)
    port map(
      preds => place_1474_preds,
      succs => place_1474_succs,
      token => place_1474_token,
      clk   => clk,
      reset => reset);

  place_1475_preds(0) <= transition_998_symbol_out;
  place_1475_succs(0) <= transition_1003_symbol_out;
  place_1475 : place
    generic map(marking => false)
    port map(
      preds => place_1475_preds,
      succs => place_1475_succs,
      token => place_1475_token,
      clk   => clk,
      reset => reset);

  place_1476_preds(0) <= transition_100_symbol_out;
  place_1476_succs(0) <= transition_107_symbol_out;
  place_1476 : place
    generic map(marking => false)
    port map(
      preds => place_1476_preds,
      succs => place_1476_succs,
      token => place_1476_token,
      clk   => clk,
      reset => reset);

  place_1477_preds(0) <= transition_1006_symbol_out;
  place_1477_succs(0) <= transition_1013_symbol_out;
  place_1477 : place
    generic map(marking => false)
    port map(
      preds => place_1477_preds,
      succs => place_1477_succs,
      token => place_1477_token,
      clk   => clk,
      reset => reset);

  place_1478_preds(0) <= transition_1013_symbol_out;
  place_1478_succs(0) <= transition_1012_symbol_out;
  place_1478 : place
    generic map(marking => false)
    port map(
      preds => place_1478_preds,
      succs => place_1478_succs,
      token => place_1478_token,
      clk   => clk,
      reset => reset);

  place_1479_preds(0) <= transition_1011_symbol_out;
  place_1479_succs(0) <= transition_1014_symbol_out;
  place_1479 : place
    generic map(marking => false)
    port map(
      preds => place_1479_preds,
      succs => place_1479_succs,
      token => place_1479_token,
      clk   => clk,
      reset => reset);

  place_1480_preds(0) <= transition_1018_symbol_out;
  place_1480_succs(0) <= transition_1036_symbol_out;
  place_1480 : place
    generic map(marking => false)
    port map(
      preds => place_1480_preds,
      succs => place_1480_succs,
      token => place_1480_token,
      clk   => clk,
      reset => reset);

  place_1481_preds(0) <= transition_3_symbol_out;
  place_1481_succs(0) <= transition_1015_symbol_out;
  place_1481 : place
    generic map(marking => false)
    port map(
      preds => place_1481_preds,
      succs => place_1481_succs,
      token => place_1481_token,
      clk   => clk,
      reset => reset);

  place_1482_preds(0) <= transition_1025_symbol_out;
  place_1482_succs(0) <= transition_1036_symbol_out;
  place_1482 : place
    generic map(marking => false)
    port map(
      preds => place_1482_preds,
      succs => place_1482_succs,
      token => place_1482_token,
      clk   => clk,
      reset => reset);

  place_1483_preds(0) <= transition_3_symbol_out;
  place_1483_succs(0) <= transition_1022_symbol_out;
  place_1483 : place
    generic map(marking => false)
    port map(
      preds => place_1483_preds,
      succs => place_1483_succs,
      token => place_1483_token,
      clk   => clk,
      reset => reset);

  place_1484_preds(0) <= transition_1036_symbol_out;
  place_1484_succs(0) <= transition_1029_symbol_out;
  place_1484 : place
    generic map(marking => false)
    port map(
      preds => place_1484_preds,
      succs => place_1484_succs,
      token => place_1484_token,
      clk   => clk,
      reset => reset);

  place_1485_preds(0) <= transition_1032_symbol_out;
  place_1485_succs(0) <= transition_1051_symbol_out;
  place_1485 : place
    generic map(marking => false)
    port map(
      preds => place_1485_preds,
      succs => place_1485_succs,
      token => place_1485_token,
      clk   => clk,
      reset => reset);

  place_1486_preds(0) <= transition_1040_symbol_out;
  place_1486_succs(0) <= transition_1051_symbol_out;
  place_1486 : place
    generic map(marking => false)
    port map(
      preds => place_1486_preds,
      succs => place_1486_succs,
      token => place_1486_token,
      clk   => clk,
      reset => reset);

  place_1487_preds(0) <= transition_3_symbol_out;
  place_1487_succs(0) <= transition_1037_symbol_out;
  place_1487 : place
    generic map(marking => false)
    port map(
      preds => place_1487_preds,
      succs => place_1487_succs,
      token => place_1487_token,
      clk   => clk,
      reset => reset);

  place_1488_preds(0) <= transition_1051_symbol_out;
  place_1488_succs(0) <= transition_1044_symbol_out;
  place_1488 : place
    generic map(marking => false)
    port map(
      preds => place_1488_preds,
      succs => place_1488_succs,
      token => place_1488_token,
      clk   => clk,
      reset => reset);

  place_1489_preds(0) <= transition_1047_symbol_out;
  place_1489_succs(0) <= transition_1052_symbol_out;
  place_1489 : place
    generic map(marking => false)
    port map(
      preds => place_1489_preds,
      succs => place_1489_succs,
      token => place_1489_token,
      clk   => clk,
      reset => reset);

  place_1490_preds(0) <= transition_107_symbol_out;
  place_1490_succs(0) <= transition_106_symbol_out;
  place_1490 : place
    generic map(marking => false)
    port map(
      preds => place_1490_preds,
      succs => place_1490_succs,
      token => place_1490_token,
      clk   => clk,
      reset => reset);

  place_1491_preds(0) <= transition_1055_symbol_out;
  place_1491_succs(0) <= transition_1062_symbol_out;
  place_1491 : place
    generic map(marking => false)
    port map(
      preds => place_1491_preds,
      succs => place_1491_succs,
      token => place_1491_token,
      clk   => clk,
      reset => reset);

  place_1492_preds(0) <= transition_1062_symbol_out;
  place_1492_succs(0) <= transition_1061_symbol_out;
  place_1492 : place
    generic map(marking => false)
    port map(
      preds => place_1492_preds,
      succs => place_1492_succs,
      token => place_1492_token,
      clk   => clk,
      reset => reset);

  place_1493_preds(0) <= transition_1060_symbol_out;
  place_1493_succs(0) <= transition_1065_symbol_out;
  place_1493 : place
    generic map(marking => false)
    port map(
      preds => place_1493_preds,
      succs => place_1493_succs,
      token => place_1493_token,
      clk   => clk,
      reset => reset);

  place_1494_preds(0) <= transition_1064_symbol_out;
  place_1494_succs(0) <= transition_1124_symbol_out;
  place_1494 : place
    generic map(marking => false)
    port map(
      preds => place_1494_preds,
      succs => place_1494_succs,
      token => place_1494_token,
      clk   => clk,
      reset => reset);

  place_1495_preds(0) <= transition_105_symbol_out;
  place_1495_succs(0) <= transition_110_symbol_out;
  place_1495 : place
    generic map(marking => false)
    port map(
      preds => place_1495_preds,
      succs => place_1495_succs,
      token => place_1495_token,
      clk   => clk,
      reset => reset);

  place_1496_preds(0) <= transition_1014_symbol_out;
  place_1496_succs(0) <= transition_1062_symbol_out;
  place_1496 : place
    generic map(marking => false)
    port map(
      preds => place_1496_preds,
      succs => place_1496_succs,
      token => place_1496_token,
      clk   => clk,
      reset => reset);

  place_1497_preds(0) <= transition_1069_symbol_out;
  place_1497_succs(0) <= transition_1087_symbol_out;
  place_1497 : place
    generic map(marking => false)
    port map(
      preds => place_1497_preds,
      succs => place_1497_succs,
      token => place_1497_token,
      clk   => clk,
      reset => reset);

  place_1498_preds(0) <= transition_3_symbol_out;
  place_1498_succs(0) <= transition_1066_symbol_out;
  place_1498 : place
    generic map(marking => false)
    port map(
      preds => place_1498_preds,
      succs => place_1498_succs,
      token => place_1498_token,
      clk   => clk,
      reset => reset);

  place_1499_preds(0) <= transition_1076_symbol_out;
  place_1499_succs(0) <= transition_1087_symbol_out;
  place_1499 : place
    generic map(marking => false)
    port map(
      preds => place_1499_preds,
      succs => place_1499_succs,
      token => place_1499_token,
      clk   => clk,
      reset => reset);

  place_1500_preds(0) <= transition_3_symbol_out;
  place_1500_succs(0) <= transition_1073_symbol_out;
  place_1500 : place
    generic map(marking => false)
    port map(
      preds => place_1500_preds,
      succs => place_1500_succs,
      token => place_1500_token,
      clk   => clk,
      reset => reset);

  place_1501_preds(0) <= transition_3_symbol_out;
  place_1501_succs(0) <= transition_8_symbol_out;
  place_1501 : place
    generic map(marking => false)
    port map(
      preds => place_1501_preds,
      succs => place_1501_succs,
      token => place_1501_token,
      clk   => clk,
      reset => reset);

  place_1502_preds(0) <= transition_1087_symbol_out;
  place_1502_succs(0) <= transition_1080_symbol_out;
  place_1502 : place
    generic map(marking => false)
    port map(
      preds => place_1502_preds,
      succs => place_1502_succs,
      token => place_1502_token,
      clk   => clk,
      reset => reset);

  place_1503_preds(0) <= transition_1083_symbol_out;
  place_1503_succs(0) <= transition_1102_symbol_out;
  place_1503 : place
    generic map(marking => false)
    port map(
      preds => place_1503_preds,
      succs => place_1503_succs,
      token => place_1503_token,
      clk   => clk,
      reset => reset);

  place_1504_preds(0) <= transition_1091_symbol_out;
  place_1504_succs(0) <= transition_1102_symbol_out;
  place_1504 : place
    generic map(marking => false)
    port map(
      preds => place_1504_preds,
      succs => place_1504_succs,
      token => place_1504_token,
      clk   => clk,
      reset => reset);

  place_1505_preds(0) <= transition_3_symbol_out;
  place_1505_succs(0) <= transition_1088_symbol_out;
  place_1505 : place
    generic map(marking => false)
    port map(
      preds => place_1505_preds,
      succs => place_1505_succs,
      token => place_1505_token,
      clk   => clk,
      reset => reset);

  place_1506_preds(0) <= transition_1102_symbol_out;
  place_1506_succs(0) <= transition_1095_symbol_out;
  place_1506 : place
    generic map(marking => false)
    port map(
      preds => place_1506_preds,
      succs => place_1506_succs,
      token => place_1506_token,
      clk   => clk,
      reset => reset);

  place_1507_preds(0) <= transition_109_symbol_out;
  place_1507_succs(0) <= transition_111_symbol_out;
  place_1507 : place
    generic map(marking => false)
    port map(
      preds => place_1507_preds,
      succs => place_1507_succs,
      token => place_1507_token,
      clk   => clk,
      reset => reset);

  place_1508_preds(0) <= transition_1098_symbol_out;
  place_1508_succs(0) <= transition_1103_symbol_out;
  place_1508 : place
    generic map(marking => false)
    port map(
      preds => place_1508_preds,
      succs => place_1508_succs,
      token => place_1508_token,
      clk   => clk,
      reset => reset);

  place_1509_preds(0) <= transition_1106_symbol_out;
  place_1509_succs(0) <= transition_1113_symbol_out;
  place_1509 : place
    generic map(marking => false)
    port map(
      preds => place_1509_preds,
      succs => place_1509_succs,
      token => place_1509_token,
      clk   => clk,
      reset => reset);

  place_1510_preds(0) <= transition_1113_symbol_out;
  place_1510_succs(0) <= transition_1112_symbol_out;
  place_1510 : place
    generic map(marking => false)
    port map(
      preds => place_1510_preds,
      succs => place_1510_succs,
      token => place_1510_token,
      clk   => clk,
      reset => reset);

  place_1511_preds(0) <= transition_1111_symbol_out;
  place_1511_succs(0) <= transition_1116_symbol_out;
  place_1511 : place
    generic map(marking => false)
    port map(
      preds => place_1511_preds,
      succs => place_1511_succs,
      token => place_1511_token,
      clk   => clk,
      reset => reset);

  place_1512_preds(0) <= transition_1115_symbol_out;
  place_1512_succs(0) <= transition_1124_symbol_out;
  place_1512 : place
    generic map(marking => false)
    port map(
      preds => place_1512_preds,
      succs => place_1512_succs,
      token => place_1512_token,
      clk   => clk,
      reset => reset);

  place_1513_preds(0) <= transition_1014_symbol_out;
  place_1513_succs(0) <= transition_1113_symbol_out;
  place_1513 : place
    generic map(marking => false)
    port map(
      preds => place_1513_preds,
      succs => place_1513_succs,
      token => place_1513_token,
      clk   => clk,
      reset => reset);

  place_1514_preds(0) <= transition_1124_symbol_out;
  place_1514_succs(0) <= transition_1117_symbol_out;
  place_1514 : place
    generic map(marking => false)
    port map(
      preds => place_1514_preds,
      succs => place_1514_succs,
      token => place_1514_token,
      clk   => clk,
      reset => reset);

  place_1515_preds(0) <= transition_1120_symbol_out;
  place_1515_succs(0) <= transition_1125_symbol_out;
  place_1515 : place
    generic map(marking => false)
    port map(
      preds => place_1515_preds,
      succs => place_1515_succs,
      token => place_1515_token,
      clk   => clk,
      reset => reset);

  place_1516_preds(0) <= transition_1128_symbol_out;
  place_1516_succs(0) <= transition_1179_symbol_out;
  place_1516 : place
    generic map(marking => false)
    port map(
      preds => place_1516_preds,
      succs => place_1516_succs,
      token => place_1516_token,
      clk   => clk,
      reset => reset);

  place_1517_preds(0) <= transition_1135_symbol_out;
  place_1517_succs(0) <= transition_1153_symbol_out;
  place_1517 : place
    generic map(marking => false)
    port map(
      preds => place_1517_preds,
      succs => place_1517_succs,
      token => place_1517_token,
      clk   => clk,
      reset => reset);

  place_1518_preds(0) <= transition_3_symbol_out;
  place_1518_succs(0) <= transition_1132_symbol_out;
  place_1518 : place
    generic map(marking => false)
    port map(
      preds => place_1518_preds,
      succs => place_1518_succs,
      token => place_1518_token,
      clk   => clk,
      reset => reset);

  place_1519_preds(0) <= transition_1142_symbol_out;
  place_1519_succs(0) <= transition_1153_symbol_out;
  place_1519 : place
    generic map(marking => false)
    port map(
      preds => place_1519_preds,
      succs => place_1519_succs,
      token => place_1519_token,
      clk   => clk,
      reset => reset);

  place_1520_preds(0) <= transition_3_symbol_out;
  place_1520_succs(0) <= transition_1139_symbol_out;
  place_1520 : place
    generic map(marking => false)
    port map(
      preds => place_1520_preds,
      succs => place_1520_succs,
      token => place_1520_token,
      clk   => clk,
      reset => reset);

  place_1521_preds(0) <= transition_1153_symbol_out;
  place_1521_succs(0) <= transition_1146_symbol_out;
  place_1521 : place
    generic map(marking => false)
    port map(
      preds => place_1521_preds,
      succs => place_1521_succs,
      token => place_1521_token,
      clk   => clk,
      reset => reset);

  place_1522_preds(0) <= transition_1149_symbol_out;
  place_1522_succs(0) <= transition_1168_symbol_out;
  place_1522 : place
    generic map(marking => false)
    port map(
      preds => place_1522_preds,
      succs => place_1522_succs,
      token => place_1522_token,
      clk   => clk,
      reset => reset);

  place_1523_preds(0) <= transition_1157_symbol_out;
  place_1523_succs(0) <= transition_1168_symbol_out;
  place_1523 : place
    generic map(marking => false)
    port map(
      preds => place_1523_preds,
      succs => place_1523_succs,
      token => place_1523_token,
      clk   => clk,
      reset => reset);

  place_1524_preds(0) <= transition_3_symbol_out;
  place_1524_succs(0) <= transition_107_symbol_out;
  place_1524 : place
    generic map(marking => false)
    port map(
      preds => place_1524_preds,
      succs => place_1524_succs,
      token => place_1524_token,
      clk   => clk,
      reset => reset);

  place_1525_preds(0) <= transition_3_symbol_out;
  place_1525_succs(0) <= transition_1154_symbol_out;
  place_1525 : place
    generic map(marking => false)
    port map(
      preds => place_1525_preds,
      succs => place_1525_succs,
      token => place_1525_token,
      clk   => clk,
      reset => reset);

  place_1526_preds(0) <= transition_1168_symbol_out;
  place_1526_succs(0) <= transition_1161_symbol_out;
  place_1526 : place
    generic map(marking => false)
    port map(
      preds => place_1526_preds,
      succs => place_1526_succs,
      token => place_1526_token,
      clk   => clk,
      reset => reset);

  place_1527_preds(0) <= transition_1164_symbol_out;
  place_1527_succs(0) <= transition_1169_symbol_out;
  place_1527 : place
    generic map(marking => false)
    port map(
      preds => place_1527_preds,
      succs => place_1527_succs,
      token => place_1527_token,
      clk   => clk,
      reset => reset);

  place_1528_preds(0) <= transition_1172_symbol_out;
  place_1528_succs(0) <= transition_1179_symbol_out;
  place_1528 : place
    generic map(marking => false)
    port map(
      preds => place_1528_preds,
      succs => place_1528_succs,
      token => place_1528_token,
      clk   => clk,
      reset => reset);

  place_1529_preds(0) <= transition_119_symbol_out;
  place_1529_succs(0) <= transition_112_symbol_out;
  place_1529 : place
    generic map(marking => false)
    port map(
      preds => place_1529_preds,
      succs => place_1529_succs,
      token => place_1529_token,
      clk   => clk,
      reset => reset);

  place_1530_preds(0) <= transition_1179_symbol_out;
  place_1530_succs(0) <= transition_1178_symbol_out;
  place_1530 : place
    generic map(marking => false)
    port map(
      preds => place_1530_preds,
      succs => place_1530_succs,
      token => place_1530_token,
      clk   => clk,
      reset => reset);

  place_1531_preds(0) <= transition_1177_symbol_out;
  place_1531_succs(0) <= transition_4_symbol_out;
  place_1531 : place
    generic map(marking => false)
    port map(
      preds => place_1531_preds,
      succs => place_1531_succs,
      token => place_1531_token,
      clk   => clk,
      reset => reset);

  place_1532_preds(0) <= transition_1187_symbol_out;
  place_1532_succs(0) <= transition_1180_symbol_out;
  place_1532 : place
    generic map(marking => false)
    port map(
      preds => place_1532_preds,
      succs => place_1532_succs,
      token => place_1532_token,
      clk   => clk,
      reset => reset);

  place_1533_preds(0) <= transition_1183_symbol_out;
  place_1533_succs(0) <= transition_1195_symbol_out;
  place_1533 : place
    generic map(marking => false)
    port map(
      preds => place_1533_preds,
      succs => place_1533_succs,
      token => place_1533_token,
      clk   => clk,
      reset => reset);

  place_1534_preds(0) <= transition_282_symbol_out;
  place_1534_succs(0) <= transition_1187_symbol_out;
  place_1534 : place
    generic map(marking => false)
    port map(
      preds => place_1534_preds,
      succs => place_1534_succs,
      token => place_1534_token,
      clk   => clk,
      reset => reset);

  place_1535_preds(0) <= transition_120_symbol_out;
  place_1535_succs(0) <= transition_1187_symbol_out;
  place_1535 : place
    generic map(marking => false)
    port map(
      preds => place_1535_preds,
      succs => place_1535_succs,
      token => place_1535_token,
      clk   => clk,
      reset => reset);

  place_1536_preds(0) <= transition_115_symbol_out;
  place_1536_succs(0) <= transition_120_symbol_out;
  place_1536 : place
    generic map(marking => false)
    port map(
      preds => place_1536_preds,
      succs => place_1536_succs,
      token => place_1536_token,
      clk   => clk,
      reset => reset);

  place_1537_preds(0) <= transition_1195_symbol_out;
  place_1537_succs(0) <= transition_1188_symbol_out;
  place_1537 : place
    generic map(marking => false)
    port map(
      preds => place_1537_preds,
      succs => place_1537_succs,
      token => place_1537_token,
      clk   => clk,
      reset => reset);

  place_1538_preds(0) <= transition_1191_symbol_out;
  place_1538_succs(0) <= transition_1196_symbol_out;
  place_1538 : place
    generic map(marking => false)
    port map(
      preds => place_1538_preds,
      succs => place_1538_succs,
      token => place_1538_token,
      clk   => clk,
      reset => reset);

  place_1539_preds(0) <= transition_444_symbol_out;
  place_1539_succs(0) <= transition_1195_symbol_out;
  place_1539 : place
    generic map(marking => false)
    port map(
      preds => place_1539_preds,
      succs => place_1539_succs,
      token => place_1539_token,
      clk   => clk,
      reset => reset);

  place_1540_preds(0) <= transition_1199_symbol_out;
  place_1540_succs(0) <= transition_4_symbol_out;
  place_1540 : place
    generic map(marking => false)
    port map(
      preds => place_1540_preds,
      succs => place_1540_succs,
      token => place_1540_token,
      clk   => clk,
      reset => reset);

  place_1541_preds(0) <= transition_4_symbol_out;
  place_1541_succs(0) <= transition_1205_symbol_out;
  place_1541 : place
    generic map(marking => false)
    port map(
      preds => place_1541_preds,
      succs => place_1541_succs,
      token => place_1541_token,
      clk   => clk,
      reset => reset);

  place_1542_preds(0) <= transition_1204_symbol_out;
  place_1542_succs(0) <= transition_2_symbol_out;
  place_1542 : place
    generic map(marking => false)
    port map(
      preds => place_1542_preds,
      succs => place_1542_succs,
      token => place_1542_token,
      clk   => clk,
      reset => reset);

  place_1543_preds(0) <= transition_59_symbol_out;
  place_1543_succs(0) <= transition_119_symbol_out;
  place_1543 : place
    generic map(marking => false)
    port map(
      preds => place_1543_preds,
      succs => place_1543_succs,
      token => place_1543_token,
      clk   => clk,
      reset => reset);

  place_1544_preds(0) <= transition_111_symbol_out;
  place_1544_succs(0) <= transition_119_symbol_out;
  place_1544 : place
    generic map(marking => false)
    port map(
      preds => place_1544_preds,
      succs => place_1544_succs,
      token => place_1544_token,
      clk   => clk,
      reset => reset);

  place_1545_preds(0) <= transition_124_symbol_out;
  place_1545_succs(0) <= transition_142_symbol_out;
  place_1545 : place
    generic map(marking => false)
    port map(
      preds => place_1545_preds,
      succs => place_1545_succs,
      token => place_1545_token,
      clk   => clk,
      reset => reset);

  place_1546_preds(0) <= transition_3_symbol_out;
  place_1546_succs(0) <= transition_121_symbol_out;
  place_1546 : place
    generic map(marking => false)
    port map(
      preds => place_1546_preds,
      succs => place_1546_succs,
      token => place_1546_token,
      clk   => clk,
      reset => reset);

  place_1547_preds(0) <= transition_131_symbol_out;
  place_1547_succs(0) <= transition_142_symbol_out;
  place_1547 : place
    generic map(marking => false)
    port map(
      preds => place_1547_preds,
      succs => place_1547_succs,
      token => place_1547_token,
      clk   => clk,
      reset => reset);

  place_1548_preds(0) <= transition_18_symbol_out;
  place_1548_succs(0) <= transition_29_symbol_out;
  place_1548 : place
    generic map(marking => false)
    port map(
      preds => place_1548_preds,
      succs => place_1548_succs,
      token => place_1548_token,
      clk   => clk,
      reset => reset);

  place_1549_preds(0) <= transition_3_symbol_out;
  place_1549_succs(0) <= transition_128_symbol_out;
  place_1549 : place
    generic map(marking => false)
    port map(
      preds => place_1549_preds,
      succs => place_1549_succs,
      token => place_1549_token,
      clk   => clk,
      reset => reset);

  place_1550_preds(0) <= transition_142_symbol_out;
  place_1550_succs(0) <= transition_135_symbol_out;
  place_1550 : place
    generic map(marking => false)
    port map(
      preds => place_1550_preds,
      succs => place_1550_succs,
      token => place_1550_token,
      clk   => clk,
      reset => reset);

  place_1551_preds(0) <= transition_138_symbol_out;
  place_1551_succs(0) <= transition_157_symbol_out;
  place_1551 : place
    generic map(marking => false)
    port map(
      preds => place_1551_preds,
      succs => place_1551_succs,
      token => place_1551_token,
      clk   => clk,
      reset => reset);

  place_1552_preds(0) <= transition_146_symbol_out;
  place_1552_succs(0) <= transition_157_symbol_out;
  place_1552 : place
    generic map(marking => false)
    port map(
      preds => place_1552_preds,
      succs => place_1552_succs,
      token => place_1552_token,
      clk   => clk,
      reset => reset);

  place_1553_preds(0) <= transition_3_symbol_out;
  place_1553_succs(0) <= transition_143_symbol_out;
  place_1553 : place
    generic map(marking => false)
    port map(
      preds => place_1553_preds,
      succs => place_1553_succs,
      token => place_1553_token,
      clk   => clk,
      reset => reset);

  transition_1_preds(0) <= place_0_token;
  transition_1 : transition
    port map(
      preds      => transition_1_preds,
      symbol_out => transition_1_symbol_out,
      symbol_in  => true);

  transition_2_preds(0) <= place_1542_token;
  transition_2 : transition
    port map(
      preds      => transition_2_preds,
      symbol_out => transition_2_symbol_out,
      symbol_in  => true);

  transition_3_preds(0) <= place_1256_token;
  transition_3 : transition
    port map(
      preds      => transition_3_preds,
      symbol_out => transition_3_symbol_out,
      symbol_in  => true);

  transition_4_preds(0) <= place_1531_token;
  transition_4_preds(1) <= place_1540_token;
  transition_4 : transition
    port map(
      preds      => transition_4_preds,
      symbol_out => transition_4_symbol_out,
      symbol_in  => true);

  transition_6_preds(0) <= place_5_token;
  transition_6 : transition
    port map(
      preds      => transition_6_preds,
      symbol_out => transition_6_symbol_out,
      symbol_in  => LambdaIn(1));

  transition_7_preds(0) <= place_1206_token;
  LambdaOut(1) <= transition_7_symbol_out;
  transition_7 : transition
    port map(
      preds      => transition_7_preds,
      symbol_out => transition_7_symbol_out,
      symbol_in  => true);

  transition_8_preds(0) <= place_1501_token;
  LambdaOut(2) <= transition_8_symbol_out;
  transition_8 : transition
    port map(
      preds      => transition_8_preds,
      symbol_out => transition_8_symbol_out,
      symbol_in  => true);

  transition_9_preds(0) <= place_12_token;
  transition_9 : transition
    port map(
      preds      => transition_9_preds,
      symbol_out => transition_9_symbol_out,
      symbol_in  => LambdaIn(2));

  transition_10_preds(0) <= place_13_token;
  LambdaOut(3) <= transition_10_symbol_out;
  transition_10 : transition
    port map(
      preds      => transition_10_preds,
      symbol_out => transition_10_symbol_out,
      symbol_in  => true);

  transition_11_preds(0) <= place_14_token;
  transition_11 : transition
    port map(
      preds      => transition_11_preds,
      symbol_out => transition_11_symbol_out,
      symbol_in  => LambdaIn(3));

  transition_15_preds(0) <= place_1220_token;
  LambdaOut(4) <= transition_15_symbol_out;
  transition_15 : transition
    port map(
      preds      => transition_15_preds,
      symbol_out => transition_15_symbol_out,
      symbol_in  => true);

  transition_16_preds(0) <= place_19_token;
  transition_16 : transition
    port map(
      preds      => transition_16_preds,
      symbol_out => transition_16_symbol_out,
      symbol_in  => LambdaIn(4));

  transition_17_preds(0) <= place_20_token;
  LambdaOut(5) <= transition_17_symbol_out;
  transition_17 : transition
    port map(
      preds      => transition_17_preds,
      symbol_out => transition_17_symbol_out,
      symbol_in  => true);

  transition_18_preds(0) <= place_21_token;
  transition_18 : transition
    port map(
      preds      => transition_18_preds,
      symbol_out => transition_18_symbol_out,
      symbol_in  => LambdaIn(5));

  transition_22_preds(0) <= place_1225_token;
  LambdaOut(6) <= transition_22_symbol_out;
  transition_22 : transition
    port map(
      preds      => transition_22_preds,
      symbol_out => transition_22_symbol_out,
      symbol_in  => true);

  transition_23_preds(0) <= place_26_token;
  transition_23 : transition
    port map(
      preds      => transition_23_preds,
      symbol_out => transition_23_symbol_out,
      symbol_in  => LambdaIn(6));

  transition_24_preds(0) <= place_27_token;
  LambdaOut(7) <= transition_24_symbol_out;
  transition_24 : transition
    port map(
      preds      => transition_24_preds,
      symbol_out => transition_24_symbol_out,
      symbol_in  => true);

  transition_25_preds(0) <= place_28_token;
  transition_25 : transition
    port map(
      preds      => transition_25_preds,
      symbol_out => transition_25_symbol_out,
      symbol_in  => LambdaIn(7));

  transition_29_preds(0) <= place_1357_token;
  transition_29_preds(1) <= place_1548_token;
  transition_29 : transition
    port map(
      preds      => transition_29_preds,
      symbol_out => transition_29_symbol_out,
      symbol_in  => true);

  transition_30_preds(0) <= place_1272_token;
  LambdaOut(8) <= transition_30_symbol_out;
  transition_30 : transition
    port map(
      preds      => transition_30_preds,
      symbol_out => transition_30_symbol_out,
      symbol_in  => true);

  transition_31_preds(0) <= place_34_token;
  transition_31 : transition
    port map(
      preds      => transition_31_preds,
      symbol_out => transition_31_symbol_out,
      symbol_in  => LambdaIn(8));

  transition_32_preds(0) <= place_35_token;
  LambdaOut(9) <= transition_32_symbol_out;
  transition_32 : transition
    port map(
      preds      => transition_32_preds,
      symbol_out => transition_32_symbol_out,
      symbol_in  => true);

  transition_33_preds(0) <= place_36_token;
  transition_33 : transition
    port map(
      preds      => transition_33_preds,
      symbol_out => transition_33_symbol_out,
      symbol_in  => LambdaIn(9));

  transition_37_preds(0) <= place_1277_token;
  LambdaOut(10) <= transition_37_symbol_out;
  transition_37 : transition
    port map(
      preds      => transition_37_preds,
      symbol_out => transition_37_symbol_out,
      symbol_in  => true);

  transition_38_preds(0) <= place_41_token;
  transition_38 : transition
    port map(
      preds      => transition_38_preds,
      symbol_out => transition_38_symbol_out,
      symbol_in  => LambdaIn(10));

  transition_39_preds(0) <= place_42_token;
  LambdaOut(11) <= transition_39_symbol_out;
  transition_39 : transition
    port map(
      preds      => transition_39_preds,
      symbol_out => transition_39_symbol_out,
      symbol_in  => true);

  transition_40_preds(0) <= place_43_token;
  transition_40 : transition
    port map(
      preds      => transition_40_preds,
      symbol_out => transition_40_symbol_out,
      symbol_in  => LambdaIn(11));

  transition_44_preds(0) <= place_1231_token;
  transition_44_preds(1) <= place_1257_token;
  transition_44 : transition
    port map(
      preds      => transition_44_preds,
      symbol_out => transition_44_symbol_out,
      symbol_in  => true);

  transition_45_preds(0) <= place_1282_token;
  LambdaOut(12) <= transition_45_symbol_out;
  transition_45 : transition
    port map(
      preds      => transition_45_preds,
      symbol_out => transition_45_symbol_out,
      symbol_in  => true);

  transition_46_preds(0) <= place_49_token;
  transition_46 : transition
    port map(
      preds      => transition_46_preds,
      symbol_out => transition_46_symbol_out,
      symbol_in  => LambdaIn(12));

  transition_47_preds(0) <= place_50_token;
  LambdaOut(13) <= transition_47_symbol_out;
  transition_47 : transition
    port map(
      preds      => transition_47_preds,
      symbol_out => transition_47_symbol_out,
      symbol_in  => true);

  transition_48_preds(0) <= place_51_token;
  transition_48 : transition
    port map(
      preds      => transition_48_preds,
      symbol_out => transition_48_symbol_out,
      symbol_in  => LambdaIn(13));

  transition_53_preds(0) <= place_52_token;
  transition_53 : transition
    port map(
      preds      => transition_53_preds,
      symbol_out => transition_53_symbol_out,
      symbol_in  => LambdaIn(14));

  transition_54_preds(0) <= place_1323_token;
  LambdaOut(14) <= transition_54_symbol_out;
  transition_54 : transition
    port map(
      preds      => transition_54_preds,
      symbol_out => transition_54_symbol_out,
      symbol_in  => true);

  transition_55_preds(0) <= place_1308_token;
  transition_55_preds(1) <= place_1358_token;
  transition_55 : transition
    port map(
      preds      => transition_55_preds,
      symbol_out => transition_55_symbol_out,
      symbol_in  => true);

  transition_57_preds(0) <= place_56_token;
  transition_57 : transition
    port map(
      preds      => transition_57_preds,
      symbol_out => transition_57_symbol_out,
      symbol_in  => LambdaIn(15));

  transition_58_preds(0) <= place_1329_token;
  LambdaOut(15) <= transition_58_symbol_out;
  transition_58 : transition
    port map(
      preds      => transition_58_preds,
      symbol_out => transition_58_symbol_out,
      symbol_in  => true);

  transition_59_preds(0) <= place_1338_token;
  transition_59 : transition
    port map(
      preds      => transition_59_preds,
      symbol_out => transition_59_symbol_out,
      symbol_in  => true);

  transition_60_preds(0) <= place_1382_token;
  LambdaOut(16) <= transition_60_symbol_out;
  transition_60 : transition
    port map(
      preds      => transition_60_preds,
      symbol_out => transition_60_symbol_out,
      symbol_in  => true);

  transition_61_preds(0) <= place_64_token;
  transition_61 : transition
    port map(
      preds      => transition_61_preds,
      symbol_out => transition_61_symbol_out,
      symbol_in  => LambdaIn(16));

  transition_62_preds(0) <= place_65_token;
  LambdaOut(17) <= transition_62_symbol_out;
  transition_62 : transition
    port map(
      preds      => transition_62_preds,
      symbol_out => transition_62_symbol_out,
      symbol_in  => true);

  transition_63_preds(0) <= place_66_token;
  transition_63 : transition
    port map(
      preds      => transition_63_preds,
      symbol_out => transition_63_symbol_out,
      symbol_in  => LambdaIn(17));

  transition_67_preds(0) <= place_1401_token;
  LambdaOut(18) <= transition_67_symbol_out;
  transition_67 : transition
    port map(
      preds      => transition_67_preds,
      symbol_out => transition_67_symbol_out,
      symbol_in  => true);

  transition_68_preds(0) <= place_71_token;
  transition_68 : transition
    port map(
      preds      => transition_68_preds,
      symbol_out => transition_68_symbol_out,
      symbol_in  => LambdaIn(18));

  transition_69_preds(0) <= place_72_token;
  LambdaOut(19) <= transition_69_symbol_out;
  transition_69 : transition
    port map(
      preds      => transition_69_preds,
      symbol_out => transition_69_symbol_out,
      symbol_in  => true);

  transition_70_preds(0) <= place_73_token;
  transition_70 : transition
    port map(
      preds      => transition_70_preds,
      symbol_out => transition_70_symbol_out,
      symbol_in  => LambdaIn(19));

  transition_74_preds(0) <= place_1406_token;
  LambdaOut(20) <= transition_74_symbol_out;
  transition_74 : transition
    port map(
      preds      => transition_74_preds,
      symbol_out => transition_74_symbol_out,
      symbol_in  => true);

  transition_75_preds(0) <= place_78_token;
  transition_75 : transition
    port map(
      preds      => transition_75_preds,
      symbol_out => transition_75_symbol_out,
      symbol_in  => LambdaIn(20));

  transition_76_preds(0) <= place_79_token;
  LambdaOut(21) <= transition_76_symbol_out;
  transition_76 : transition
    port map(
      preds      => transition_76_preds,
      symbol_out => transition_76_symbol_out,
      symbol_in  => true);

  transition_77_preds(0) <= place_80_token;
  transition_77 : transition
    port map(
      preds      => transition_77_preds,
      symbol_out => transition_77_symbol_out,
      symbol_in  => LambdaIn(21));

  transition_81_preds(0) <= place_1369_token;
  transition_81_preds(1) <= place_1391_token;
  transition_81 : transition
    port map(
      preds      => transition_81_preds,
      symbol_out => transition_81_symbol_out,
      symbol_in  => true);

  transition_82_preds(0) <= place_1444_token;
  LambdaOut(22) <= transition_82_symbol_out;
  transition_82 : transition
    port map(
      preds      => transition_82_preds,
      symbol_out => transition_82_symbol_out,
      symbol_in  => true);

  transition_83_preds(0) <= place_86_token;
  transition_83 : transition
    port map(
      preds      => transition_83_preds,
      symbol_out => transition_83_symbol_out,
      symbol_in  => LambdaIn(22));

  transition_84_preds(0) <= place_87_token;
  LambdaOut(23) <= transition_84_symbol_out;
  transition_84 : transition
    port map(
      preds      => transition_84_preds,
      symbol_out => transition_84_symbol_out,
      symbol_in  => true);

  transition_85_preds(0) <= place_88_token;
  transition_85 : transition
    port map(
      preds      => transition_85_preds,
      symbol_out => transition_85_symbol_out,
      symbol_in  => LambdaIn(23));

  transition_89_preds(0) <= place_1449_token;
  LambdaOut(24) <= transition_89_symbol_out;
  transition_89 : transition
    port map(
      preds      => transition_89_preds,
      symbol_out => transition_89_symbol_out,
      symbol_in  => true);

  transition_90_preds(0) <= place_93_token;
  transition_90 : transition
    port map(
      preds      => transition_90_preds,
      symbol_out => transition_90_symbol_out,
      symbol_in  => LambdaIn(24));

  transition_91_preds(0) <= place_94_token;
  LambdaOut(25) <= transition_91_symbol_out;
  transition_91 : transition
    port map(
      preds      => transition_91_preds,
      symbol_out => transition_91_symbol_out,
      symbol_in  => true);

  transition_92_preds(0) <= place_95_token;
  transition_92 : transition
    port map(
      preds      => transition_92_preds,
      symbol_out => transition_92_symbol_out,
      symbol_in  => LambdaIn(25));

  transition_96_preds(0) <= place_1411_token;
  transition_96_preds(1) <= place_1435_token;
  transition_96 : transition
    port map(
      preds      => transition_96_preds,
      symbol_out => transition_96_symbol_out,
      symbol_in  => true);

  transition_97_preds(0) <= place_1454_token;
  LambdaOut(26) <= transition_97_symbol_out;
  transition_97 : transition
    port map(
      preds      => transition_97_preds,
      symbol_out => transition_97_symbol_out,
      symbol_in  => true);

  transition_98_preds(0) <= place_101_token;
  transition_98 : transition
    port map(
      preds      => transition_98_preds,
      symbol_out => transition_98_symbol_out,
      symbol_in  => LambdaIn(26));

  transition_99_preds(0) <= place_102_token;
  LambdaOut(27) <= transition_99_symbol_out;
  transition_99 : transition
    port map(
      preds      => transition_99_preds,
      symbol_out => transition_99_symbol_out,
      symbol_in  => true);

  transition_100_preds(0) <= place_103_token;
  transition_100 : transition
    port map(
      preds      => transition_100_preds,
      symbol_out => transition_100_symbol_out,
      symbol_in  => LambdaIn(27));

  transition_105_preds(0) <= place_104_token;
  transition_105 : transition
    port map(
      preds      => transition_105_preds,
      symbol_out => transition_105_symbol_out,
      symbol_in  => LambdaIn(28));

  transition_106_preds(0) <= place_1490_token;
  LambdaOut(28) <= transition_106_symbol_out;
  transition_106 : transition
    port map(
      preds      => transition_106_preds,
      symbol_out => transition_106_symbol_out,
      symbol_in  => true);

  transition_107_preds(0) <= place_1476_token;
  transition_107_preds(1) <= place_1524_token;
  transition_107 : transition
    port map(
      preds      => transition_107_preds,
      symbol_out => transition_107_symbol_out,
      symbol_in  => true);

  transition_109_preds(0) <= place_108_token;
  transition_109 : transition
    port map(
      preds      => transition_109_preds,
      symbol_out => transition_109_symbol_out,
      symbol_in  => LambdaIn(29));

  transition_110_preds(0) <= place_1495_token;
  LambdaOut(29) <= transition_110_symbol_out;
  transition_110 : transition
    port map(
      preds      => transition_110_preds,
      symbol_out => transition_110_symbol_out,
      symbol_in  => true);

  transition_111_preds(0) <= place_1507_token;
  transition_111 : transition
    port map(
      preds      => transition_111_preds,
      symbol_out => transition_111_symbol_out,
      symbol_in  => true);

  transition_112_preds(0) <= place_1529_token;
  LambdaOut(30) <= transition_112_symbol_out;
  transition_112 : transition
    port map(
      preds      => transition_112_preds,
      symbol_out => transition_112_symbol_out,
      symbol_in  => true);

  transition_113_preds(0) <= place_116_token;
  transition_113 : transition
    port map(
      preds      => transition_113_preds,
      symbol_out => transition_113_symbol_out,
      symbol_in  => LambdaIn(30));

  transition_114_preds(0) <= place_117_token;
  LambdaOut(31) <= transition_114_symbol_out;
  transition_114 : transition
    port map(
      preds      => transition_114_preds,
      symbol_out => transition_114_symbol_out,
      symbol_in  => true);

  transition_115_preds(0) <= place_118_token;
  transition_115 : transition
    port map(
      preds      => transition_115_preds,
      symbol_out => transition_115_symbol_out,
      symbol_in  => LambdaIn(31));

  transition_119_preds(0) <= place_1544_token;
  transition_119_preds(1) <= place_1543_token;
  transition_119 : transition
    port map(
      preds      => transition_119_preds,
      symbol_out => transition_119_symbol_out,
      symbol_in  => true);

  transition_120_preds(0) <= place_1536_token;
  transition_120 : transition
    port map(
      preds      => transition_120_preds,
      symbol_out => transition_120_symbol_out,
      symbol_in  => true);

  transition_121_preds(0) <= place_1546_token;
  LambdaOut(32) <= transition_121_symbol_out;
  transition_121 : transition
    port map(
      preds      => transition_121_preds,
      symbol_out => transition_121_symbol_out,
      symbol_in  => true);

  transition_122_preds(0) <= place_125_token;
  transition_122 : transition
    port map(
      preds      => transition_122_preds,
      symbol_out => transition_122_symbol_out,
      symbol_in  => LambdaIn(32));

  transition_123_preds(0) <= place_126_token;
  LambdaOut(33) <= transition_123_symbol_out;
  transition_123 : transition
    port map(
      preds      => transition_123_preds,
      symbol_out => transition_123_symbol_out,
      symbol_in  => true);

  transition_124_preds(0) <= place_127_token;
  transition_124 : transition
    port map(
      preds      => transition_124_preds,
      symbol_out => transition_124_symbol_out,
      symbol_in  => LambdaIn(33));

  transition_128_preds(0) <= place_1549_token;
  LambdaOut(34) <= transition_128_symbol_out;
  transition_128 : transition
    port map(
      preds      => transition_128_preds,
      symbol_out => transition_128_symbol_out,
      symbol_in  => true);

  transition_129_preds(0) <= place_132_token;
  transition_129 : transition
    port map(
      preds      => transition_129_preds,
      symbol_out => transition_129_symbol_out,
      symbol_in  => LambdaIn(34));

  transition_130_preds(0) <= place_133_token;
  LambdaOut(35) <= transition_130_symbol_out;
  transition_130 : transition
    port map(
      preds      => transition_130_preds,
      symbol_out => transition_130_symbol_out,
      symbol_in  => true);

  transition_131_preds(0) <= place_134_token;
  transition_131 : transition
    port map(
      preds      => transition_131_preds,
      symbol_out => transition_131_symbol_out,
      symbol_in  => LambdaIn(35));

  transition_135_preds(0) <= place_1550_token;
  LambdaOut(36) <= transition_135_symbol_out;
  transition_135 : transition
    port map(
      preds      => transition_135_preds,
      symbol_out => transition_135_symbol_out,
      symbol_in  => true);

  transition_136_preds(0) <= place_139_token;
  transition_136 : transition
    port map(
      preds      => transition_136_preds,
      symbol_out => transition_136_symbol_out,
      symbol_in  => LambdaIn(36));

  transition_137_preds(0) <= place_140_token;
  LambdaOut(37) <= transition_137_symbol_out;
  transition_137 : transition
    port map(
      preds      => transition_137_preds,
      symbol_out => transition_137_symbol_out,
      symbol_in  => true);

  transition_138_preds(0) <= place_141_token;
  transition_138 : transition
    port map(
      preds      => transition_138_preds,
      symbol_out => transition_138_symbol_out,
      symbol_in  => LambdaIn(37));

  transition_142_preds(0) <= place_1545_token;
  transition_142_preds(1) <= place_1547_token;
  transition_142 : transition
    port map(
      preds      => transition_142_preds,
      symbol_out => transition_142_symbol_out,
      symbol_in  => true);

  transition_143_preds(0) <= place_1553_token;
  LambdaOut(38) <= transition_143_symbol_out;
  transition_143 : transition
    port map(
      preds      => transition_143_preds,
      symbol_out => transition_143_symbol_out,
      symbol_in  => true);

  transition_144_preds(0) <= place_147_token;
  transition_144 : transition
    port map(
      preds      => transition_144_preds,
      symbol_out => transition_144_symbol_out,
      symbol_in  => LambdaIn(38));

  transition_145_preds(0) <= place_148_token;
  LambdaOut(39) <= transition_145_symbol_out;
  transition_145 : transition
    port map(
      preds      => transition_145_preds,
      symbol_out => transition_145_symbol_out,
      symbol_in  => true);

  transition_146_preds(0) <= place_149_token;
  transition_146 : transition
    port map(
      preds      => transition_146_preds,
      symbol_out => transition_146_symbol_out,
      symbol_in  => LambdaIn(39));

  transition_150_preds(0) <= place_1207_token;
  LambdaOut(40) <= transition_150_symbol_out;
  transition_150 : transition
    port map(
      preds      => transition_150_preds,
      symbol_out => transition_150_symbol_out,
      symbol_in  => true);

  transition_151_preds(0) <= place_154_token;
  transition_151 : transition
    port map(
      preds      => transition_151_preds,
      symbol_out => transition_151_symbol_out,
      symbol_in  => LambdaIn(40));

  transition_152_preds(0) <= place_155_token;
  LambdaOut(41) <= transition_152_symbol_out;
  transition_152 : transition
    port map(
      preds      => transition_152_preds,
      symbol_out => transition_152_symbol_out,
      symbol_in  => true);

  transition_153_preds(0) <= place_156_token;
  transition_153 : transition
    port map(
      preds      => transition_153_preds,
      symbol_out => transition_153_symbol_out,
      symbol_in  => LambdaIn(41));

  transition_157_preds(0) <= place_1551_token;
  transition_157_preds(1) <= place_1552_token;
  transition_157 : transition
    port map(
      preds      => transition_157_preds,
      symbol_out => transition_157_symbol_out,
      symbol_in  => true);

  transition_158_preds(0) <= place_1208_token;
  LambdaOut(42) <= transition_158_symbol_out;
  transition_158 : transition
    port map(
      preds      => transition_158_preds,
      symbol_out => transition_158_symbol_out,
      symbol_in  => true);

  transition_159_preds(0) <= place_162_token;
  transition_159 : transition
    port map(
      preds      => transition_159_preds,
      symbol_out => transition_159_symbol_out,
      symbol_in  => LambdaIn(42));

  transition_160_preds(0) <= place_163_token;
  LambdaOut(43) <= transition_160_symbol_out;
  transition_160 : transition
    port map(
      preds      => transition_160_preds,
      symbol_out => transition_160_symbol_out,
      symbol_in  => true);

  transition_161_preds(0) <= place_164_token;
  transition_161 : transition
    port map(
      preds      => transition_161_preds,
      symbol_out => transition_161_symbol_out,
      symbol_in  => LambdaIn(43));

  transition_166_preds(0) <= place_165_token;
  transition_166 : transition
    port map(
      preds      => transition_166_preds,
      symbol_out => transition_166_symbol_out,
      symbol_in  => LambdaIn(44));

  transition_167_preds(0) <= place_1210_token;
  LambdaOut(44) <= transition_167_symbol_out;
  transition_167 : transition
    port map(
      preds      => transition_167_preds,
      symbol_out => transition_167_symbol_out,
      symbol_in  => true);

  transition_168_preds(0) <= place_1209_token;
  transition_168_preds(1) <= place_1212_token;
  transition_168 : transition
    port map(
      preds      => transition_168_preds,
      symbol_out => transition_168_symbol_out,
      symbol_in  => true);

  transition_169_preds(0) <= place_1211_token;
  transition_169 : transition
    port map(
      preds      => transition_169_preds,
      symbol_out => transition_169_symbol_out,
      symbol_in  => true);

  transition_170_preds(0) <= place_1214_token;
  LambdaOut(45) <= transition_170_symbol_out;
  transition_170 : transition
    port map(
      preds      => transition_170_preds,
      symbol_out => transition_170_symbol_out,
      symbol_in  => true);

  transition_171_preds(0) <= place_174_token;
  transition_171 : transition
    port map(
      preds      => transition_171_preds,
      symbol_out => transition_171_symbol_out,
      symbol_in  => LambdaIn(45));

  transition_172_preds(0) <= place_175_token;
  LambdaOut(46) <= transition_172_symbol_out;
  transition_172 : transition
    port map(
      preds      => transition_172_preds,
      symbol_out => transition_172_symbol_out,
      symbol_in  => true);

  transition_173_preds(0) <= place_176_token;
  transition_173 : transition
    port map(
      preds      => transition_173_preds,
      symbol_out => transition_173_symbol_out,
      symbol_in  => LambdaIn(46));

  transition_177_preds(0) <= place_1216_token;
  LambdaOut(47) <= transition_177_symbol_out;
  transition_177 : transition
    port map(
      preds      => transition_177_preds,
      symbol_out => transition_177_symbol_out,
      symbol_in  => true);

  transition_178_preds(0) <= place_181_token;
  transition_178 : transition
    port map(
      preds      => transition_178_preds,
      symbol_out => transition_178_symbol_out,
      symbol_in  => LambdaIn(47));

  transition_179_preds(0) <= place_182_token;
  LambdaOut(48) <= transition_179_symbol_out;
  transition_179 : transition
    port map(
      preds      => transition_179_preds,
      symbol_out => transition_179_symbol_out,
      symbol_in  => true);

  transition_180_preds(0) <= place_183_token;
  transition_180 : transition
    port map(
      preds      => transition_180_preds,
      symbol_out => transition_180_symbol_out,
      symbol_in  => LambdaIn(48));

  transition_184_preds(0) <= place_1217_token;
  LambdaOut(49) <= transition_184_symbol_out;
  transition_184 : transition
    port map(
      preds      => transition_184_preds,
      symbol_out => transition_184_symbol_out,
      symbol_in  => true);

  transition_185_preds(0) <= place_188_token;
  transition_185 : transition
    port map(
      preds      => transition_185_preds,
      symbol_out => transition_185_symbol_out,
      symbol_in  => LambdaIn(49));

  transition_186_preds(0) <= place_189_token;
  LambdaOut(50) <= transition_186_symbol_out;
  transition_186 : transition
    port map(
      preds      => transition_186_preds,
      symbol_out => transition_186_symbol_out,
      symbol_in  => true);

  transition_187_preds(0) <= place_190_token;
  transition_187 : transition
    port map(
      preds      => transition_187_preds,
      symbol_out => transition_187_symbol_out,
      symbol_in  => LambdaIn(50));

  transition_191_preds(0) <= place_1213_token;
  transition_191_preds(1) <= place_1215_token;
  transition_191 : transition
    port map(
      preds      => transition_191_preds,
      symbol_out => transition_191_symbol_out,
      symbol_in  => true);

  transition_192_preds(0) <= place_1221_token;
  LambdaOut(51) <= transition_192_symbol_out;
  transition_192 : transition
    port map(
      preds      => transition_192_preds,
      symbol_out => transition_192_symbol_out,
      symbol_in  => true);

  transition_193_preds(0) <= place_196_token;
  transition_193 : transition
    port map(
      preds      => transition_193_preds,
      symbol_out => transition_193_symbol_out,
      symbol_in  => LambdaIn(51));

  transition_194_preds(0) <= place_197_token;
  LambdaOut(52) <= transition_194_symbol_out;
  transition_194 : transition
    port map(
      preds      => transition_194_preds,
      symbol_out => transition_194_symbol_out,
      symbol_in  => true);

  transition_195_preds(0) <= place_198_token;
  transition_195 : transition
    port map(
      preds      => transition_195_preds,
      symbol_out => transition_195_symbol_out,
      symbol_in  => LambdaIn(52));

  transition_199_preds(0) <= place_1222_token;
  LambdaOut(53) <= transition_199_symbol_out;
  transition_199 : transition
    port map(
      preds      => transition_199_preds,
      symbol_out => transition_199_symbol_out,
      symbol_in  => true);

  transition_200_preds(0) <= place_203_token;
  transition_200 : transition
    port map(
      preds      => transition_200_preds,
      symbol_out => transition_200_symbol_out,
      symbol_in  => LambdaIn(53));

  transition_201_preds(0) <= place_204_token;
  LambdaOut(54) <= transition_201_symbol_out;
  transition_201 : transition
    port map(
      preds      => transition_201_preds,
      symbol_out => transition_201_symbol_out,
      symbol_in  => true);

  transition_202_preds(0) <= place_205_token;
  transition_202 : transition
    port map(
      preds      => transition_202_preds,
      symbol_out => transition_202_symbol_out,
      symbol_in  => LambdaIn(54));

  transition_206_preds(0) <= place_1218_token;
  transition_206_preds(1) <= place_1219_token;
  transition_206 : transition
    port map(
      preds      => transition_206_preds,
      symbol_out => transition_206_symbol_out,
      symbol_in  => true);

  transition_207_preds(0) <= place_1223_token;
  LambdaOut(55) <= transition_207_symbol_out;
  transition_207 : transition
    port map(
      preds      => transition_207_preds,
      symbol_out => transition_207_symbol_out,
      symbol_in  => true);

  transition_208_preds(0) <= place_211_token;
  transition_208 : transition
    port map(
      preds      => transition_208_preds,
      symbol_out => transition_208_symbol_out,
      symbol_in  => LambdaIn(55));

  transition_209_preds(0) <= place_212_token;
  LambdaOut(56) <= transition_209_symbol_out;
  transition_209 : transition
    port map(
      preds      => transition_209_preds,
      symbol_out => transition_209_symbol_out,
      symbol_in  => true);

  transition_210_preds(0) <= place_213_token;
  transition_210 : transition
    port map(
      preds      => transition_210_preds,
      symbol_out => transition_210_symbol_out,
      symbol_in  => LambdaIn(56));

  transition_215_preds(0) <= place_214_token;
  transition_215 : transition
    port map(
      preds      => transition_215_preds,
      symbol_out => transition_215_symbol_out,
      symbol_in  => LambdaIn(57));

  transition_216_preds(0) <= place_1226_token;
  LambdaOut(57) <= transition_216_symbol_out;
  transition_216 : transition
    port map(
      preds      => transition_216_preds,
      symbol_out => transition_216_symbol_out,
      symbol_in  => true);

  transition_217_preds(0) <= place_1224_token;
  transition_217_preds(1) <= place_1229_token;
  transition_217 : transition
    port map(
      preds      => transition_217_preds,
      symbol_out => transition_217_symbol_out,
      symbol_in  => true);

  transition_219_preds(0) <= place_218_token;
  transition_219 : transition
    port map(
      preds      => transition_219_preds,
      symbol_out => transition_219_symbol_out,
      symbol_in  => LambdaIn(58));

  transition_220_preds(0) <= place_1227_token;
  LambdaOut(58) <= transition_220_symbol_out;
  transition_220 : transition
    port map(
      preds      => transition_220_preds,
      symbol_out => transition_220_symbol_out,
      symbol_in  => true);

  transition_221_preds(0) <= place_1228_token;
  transition_221 : transition
    port map(
      preds      => transition_221_preds,
      symbol_out => transition_221_symbol_out,
      symbol_in  => true);

  transition_222_preds(0) <= place_1232_token;
  LambdaOut(59) <= transition_222_symbol_out;
  transition_222 : transition
    port map(
      preds      => transition_222_preds,
      symbol_out => transition_222_symbol_out,
      symbol_in  => true);

  transition_223_preds(0) <= place_226_token;
  transition_223 : transition
    port map(
      preds      => transition_223_preds,
      symbol_out => transition_223_symbol_out,
      symbol_in  => LambdaIn(59));

  transition_224_preds(0) <= place_227_token;
  LambdaOut(60) <= transition_224_symbol_out;
  transition_224 : transition
    port map(
      preds      => transition_224_preds,
      symbol_out => transition_224_symbol_out,
      symbol_in  => true);

  transition_225_preds(0) <= place_228_token;
  transition_225 : transition
    port map(
      preds      => transition_225_preds,
      symbol_out => transition_225_symbol_out,
      symbol_in  => LambdaIn(60));

  transition_229_preds(0) <= place_1234_token;
  LambdaOut(61) <= transition_229_symbol_out;
  transition_229 : transition
    port map(
      preds      => transition_229_preds,
      symbol_out => transition_229_symbol_out,
      symbol_in  => true);

  transition_230_preds(0) <= place_233_token;
  transition_230 : transition
    port map(
      preds      => transition_230_preds,
      symbol_out => transition_230_symbol_out,
      symbol_in  => LambdaIn(61));

  transition_231_preds(0) <= place_234_token;
  LambdaOut(62) <= transition_231_symbol_out;
  transition_231 : transition
    port map(
      preds      => transition_231_preds,
      symbol_out => transition_231_symbol_out,
      symbol_in  => true);

  transition_232_preds(0) <= place_235_token;
  transition_232 : transition
    port map(
      preds      => transition_232_preds,
      symbol_out => transition_232_symbol_out,
      symbol_in  => LambdaIn(62));

  transition_236_preds(0) <= place_1235_token;
  LambdaOut(63) <= transition_236_symbol_out;
  transition_236 : transition
    port map(
      preds      => transition_236_preds,
      symbol_out => transition_236_symbol_out,
      symbol_in  => true);

  transition_237_preds(0) <= place_240_token;
  transition_237 : transition
    port map(
      preds      => transition_237_preds,
      symbol_out => transition_237_symbol_out,
      symbol_in  => LambdaIn(63));

  transition_238_preds(0) <= place_241_token;
  LambdaOut(64) <= transition_238_symbol_out;
  transition_238 : transition
    port map(
      preds      => transition_238_preds,
      symbol_out => transition_238_symbol_out,
      symbol_in  => true);

  transition_239_preds(0) <= place_242_token;
  transition_239 : transition
    port map(
      preds      => transition_239_preds,
      symbol_out => transition_239_symbol_out,
      symbol_in  => LambdaIn(64));

  transition_243_preds(0) <= place_1230_token;
  transition_243_preds(1) <= place_1233_token;
  transition_243 : transition
    port map(
      preds      => transition_243_preds,
      symbol_out => transition_243_symbol_out,
      symbol_in  => true);

  transition_244_preds(0) <= place_1238_token;
  LambdaOut(65) <= transition_244_symbol_out;
  transition_244 : transition
    port map(
      preds      => transition_244_preds,
      symbol_out => transition_244_symbol_out,
      symbol_in  => true);

  transition_245_preds(0) <= place_248_token;
  transition_245 : transition
    port map(
      preds      => transition_245_preds,
      symbol_out => transition_245_symbol_out,
      symbol_in  => LambdaIn(65));

  transition_246_preds(0) <= place_249_token;
  LambdaOut(66) <= transition_246_symbol_out;
  transition_246 : transition
    port map(
      preds      => transition_246_preds,
      symbol_out => transition_246_symbol_out,
      symbol_in  => true);

  transition_247_preds(0) <= place_250_token;
  transition_247 : transition
    port map(
      preds      => transition_247_preds,
      symbol_out => transition_247_symbol_out,
      symbol_in  => LambdaIn(66));

  transition_251_preds(0) <= place_1239_token;
  LambdaOut(67) <= transition_251_symbol_out;
  transition_251 : transition
    port map(
      preds      => transition_251_preds,
      symbol_out => transition_251_symbol_out,
      symbol_in  => true);

  transition_252_preds(0) <= place_255_token;
  transition_252 : transition
    port map(
      preds      => transition_252_preds,
      symbol_out => transition_252_symbol_out,
      symbol_in  => LambdaIn(67));

  transition_253_preds(0) <= place_256_token;
  LambdaOut(68) <= transition_253_symbol_out;
  transition_253 : transition
    port map(
      preds      => transition_253_preds,
      symbol_out => transition_253_symbol_out,
      symbol_in  => true);

  transition_254_preds(0) <= place_257_token;
  transition_254 : transition
    port map(
      preds      => transition_254_preds,
      symbol_out => transition_254_symbol_out,
      symbol_in  => LambdaIn(68));

  transition_258_preds(0) <= place_1236_token;
  transition_258_preds(1) <= place_1237_token;
  transition_258 : transition
    port map(
      preds      => transition_258_preds,
      symbol_out => transition_258_symbol_out,
      symbol_in  => true);

  transition_259_preds(0) <= place_1240_token;
  LambdaOut(69) <= transition_259_symbol_out;
  transition_259 : transition
    port map(
      preds      => transition_259_preds,
      symbol_out => transition_259_symbol_out,
      symbol_in  => true);

  transition_260_preds(0) <= place_263_token;
  transition_260 : transition
    port map(
      preds      => transition_260_preds,
      symbol_out => transition_260_symbol_out,
      symbol_in  => LambdaIn(69));

  transition_261_preds(0) <= place_264_token;
  LambdaOut(70) <= transition_261_symbol_out;
  transition_261 : transition
    port map(
      preds      => transition_261_preds,
      symbol_out => transition_261_symbol_out,
      symbol_in  => true);

  transition_262_preds(0) <= place_265_token;
  transition_262 : transition
    port map(
      preds      => transition_262_preds,
      symbol_out => transition_262_symbol_out,
      symbol_in  => LambdaIn(70));

  transition_267_preds(0) <= place_266_token;
  transition_267 : transition
    port map(
      preds      => transition_267_preds,
      symbol_out => transition_267_symbol_out,
      symbol_in  => LambdaIn(71));

  transition_268_preds(0) <= place_1242_token;
  LambdaOut(71) <= transition_268_symbol_out;
  transition_268 : transition
    port map(
      preds      => transition_268_preds,
      symbol_out => transition_268_symbol_out,
      symbol_in  => true);

  transition_269_preds(0) <= place_1241_token;
  transition_269_preds(1) <= place_1245_token;
  transition_269 : transition
    port map(
      preds      => transition_269_preds,
      symbol_out => transition_269_symbol_out,
      symbol_in  => true);

  transition_271_preds(0) <= place_270_token;
  transition_271 : transition
    port map(
      preds      => transition_271_preds,
      symbol_out => transition_271_symbol_out,
      symbol_in  => LambdaIn(72));

  transition_272_preds(0) <= place_1243_token;
  LambdaOut(72) <= transition_272_symbol_out;
  transition_272 : transition
    port map(
      preds      => transition_272_preds,
      symbol_out => transition_272_symbol_out,
      symbol_in  => true);

  transition_273_preds(0) <= place_1244_token;
  transition_273 : transition
    port map(
      preds      => transition_273_preds,
      symbol_out => transition_273_symbol_out,
      symbol_in  => true);

  transition_274_preds(0) <= place_1246_token;
  LambdaOut(73) <= transition_274_symbol_out;
  transition_274 : transition
    port map(
      preds      => transition_274_preds,
      symbol_out => transition_274_symbol_out,
      symbol_in  => true);

  transition_275_preds(0) <= place_278_token;
  transition_275 : transition
    port map(
      preds      => transition_275_preds,
      symbol_out => transition_275_symbol_out,
      symbol_in  => LambdaIn(73));

  transition_276_preds(0) <= place_279_token;
  LambdaOut(74) <= transition_276_symbol_out;
  transition_276 : transition
    port map(
      preds      => transition_276_preds,
      symbol_out => transition_276_symbol_out,
      symbol_in  => true);

  transition_277_preds(0) <= place_280_token;
  transition_277 : transition
    port map(
      preds      => transition_277_preds,
      symbol_out => transition_277_symbol_out,
      symbol_in  => LambdaIn(74));

  transition_281_preds(0) <= place_1248_token;
  transition_281_preds(1) <= place_1249_token;
  transition_281 : transition
    port map(
      preds      => transition_281_preds,
      symbol_out => transition_281_symbol_out,
      symbol_in  => true);

  transition_282_preds(0) <= place_1247_token;
  transition_282 : transition
    port map(
      preds      => transition_282_preds,
      symbol_out => transition_282_symbol_out,
      symbol_in  => true);

  transition_283_preds(0) <= place_1251_token;
  LambdaOut(75) <= transition_283_symbol_out;
  transition_283 : transition
    port map(
      preds      => transition_283_preds,
      symbol_out => transition_283_symbol_out,
      symbol_in  => true);

  transition_284_preds(0) <= place_287_token;
  transition_284 : transition
    port map(
      preds      => transition_284_preds,
      symbol_out => transition_284_symbol_out,
      symbol_in  => LambdaIn(75));

  transition_285_preds(0) <= place_288_token;
  LambdaOut(76) <= transition_285_symbol_out;
  transition_285 : transition
    port map(
      preds      => transition_285_preds,
      symbol_out => transition_285_symbol_out,
      symbol_in  => true);

  transition_286_preds(0) <= place_289_token;
  transition_286 : transition
    port map(
      preds      => transition_286_preds,
      symbol_out => transition_286_symbol_out,
      symbol_in  => LambdaIn(76));

  transition_290_preds(0) <= place_1253_token;
  LambdaOut(77) <= transition_290_symbol_out;
  transition_290 : transition
    port map(
      preds      => transition_290_preds,
      symbol_out => transition_290_symbol_out,
      symbol_in  => true);

  transition_291_preds(0) <= place_294_token;
  transition_291 : transition
    port map(
      preds      => transition_291_preds,
      symbol_out => transition_291_symbol_out,
      symbol_in  => LambdaIn(77));

  transition_292_preds(0) <= place_295_token;
  LambdaOut(78) <= transition_292_symbol_out;
  transition_292 : transition
    port map(
      preds      => transition_292_preds,
      symbol_out => transition_292_symbol_out,
      symbol_in  => true);

  transition_293_preds(0) <= place_296_token;
  transition_293 : transition
    port map(
      preds      => transition_293_preds,
      symbol_out => transition_293_symbol_out,
      symbol_in  => LambdaIn(78));

  transition_297_preds(0) <= place_1254_token;
  LambdaOut(79) <= transition_297_symbol_out;
  transition_297 : transition
    port map(
      preds      => transition_297_preds,
      symbol_out => transition_297_symbol_out,
      symbol_in  => true);

  transition_298_preds(0) <= place_301_token;
  transition_298 : transition
    port map(
      preds      => transition_298_preds,
      symbol_out => transition_298_symbol_out,
      symbol_in  => LambdaIn(79));

  transition_299_preds(0) <= place_302_token;
  LambdaOut(80) <= transition_299_symbol_out;
  transition_299 : transition
    port map(
      preds      => transition_299_preds,
      symbol_out => transition_299_symbol_out,
      symbol_in  => true);

  transition_300_preds(0) <= place_303_token;
  transition_300 : transition
    port map(
      preds      => transition_300_preds,
      symbol_out => transition_300_symbol_out,
      symbol_in  => LambdaIn(80));

  transition_304_preds(0) <= place_1252_token;
  transition_304_preds(1) <= place_1250_token;
  transition_304 : transition
    port map(
      preds      => transition_304_preds,
      symbol_out => transition_304_symbol_out,
      symbol_in  => true);

  transition_305_preds(0) <= place_1259_token;
  LambdaOut(81) <= transition_305_symbol_out;
  transition_305 : transition
    port map(
      preds      => transition_305_preds,
      symbol_out => transition_305_symbol_out,
      symbol_in  => true);

  transition_306_preds(0) <= place_309_token;
  transition_306 : transition
    port map(
      preds      => transition_306_preds,
      symbol_out => transition_306_symbol_out,
      symbol_in  => LambdaIn(81));

  transition_307_preds(0) <= place_310_token;
  LambdaOut(82) <= transition_307_symbol_out;
  transition_307 : transition
    port map(
      preds      => transition_307_preds,
      symbol_out => transition_307_symbol_out,
      symbol_in  => true);

  transition_308_preds(0) <= place_311_token;
  transition_308 : transition
    port map(
      preds      => transition_308_preds,
      symbol_out => transition_308_symbol_out,
      symbol_in  => LambdaIn(82));

  transition_312_preds(0) <= place_1260_token;
  LambdaOut(83) <= transition_312_symbol_out;
  transition_312 : transition
    port map(
      preds      => transition_312_preds,
      symbol_out => transition_312_symbol_out,
      symbol_in  => true);

  transition_313_preds(0) <= place_316_token;
  transition_313 : transition
    port map(
      preds      => transition_313_preds,
      symbol_out => transition_313_symbol_out,
      symbol_in  => LambdaIn(83));

  transition_314_preds(0) <= place_317_token;
  LambdaOut(84) <= transition_314_symbol_out;
  transition_314 : transition
    port map(
      preds      => transition_314_preds,
      symbol_out => transition_314_symbol_out,
      symbol_in  => true);

  transition_315_preds(0) <= place_318_token;
  transition_315 : transition
    port map(
      preds      => transition_315_preds,
      symbol_out => transition_315_symbol_out,
      symbol_in  => LambdaIn(84));

  transition_319_preds(0) <= place_1255_token;
  transition_319_preds(1) <= place_1258_token;
  transition_319 : transition
    port map(
      preds      => transition_319_preds,
      symbol_out => transition_319_symbol_out,
      symbol_in  => true);

  transition_320_preds(0) <= place_1261_token;
  LambdaOut(85) <= transition_320_symbol_out;
  transition_320 : transition
    port map(
      preds      => transition_320_preds,
      symbol_out => transition_320_symbol_out,
      symbol_in  => true);

  transition_321_preds(0) <= place_324_token;
  transition_321 : transition
    port map(
      preds      => transition_321_preds,
      symbol_out => transition_321_symbol_out,
      symbol_in  => LambdaIn(85));

  transition_322_preds(0) <= place_325_token;
  LambdaOut(86) <= transition_322_symbol_out;
  transition_322 : transition
    port map(
      preds      => transition_322_preds,
      symbol_out => transition_322_symbol_out,
      symbol_in  => true);

  transition_323_preds(0) <= place_326_token;
  transition_323 : transition
    port map(
      preds      => transition_323_preds,
      symbol_out => transition_323_symbol_out,
      symbol_in  => LambdaIn(86));

  transition_328_preds(0) <= place_327_token;
  transition_328 : transition
    port map(
      preds      => transition_328_preds,
      symbol_out => transition_328_symbol_out,
      symbol_in  => LambdaIn(87));

  transition_329_preds(0) <= place_1263_token;
  LambdaOut(87) <= transition_329_symbol_out;
  transition_329 : transition
    port map(
      preds      => transition_329_preds,
      symbol_out => transition_329_symbol_out,
      symbol_in  => true);

  transition_330_preds(0) <= place_1262_token;
  transition_330_preds(1) <= place_1265_token;
  transition_330 : transition
    port map(
      preds      => transition_330_preds,
      symbol_out => transition_330_symbol_out,
      symbol_in  => true);

  transition_331_preds(0) <= place_1264_token;
  transition_331 : transition
    port map(
      preds      => transition_331_preds,
      symbol_out => transition_331_symbol_out,
      symbol_in  => true);

  transition_332_preds(0) <= place_1267_token;
  LambdaOut(88) <= transition_332_symbol_out;
  transition_332 : transition
    port map(
      preds      => transition_332_preds,
      symbol_out => transition_332_symbol_out,
      symbol_in  => true);

  transition_333_preds(0) <= place_336_token;
  transition_333 : transition
    port map(
      preds      => transition_333_preds,
      symbol_out => transition_333_symbol_out,
      symbol_in  => LambdaIn(88));

  transition_334_preds(0) <= place_337_token;
  LambdaOut(89) <= transition_334_symbol_out;
  transition_334 : transition
    port map(
      preds      => transition_334_preds,
      symbol_out => transition_334_symbol_out,
      symbol_in  => true);

  transition_335_preds(0) <= place_338_token;
  transition_335 : transition
    port map(
      preds      => transition_335_preds,
      symbol_out => transition_335_symbol_out,
      symbol_in  => LambdaIn(89));

  transition_339_preds(0) <= place_1269_token;
  LambdaOut(90) <= transition_339_symbol_out;
  transition_339 : transition
    port map(
      preds      => transition_339_preds,
      symbol_out => transition_339_symbol_out,
      symbol_in  => true);

  transition_340_preds(0) <= place_343_token;
  transition_340 : transition
    port map(
      preds      => transition_340_preds,
      symbol_out => transition_340_symbol_out,
      symbol_in  => LambdaIn(90));

  transition_341_preds(0) <= place_344_token;
  LambdaOut(91) <= transition_341_symbol_out;
  transition_341 : transition
    port map(
      preds      => transition_341_preds,
      symbol_out => transition_341_symbol_out,
      symbol_in  => true);

  transition_342_preds(0) <= place_345_token;
  transition_342 : transition
    port map(
      preds      => transition_342_preds,
      symbol_out => transition_342_symbol_out,
      symbol_in  => LambdaIn(91));

  transition_346_preds(0) <= place_1270_token;
  LambdaOut(92) <= transition_346_symbol_out;
  transition_346 : transition
    port map(
      preds      => transition_346_preds,
      symbol_out => transition_346_symbol_out,
      symbol_in  => true);

  transition_347_preds(0) <= place_350_token;
  transition_347 : transition
    port map(
      preds      => transition_347_preds,
      symbol_out => transition_347_symbol_out,
      symbol_in  => LambdaIn(92));

  transition_348_preds(0) <= place_351_token;
  LambdaOut(93) <= transition_348_symbol_out;
  transition_348 : transition
    port map(
      preds      => transition_348_preds,
      symbol_out => transition_348_symbol_out,
      symbol_in  => true);

  transition_349_preds(0) <= place_352_token;
  transition_349 : transition
    port map(
      preds      => transition_349_preds,
      symbol_out => transition_349_symbol_out,
      symbol_in  => LambdaIn(93));

  transition_353_preds(0) <= place_1266_token;
  transition_353_preds(1) <= place_1268_token;
  transition_353 : transition
    port map(
      preds      => transition_353_preds,
      symbol_out => transition_353_symbol_out,
      symbol_in  => true);

  transition_354_preds(0) <= place_1274_token;
  LambdaOut(94) <= transition_354_symbol_out;
  transition_354 : transition
    port map(
      preds      => transition_354_preds,
      symbol_out => transition_354_symbol_out,
      symbol_in  => true);

  transition_355_preds(0) <= place_358_token;
  transition_355 : transition
    port map(
      preds      => transition_355_preds,
      symbol_out => transition_355_symbol_out,
      symbol_in  => LambdaIn(94));

  transition_356_preds(0) <= place_359_token;
  LambdaOut(95) <= transition_356_symbol_out;
  transition_356 : transition
    port map(
      preds      => transition_356_preds,
      symbol_out => transition_356_symbol_out,
      symbol_in  => true);

  transition_357_preds(0) <= place_360_token;
  transition_357 : transition
    port map(
      preds      => transition_357_preds,
      symbol_out => transition_357_symbol_out,
      symbol_in  => LambdaIn(95));

  transition_361_preds(0) <= place_1275_token;
  LambdaOut(96) <= transition_361_symbol_out;
  transition_361 : transition
    port map(
      preds      => transition_361_preds,
      symbol_out => transition_361_symbol_out,
      symbol_in  => true);

  transition_362_preds(0) <= place_365_token;
  transition_362 : transition
    port map(
      preds      => transition_362_preds,
      symbol_out => transition_362_symbol_out,
      symbol_in  => LambdaIn(96));

  transition_363_preds(0) <= place_366_token;
  LambdaOut(97) <= transition_363_symbol_out;
  transition_363 : transition
    port map(
      preds      => transition_363_preds,
      symbol_out => transition_363_symbol_out,
      symbol_in  => true);

  transition_364_preds(0) <= place_367_token;
  transition_364 : transition
    port map(
      preds      => transition_364_preds,
      symbol_out => transition_364_symbol_out,
      symbol_in  => LambdaIn(97));

  transition_368_preds(0) <= place_1273_token;
  transition_368_preds(1) <= place_1271_token;
  transition_368 : transition
    port map(
      preds      => transition_368_preds,
      symbol_out => transition_368_symbol_out,
      symbol_in  => true);

  transition_369_preds(0) <= place_1276_token;
  LambdaOut(98) <= transition_369_symbol_out;
  transition_369 : transition
    port map(
      preds      => transition_369_preds,
      symbol_out => transition_369_symbol_out,
      symbol_in  => true);

  transition_370_preds(0) <= place_373_token;
  transition_370 : transition
    port map(
      preds      => transition_370_preds,
      symbol_out => transition_370_symbol_out,
      symbol_in  => LambdaIn(98));

  transition_371_preds(0) <= place_374_token;
  LambdaOut(99) <= transition_371_symbol_out;
  transition_371 : transition
    port map(
      preds      => transition_371_preds,
      symbol_out => transition_371_symbol_out,
      symbol_in  => true);

  transition_372_preds(0) <= place_375_token;
  transition_372 : transition
    port map(
      preds      => transition_372_preds,
      symbol_out => transition_372_symbol_out,
      symbol_in  => LambdaIn(99));

  transition_377_preds(0) <= place_376_token;
  transition_377 : transition
    port map(
      preds      => transition_377_preds,
      symbol_out => transition_377_symbol_out,
      symbol_in  => LambdaIn(100));

  transition_378_preds(0) <= place_1279_token;
  LambdaOut(100) <= transition_378_symbol_out;
  transition_378 : transition
    port map(
      preds      => transition_378_preds,
      symbol_out => transition_378_symbol_out,
      symbol_in  => true);

  transition_379_preds(0) <= place_1278_token;
  transition_379_preds(1) <= place_1283_token;
  transition_379 : transition
    port map(
      preds      => transition_379_preds,
      symbol_out => transition_379_symbol_out,
      symbol_in  => true);

  transition_381_preds(0) <= place_380_token;
  transition_381 : transition
    port map(
      preds      => transition_381_preds,
      symbol_out => transition_381_symbol_out,
      symbol_in  => LambdaIn(101));

  transition_382_preds(0) <= place_1280_token;
  LambdaOut(101) <= transition_382_symbol_out;
  transition_382 : transition
    port map(
      preds      => transition_382_preds,
      symbol_out => transition_382_symbol_out,
      symbol_in  => true);

  transition_383_preds(0) <= place_1281_token;
  transition_383 : transition
    port map(
      preds      => transition_383_preds,
      symbol_out => transition_383_symbol_out,
      symbol_in  => true);

  transition_384_preds(0) <= place_1285_token;
  LambdaOut(102) <= transition_384_symbol_out;
  transition_384 : transition
    port map(
      preds      => transition_384_preds,
      symbol_out => transition_384_symbol_out,
      symbol_in  => true);

  transition_385_preds(0) <= place_388_token;
  transition_385 : transition
    port map(
      preds      => transition_385_preds,
      symbol_out => transition_385_symbol_out,
      symbol_in  => LambdaIn(102));

  transition_386_preds(0) <= place_389_token;
  LambdaOut(103) <= transition_386_symbol_out;
  transition_386 : transition
    port map(
      preds      => transition_386_preds,
      symbol_out => transition_386_symbol_out,
      symbol_in  => true);

  transition_387_preds(0) <= place_390_token;
  transition_387 : transition
    port map(
      preds      => transition_387_preds,
      symbol_out => transition_387_symbol_out,
      symbol_in  => LambdaIn(103));

  transition_391_preds(0) <= place_1287_token;
  LambdaOut(104) <= transition_391_symbol_out;
  transition_391 : transition
    port map(
      preds      => transition_391_preds,
      symbol_out => transition_391_symbol_out,
      symbol_in  => true);

  transition_392_preds(0) <= place_395_token;
  transition_392 : transition
    port map(
      preds      => transition_392_preds,
      symbol_out => transition_392_symbol_out,
      symbol_in  => LambdaIn(104));

  transition_393_preds(0) <= place_396_token;
  LambdaOut(105) <= transition_393_symbol_out;
  transition_393 : transition
    port map(
      preds      => transition_393_preds,
      symbol_out => transition_393_symbol_out,
      symbol_in  => true);

  transition_394_preds(0) <= place_397_token;
  transition_394 : transition
    port map(
      preds      => transition_394_preds,
      symbol_out => transition_394_symbol_out,
      symbol_in  => LambdaIn(105));

  transition_398_preds(0) <= place_1288_token;
  LambdaOut(106) <= transition_398_symbol_out;
  transition_398 : transition
    port map(
      preds      => transition_398_preds,
      symbol_out => transition_398_symbol_out,
      symbol_in  => true);

  transition_399_preds(0) <= place_402_token;
  transition_399 : transition
    port map(
      preds      => transition_399_preds,
      symbol_out => transition_399_symbol_out,
      symbol_in  => LambdaIn(106));

  transition_400_preds(0) <= place_403_token;
  LambdaOut(107) <= transition_400_symbol_out;
  transition_400 : transition
    port map(
      preds      => transition_400_preds,
      symbol_out => transition_400_symbol_out,
      symbol_in  => true);

  transition_401_preds(0) <= place_404_token;
  transition_401 : transition
    port map(
      preds      => transition_401_preds,
      symbol_out => transition_401_symbol_out,
      symbol_in  => LambdaIn(107));

  transition_405_preds(0) <= place_1286_token;
  transition_405_preds(1) <= place_1284_token;
  transition_405 : transition
    port map(
      preds      => transition_405_preds,
      symbol_out => transition_405_symbol_out,
      symbol_in  => true);

  transition_406_preds(0) <= place_1291_token;
  LambdaOut(108) <= transition_406_symbol_out;
  transition_406 : transition
    port map(
      preds      => transition_406_preds,
      symbol_out => transition_406_symbol_out,
      symbol_in  => true);

  transition_407_preds(0) <= place_410_token;
  transition_407 : transition
    port map(
      preds      => transition_407_preds,
      symbol_out => transition_407_symbol_out,
      symbol_in  => LambdaIn(108));

  transition_408_preds(0) <= place_411_token;
  LambdaOut(109) <= transition_408_symbol_out;
  transition_408 : transition
    port map(
      preds      => transition_408_preds,
      symbol_out => transition_408_symbol_out,
      symbol_in  => true);

  transition_409_preds(0) <= place_412_token;
  transition_409 : transition
    port map(
      preds      => transition_409_preds,
      symbol_out => transition_409_symbol_out,
      symbol_in  => LambdaIn(109));

  transition_413_preds(0) <= place_1292_token;
  LambdaOut(110) <= transition_413_symbol_out;
  transition_413 : transition
    port map(
      preds      => transition_413_preds,
      symbol_out => transition_413_symbol_out,
      symbol_in  => true);

  transition_414_preds(0) <= place_417_token;
  transition_414 : transition
    port map(
      preds      => transition_414_preds,
      symbol_out => transition_414_symbol_out,
      symbol_in  => LambdaIn(110));

  transition_415_preds(0) <= place_418_token;
  LambdaOut(111) <= transition_415_symbol_out;
  transition_415 : transition
    port map(
      preds      => transition_415_preds,
      symbol_out => transition_415_symbol_out,
      symbol_in  => true);

  transition_416_preds(0) <= place_419_token;
  transition_416 : transition
    port map(
      preds      => transition_416_preds,
      symbol_out => transition_416_symbol_out,
      symbol_in  => LambdaIn(111));

  transition_420_preds(0) <= place_1289_token;
  transition_420_preds(1) <= place_1290_token;
  transition_420 : transition
    port map(
      preds      => transition_420_preds,
      symbol_out => transition_420_symbol_out,
      symbol_in  => true);

  transition_421_preds(0) <= place_1293_token;
  LambdaOut(112) <= transition_421_symbol_out;
  transition_421 : transition
    port map(
      preds      => transition_421_preds,
      symbol_out => transition_421_symbol_out,
      symbol_in  => true);

  transition_422_preds(0) <= place_425_token;
  transition_422 : transition
    port map(
      preds      => transition_422_preds,
      symbol_out => transition_422_symbol_out,
      symbol_in  => LambdaIn(112));

  transition_423_preds(0) <= place_426_token;
  LambdaOut(113) <= transition_423_symbol_out;
  transition_423 : transition
    port map(
      preds      => transition_423_preds,
      symbol_out => transition_423_symbol_out,
      symbol_in  => true);

  transition_424_preds(0) <= place_427_token;
  transition_424 : transition
    port map(
      preds      => transition_424_preds,
      symbol_out => transition_424_symbol_out,
      symbol_in  => LambdaIn(113));

  transition_429_preds(0) <= place_428_token;
  transition_429 : transition
    port map(
      preds      => transition_429_preds,
      symbol_out => transition_429_symbol_out,
      symbol_in  => LambdaIn(114));

  transition_430_preds(0) <= place_1295_token;
  LambdaOut(114) <= transition_430_symbol_out;
  transition_430 : transition
    port map(
      preds      => transition_430_preds,
      symbol_out => transition_430_symbol_out,
      symbol_in  => true);

  transition_431_preds(0) <= place_1298_token;
  transition_431_preds(1) <= place_1294_token;
  transition_431 : transition
    port map(
      preds      => transition_431_preds,
      symbol_out => transition_431_symbol_out,
      symbol_in  => true);

  transition_433_preds(0) <= place_432_token;
  transition_433 : transition
    port map(
      preds      => transition_433_preds,
      symbol_out => transition_433_symbol_out,
      symbol_in  => LambdaIn(115));

  transition_434_preds(0) <= place_1296_token;
  LambdaOut(115) <= transition_434_symbol_out;
  transition_434 : transition
    port map(
      preds      => transition_434_preds,
      symbol_out => transition_434_symbol_out,
      symbol_in  => true);

  transition_435_preds(0) <= place_1297_token;
  transition_435 : transition
    port map(
      preds      => transition_435_preds,
      symbol_out => transition_435_symbol_out,
      symbol_in  => true);

  transition_436_preds(0) <= place_1299_token;
  LambdaOut(116) <= transition_436_symbol_out;
  transition_436 : transition
    port map(
      preds      => transition_436_preds,
      symbol_out => transition_436_symbol_out,
      symbol_in  => true);

  transition_437_preds(0) <= place_440_token;
  transition_437 : transition
    port map(
      preds      => transition_437_preds,
      symbol_out => transition_437_symbol_out,
      symbol_in  => LambdaIn(116));

  transition_438_preds(0) <= place_441_token;
  LambdaOut(117) <= transition_438_symbol_out;
  transition_438 : transition
    port map(
      preds      => transition_438_preds,
      symbol_out => transition_438_symbol_out,
      symbol_in  => true);

  transition_439_preds(0) <= place_442_token;
  transition_439 : transition
    port map(
      preds      => transition_439_preds,
      symbol_out => transition_439_symbol_out,
      symbol_in  => LambdaIn(117));

  transition_443_preds(0) <= place_1301_token;
  transition_443_preds(1) <= place_1302_token;
  transition_443 : transition
    port map(
      preds      => transition_443_preds,
      symbol_out => transition_443_symbol_out,
      symbol_in  => true);

  transition_444_preds(0) <= place_1300_token;
  transition_444 : transition
    port map(
      preds      => transition_444_preds,
      symbol_out => transition_444_symbol_out,
      symbol_in  => true);

  transition_445_preds(0) <= place_1304_token;
  LambdaOut(118) <= transition_445_symbol_out;
  transition_445 : transition
    port map(
      preds      => transition_445_preds,
      symbol_out => transition_445_symbol_out,
      symbol_in  => true);

  transition_446_preds(0) <= place_449_token;
  transition_446 : transition
    port map(
      preds      => transition_446_preds,
      symbol_out => transition_446_symbol_out,
      symbol_in  => LambdaIn(118));

  transition_447_preds(0) <= place_450_token;
  LambdaOut(119) <= transition_447_symbol_out;
  transition_447 : transition
    port map(
      preds      => transition_447_preds,
      symbol_out => transition_447_symbol_out,
      symbol_in  => true);

  transition_448_preds(0) <= place_451_token;
  transition_448 : transition
    port map(
      preds      => transition_448_preds,
      symbol_out => transition_448_symbol_out,
      symbol_in  => LambdaIn(119));

  transition_452_preds(0) <= place_1306_token;
  LambdaOut(120) <= transition_452_symbol_out;
  transition_452 : transition
    port map(
      preds      => transition_452_preds,
      symbol_out => transition_452_symbol_out,
      symbol_in  => true);

  transition_453_preds(0) <= place_456_token;
  transition_453 : transition
    port map(
      preds      => transition_453_preds,
      symbol_out => transition_453_symbol_out,
      symbol_in  => LambdaIn(120));

  transition_454_preds(0) <= place_457_token;
  LambdaOut(121) <= transition_454_symbol_out;
  transition_454 : transition
    port map(
      preds      => transition_454_preds,
      symbol_out => transition_454_symbol_out,
      symbol_in  => true);

  transition_455_preds(0) <= place_458_token;
  transition_455 : transition
    port map(
      preds      => transition_455_preds,
      symbol_out => transition_455_symbol_out,
      symbol_in  => LambdaIn(121));

  transition_459_preds(0) <= place_1307_token;
  LambdaOut(122) <= transition_459_symbol_out;
  transition_459 : transition
    port map(
      preds      => transition_459_preds,
      symbol_out => transition_459_symbol_out,
      symbol_in  => true);

  transition_460_preds(0) <= place_463_token;
  transition_460 : transition
    port map(
      preds      => transition_460_preds,
      symbol_out => transition_460_symbol_out,
      symbol_in  => LambdaIn(122));

  transition_461_preds(0) <= place_464_token;
  LambdaOut(123) <= transition_461_symbol_out;
  transition_461 : transition
    port map(
      preds      => transition_461_preds,
      symbol_out => transition_461_symbol_out,
      symbol_in  => true);

  transition_462_preds(0) <= place_465_token;
  transition_462 : transition
    port map(
      preds      => transition_462_preds,
      symbol_out => transition_462_symbol_out,
      symbol_in  => LambdaIn(123));

  transition_466_preds(0) <= place_1305_token;
  transition_466_preds(1) <= place_1303_token;
  transition_466 : transition
    port map(
      preds      => transition_466_preds,
      symbol_out => transition_466_symbol_out,
      symbol_in  => true);

  transition_467_preds(0) <= place_1311_token;
  LambdaOut(124) <= transition_467_symbol_out;
  transition_467 : transition
    port map(
      preds      => transition_467_preds,
      symbol_out => transition_467_symbol_out,
      symbol_in  => true);

  transition_468_preds(0) <= place_471_token;
  transition_468 : transition
    port map(
      preds      => transition_468_preds,
      symbol_out => transition_468_symbol_out,
      symbol_in  => LambdaIn(124));

  transition_469_preds(0) <= place_472_token;
  LambdaOut(125) <= transition_469_symbol_out;
  transition_469 : transition
    port map(
      preds      => transition_469_preds,
      symbol_out => transition_469_symbol_out,
      symbol_in  => true);

  transition_470_preds(0) <= place_473_token;
  transition_470 : transition
    port map(
      preds      => transition_470_preds,
      symbol_out => transition_470_symbol_out,
      symbol_in  => LambdaIn(125));

  transition_474_preds(0) <= place_1312_token;
  LambdaOut(126) <= transition_474_symbol_out;
  transition_474 : transition
    port map(
      preds      => transition_474_preds,
      symbol_out => transition_474_symbol_out,
      symbol_in  => true);

  transition_475_preds(0) <= place_478_token;
  transition_475 : transition
    port map(
      preds      => transition_475_preds,
      symbol_out => transition_475_symbol_out,
      symbol_in  => LambdaIn(126));

  transition_476_preds(0) <= place_479_token;
  LambdaOut(127) <= transition_476_symbol_out;
  transition_476 : transition
    port map(
      preds      => transition_476_preds,
      symbol_out => transition_476_symbol_out,
      symbol_in  => true);

  transition_477_preds(0) <= place_480_token;
  transition_477 : transition
    port map(
      preds      => transition_477_preds,
      symbol_out => transition_477_symbol_out,
      symbol_in  => LambdaIn(127));

  transition_481_preds(0) <= place_1309_token;
  transition_481_preds(1) <= place_1310_token;
  transition_481 : transition
    port map(
      preds      => transition_481_preds,
      symbol_out => transition_481_symbol_out,
      symbol_in  => true);

  transition_482_preds(0) <= place_1313_token;
  LambdaOut(128) <= transition_482_symbol_out;
  transition_482 : transition
    port map(
      preds      => transition_482_preds,
      symbol_out => transition_482_symbol_out,
      symbol_in  => true);

  transition_483_preds(0) <= place_486_token;
  transition_483 : transition
    port map(
      preds      => transition_483_preds,
      symbol_out => transition_483_symbol_out,
      symbol_in  => LambdaIn(128));

  transition_484_preds(0) <= place_487_token;
  LambdaOut(129) <= transition_484_symbol_out;
  transition_484 : transition
    port map(
      preds      => transition_484_preds,
      symbol_out => transition_484_symbol_out,
      symbol_in  => true);

  transition_485_preds(0) <= place_488_token;
  transition_485 : transition
    port map(
      preds      => transition_485_preds,
      symbol_out => transition_485_symbol_out,
      symbol_in  => LambdaIn(129));

  transition_490_preds(0) <= place_489_token;
  transition_490 : transition
    port map(
      preds      => transition_490_preds,
      symbol_out => transition_490_symbol_out,
      symbol_in  => LambdaIn(130));

  transition_491_preds(0) <= place_1315_token;
  LambdaOut(130) <= transition_491_symbol_out;
  transition_491 : transition
    port map(
      preds      => transition_491_preds,
      symbol_out => transition_491_symbol_out,
      symbol_in  => true);

  transition_492_preds(0) <= place_1314_token;
  transition_492_preds(1) <= place_1317_token;
  transition_492 : transition
    port map(
      preds      => transition_492_preds,
      symbol_out => transition_492_symbol_out,
      symbol_in  => true);

  transition_493_preds(0) <= place_1318_token;
  LambdaOut(131) <= transition_493_symbol_out;
  transition_493 : transition
    port map(
      preds      => transition_493_preds,
      symbol_out => transition_493_symbol_out,
      symbol_in  => true);

  transition_494_preds(0) <= place_497_token;
  transition_494 : transition
    port map(
      preds      => transition_494_preds,
      symbol_out => transition_494_symbol_out,
      symbol_in  => LambdaIn(131));

  transition_495_preds(0) <= place_498_token;
  LambdaOut(132) <= transition_495_symbol_out;
  transition_495 : transition
    port map(
      preds      => transition_495_preds,
      symbol_out => transition_495_symbol_out,
      symbol_in  => true);

  transition_496_preds(0) <= place_499_token;
  transition_496 : transition
    port map(
      preds      => transition_496_preds,
      symbol_out => transition_496_symbol_out,
      symbol_in  => LambdaIn(132));

  transition_500_preds(0) <= place_1320_token;
  transition_500_preds(1) <= place_1321_token;
  transition_500 : transition
    port map(
      preds      => transition_500_preds,
      symbol_out => transition_500_symbol_out,
      symbol_in  => true);

  transition_501_preds(0) <= place_1319_token;
  LambdaOut(133) <= transition_501_symbol_out;
  transition_501 : transition
    port map(
      preds      => transition_501_preds,
      symbol_out => transition_501_symbol_out,
      symbol_in  => true);

  transition_502_preds(0) <= place_505_token;
  transition_502 : transition
    port map(
      preds      => transition_502_preds,
      symbol_out => transition_502_symbol_out,
      symbol_in  => LambdaIn(133));

  transition_503_preds(0) <= place_506_token;
  LambdaOut(134) <= transition_503_symbol_out;
  transition_503 : transition
    port map(
      preds      => transition_503_preds,
      symbol_out => transition_503_symbol_out,
      symbol_in  => true);

  transition_504_preds(0) <= place_507_token;
  transition_504 : transition
    port map(
      preds      => transition_504_preds,
      symbol_out => transition_504_symbol_out,
      symbol_in  => LambdaIn(134));

  transition_508_preds(0) <= place_1325_token;
  LambdaOut(135) <= transition_508_symbol_out;
  transition_508 : transition
    port map(
      preds      => transition_508_preds,
      symbol_out => transition_508_symbol_out,
      symbol_in  => true);

  transition_509_preds(0) <= place_512_token;
  transition_509 : transition
    port map(
      preds      => transition_509_preds,
      symbol_out => transition_509_symbol_out,
      symbol_in  => LambdaIn(135));

  transition_510_preds(0) <= place_513_token;
  LambdaOut(136) <= transition_510_symbol_out;
  transition_510 : transition
    port map(
      preds      => transition_510_preds,
      symbol_out => transition_510_symbol_out,
      symbol_in  => true);

  transition_511_preds(0) <= place_514_token;
  transition_511 : transition
    port map(
      preds      => transition_511_preds,
      symbol_out => transition_511_symbol_out,
      symbol_in  => LambdaIn(136));

  transition_515_preds(0) <= place_1327_token;
  LambdaOut(137) <= transition_515_symbol_out;
  transition_515 : transition
    port map(
      preds      => transition_515_preds,
      symbol_out => transition_515_symbol_out,
      symbol_in  => true);

  transition_516_preds(0) <= place_519_token;
  transition_516 : transition
    port map(
      preds      => transition_516_preds,
      symbol_out => transition_516_symbol_out,
      symbol_in  => LambdaIn(137));

  transition_517_preds(0) <= place_520_token;
  LambdaOut(138) <= transition_517_symbol_out;
  transition_517 : transition
    port map(
      preds      => transition_517_preds,
      symbol_out => transition_517_symbol_out,
      symbol_in  => true);

  transition_518_preds(0) <= place_521_token;
  transition_518 : transition
    port map(
      preds      => transition_518_preds,
      symbol_out => transition_518_symbol_out,
      symbol_in  => LambdaIn(138));

  transition_522_preds(0) <= place_1328_token;
  LambdaOut(139) <= transition_522_symbol_out;
  transition_522 : transition
    port map(
      preds      => transition_522_preds,
      symbol_out => transition_522_symbol_out,
      symbol_in  => true);

  transition_523_preds(0) <= place_526_token;
  transition_523 : transition
    port map(
      preds      => transition_523_preds,
      symbol_out => transition_523_symbol_out,
      symbol_in  => LambdaIn(139));

  transition_524_preds(0) <= place_527_token;
  LambdaOut(140) <= transition_524_symbol_out;
  transition_524 : transition
    port map(
      preds      => transition_524_preds,
      symbol_out => transition_524_symbol_out,
      symbol_in  => true);

  transition_525_preds(0) <= place_528_token;
  transition_525 : transition
    port map(
      preds      => transition_525_preds,
      symbol_out => transition_525_symbol_out,
      symbol_in  => LambdaIn(140));

  transition_529_preds(0) <= place_1324_token;
  transition_529_preds(1) <= place_1326_token;
  transition_529 : transition
    port map(
      preds      => transition_529_preds,
      symbol_out => transition_529_symbol_out,
      symbol_in  => true);

  transition_530_preds(0) <= place_1332_token;
  LambdaOut(141) <= transition_530_symbol_out;
  transition_530 : transition
    port map(
      preds      => transition_530_preds,
      symbol_out => transition_530_symbol_out,
      symbol_in  => true);

  transition_531_preds(0) <= place_534_token;
  transition_531 : transition
    port map(
      preds      => transition_531_preds,
      symbol_out => transition_531_symbol_out,
      symbol_in  => LambdaIn(141));

  transition_532_preds(0) <= place_535_token;
  LambdaOut(142) <= transition_532_symbol_out;
  transition_532 : transition
    port map(
      preds      => transition_532_preds,
      symbol_out => transition_532_symbol_out,
      symbol_in  => true);

  transition_533_preds(0) <= place_536_token;
  transition_533 : transition
    port map(
      preds      => transition_533_preds,
      symbol_out => transition_533_symbol_out,
      symbol_in  => LambdaIn(142));

  transition_537_preds(0) <= place_1333_token;
  LambdaOut(143) <= transition_537_symbol_out;
  transition_537 : transition
    port map(
      preds      => transition_537_preds,
      symbol_out => transition_537_symbol_out,
      symbol_in  => true);

  transition_538_preds(0) <= place_541_token;
  transition_538 : transition
    port map(
      preds      => transition_538_preds,
      symbol_out => transition_538_symbol_out,
      symbol_in  => LambdaIn(143));

  transition_539_preds(0) <= place_542_token;
  LambdaOut(144) <= transition_539_symbol_out;
  transition_539 : transition
    port map(
      preds      => transition_539_preds,
      symbol_out => transition_539_symbol_out,
      symbol_in  => true);

  transition_540_preds(0) <= place_543_token;
  transition_540 : transition
    port map(
      preds      => transition_540_preds,
      symbol_out => transition_540_symbol_out,
      symbol_in  => LambdaIn(144));

  transition_544_preds(0) <= place_1330_token;
  transition_544_preds(1) <= place_1331_token;
  transition_544 : transition
    port map(
      preds      => transition_544_preds,
      symbol_out => transition_544_symbol_out,
      symbol_in  => true);

  transition_545_preds(0) <= place_1334_token;
  LambdaOut(145) <= transition_545_symbol_out;
  transition_545 : transition
    port map(
      preds      => transition_545_preds,
      symbol_out => transition_545_symbol_out,
      symbol_in  => true);

  transition_546_preds(0) <= place_549_token;
  transition_546 : transition
    port map(
      preds      => transition_546_preds,
      symbol_out => transition_546_symbol_out,
      symbol_in  => LambdaIn(145));

  transition_547_preds(0) <= place_550_token;
  LambdaOut(146) <= transition_547_symbol_out;
  transition_547 : transition
    port map(
      preds      => transition_547_preds,
      symbol_out => transition_547_symbol_out,
      symbol_in  => true);

  transition_548_preds(0) <= place_551_token;
  transition_548 : transition
    port map(
      preds      => transition_548_preds,
      symbol_out => transition_548_symbol_out,
      symbol_in  => LambdaIn(146));

  transition_553_preds(0) <= place_552_token;
  transition_553 : transition
    port map(
      preds      => transition_553_preds,
      symbol_out => transition_553_symbol_out,
      symbol_in  => LambdaIn(147));

  transition_554_preds(0) <= place_1336_token;
  LambdaOut(147) <= transition_554_symbol_out;
  transition_554 : transition
    port map(
      preds      => transition_554_preds,
      symbol_out => transition_554_symbol_out,
      symbol_in  => true);

  transition_555_preds(0) <= place_1316_token;
  transition_555_preds(1) <= place_1322_token;
  transition_555_preds(2) <= place_1335_token;
  transition_555 : transition
    port map(
      preds      => transition_555_preds,
      symbol_out => transition_555_symbol_out,
      symbol_in  => true);

  transition_556_preds(0) <= place_1339_token;
  LambdaOut(148) <= transition_556_symbol_out;
  transition_556 : transition
    port map(
      preds      => transition_556_preds,
      symbol_out => transition_556_symbol_out,
      symbol_in  => true);

  transition_557_preds(0) <= place_560_token;
  transition_557 : transition
    port map(
      preds      => transition_557_preds,
      symbol_out => transition_557_symbol_out,
      symbol_in  => LambdaIn(148));

  transition_558_preds(0) <= place_561_token;
  LambdaOut(149) <= transition_558_symbol_out;
  transition_558 : transition
    port map(
      preds      => transition_558_preds,
      symbol_out => transition_558_symbol_out,
      symbol_in  => true);

  transition_559_preds(0) <= place_562_token;
  transition_559 : transition
    port map(
      preds      => transition_559_preds,
      symbol_out => transition_559_symbol_out,
      symbol_in  => LambdaIn(149));

  transition_563_preds(0) <= place_1341_token;
  transition_563_preds(1) <= place_1342_token;
  transition_563 : transition
    port map(
      preds      => transition_563_preds,
      symbol_out => transition_563_symbol_out,
      symbol_in  => true);

  transition_564_preds(0) <= place_1340_token;
  LambdaOut(150) <= transition_564_symbol_out;
  transition_564 : transition
    port map(
      preds      => transition_564_preds,
      symbol_out => transition_564_symbol_out,
      symbol_in  => true);

  transition_565_preds(0) <= place_568_token;
  transition_565 : transition
    port map(
      preds      => transition_565_preds,
      symbol_out => transition_565_symbol_out,
      symbol_in  => LambdaIn(150));

  transition_566_preds(0) <= place_569_token;
  LambdaOut(151) <= transition_566_symbol_out;
  transition_566 : transition
    port map(
      preds      => transition_566_preds,
      symbol_out => transition_566_symbol_out,
      symbol_in  => true);

  transition_567_preds(0) <= place_570_token;
  transition_567 : transition
    port map(
      preds      => transition_567_preds,
      symbol_out => transition_567_symbol_out,
      symbol_in  => LambdaIn(151));

  transition_571_preds(0) <= place_1345_token;
  LambdaOut(152) <= transition_571_symbol_out;
  transition_571 : transition
    port map(
      preds      => transition_571_preds,
      symbol_out => transition_571_symbol_out,
      symbol_in  => true);

  transition_572_preds(0) <= place_575_token;
  transition_572 : transition
    port map(
      preds      => transition_572_preds,
      symbol_out => transition_572_symbol_out,
      symbol_in  => LambdaIn(152));

  transition_573_preds(0) <= place_576_token;
  LambdaOut(153) <= transition_573_symbol_out;
  transition_573 : transition
    port map(
      preds      => transition_573_preds,
      symbol_out => transition_573_symbol_out,
      symbol_in  => true);

  transition_574_preds(0) <= place_577_token;
  transition_574 : transition
    port map(
      preds      => transition_574_preds,
      symbol_out => transition_574_symbol_out,
      symbol_in  => LambdaIn(153));

  transition_578_preds(0) <= place_1347_token;
  LambdaOut(154) <= transition_578_symbol_out;
  transition_578 : transition
    port map(
      preds      => transition_578_preds,
      symbol_out => transition_578_symbol_out,
      symbol_in  => true);

  transition_579_preds(0) <= place_582_token;
  transition_579 : transition
    port map(
      preds      => transition_579_preds,
      symbol_out => transition_579_symbol_out,
      symbol_in  => LambdaIn(154));

  transition_580_preds(0) <= place_583_token;
  LambdaOut(155) <= transition_580_symbol_out;
  transition_580 : transition
    port map(
      preds      => transition_580_preds,
      symbol_out => transition_580_symbol_out,
      symbol_in  => true);

  transition_581_preds(0) <= place_584_token;
  transition_581 : transition
    port map(
      preds      => transition_581_preds,
      symbol_out => transition_581_symbol_out,
      symbol_in  => LambdaIn(155));

  transition_585_preds(0) <= place_1348_token;
  LambdaOut(156) <= transition_585_symbol_out;
  transition_585 : transition
    port map(
      preds      => transition_585_preds,
      symbol_out => transition_585_symbol_out,
      symbol_in  => true);

  transition_586_preds(0) <= place_589_token;
  transition_586 : transition
    port map(
      preds      => transition_586_preds,
      symbol_out => transition_586_symbol_out,
      symbol_in  => LambdaIn(156));

  transition_587_preds(0) <= place_590_token;
  LambdaOut(157) <= transition_587_symbol_out;
  transition_587 : transition
    port map(
      preds      => transition_587_preds,
      symbol_out => transition_587_symbol_out,
      symbol_in  => true);

  transition_588_preds(0) <= place_591_token;
  transition_588 : transition
    port map(
      preds      => transition_588_preds,
      symbol_out => transition_588_symbol_out,
      symbol_in  => LambdaIn(157));

  transition_592_preds(0) <= place_1346_token;
  transition_592_preds(1) <= place_1344_token;
  transition_592 : transition
    port map(
      preds      => transition_592_preds,
      symbol_out => transition_592_symbol_out,
      symbol_in  => true);

  transition_593_preds(0) <= place_1351_token;
  LambdaOut(158) <= transition_593_symbol_out;
  transition_593 : transition
    port map(
      preds      => transition_593_preds,
      symbol_out => transition_593_symbol_out,
      symbol_in  => true);

  transition_594_preds(0) <= place_597_token;
  transition_594 : transition
    port map(
      preds      => transition_594_preds,
      symbol_out => transition_594_symbol_out,
      symbol_in  => LambdaIn(158));

  transition_595_preds(0) <= place_598_token;
  LambdaOut(159) <= transition_595_symbol_out;
  transition_595 : transition
    port map(
      preds      => transition_595_preds,
      symbol_out => transition_595_symbol_out,
      symbol_in  => true);

  transition_596_preds(0) <= place_599_token;
  transition_596 : transition
    port map(
      preds      => transition_596_preds,
      symbol_out => transition_596_symbol_out,
      symbol_in  => LambdaIn(159));

  transition_600_preds(0) <= place_1352_token;
  LambdaOut(160) <= transition_600_symbol_out;
  transition_600 : transition
    port map(
      preds      => transition_600_preds,
      symbol_out => transition_600_symbol_out,
      symbol_in  => true);

  transition_601_preds(0) <= place_604_token;
  transition_601 : transition
    port map(
      preds      => transition_601_preds,
      symbol_out => transition_601_symbol_out,
      symbol_in  => LambdaIn(160));

  transition_602_preds(0) <= place_605_token;
  LambdaOut(161) <= transition_602_symbol_out;
  transition_602 : transition
    port map(
      preds      => transition_602_preds,
      symbol_out => transition_602_symbol_out,
      symbol_in  => true);

  transition_603_preds(0) <= place_606_token;
  transition_603 : transition
    port map(
      preds      => transition_603_preds,
      symbol_out => transition_603_symbol_out,
      symbol_in  => LambdaIn(161));

  transition_607_preds(0) <= place_1349_token;
  transition_607_preds(1) <= place_1350_token;
  transition_607 : transition
    port map(
      preds      => transition_607_preds,
      symbol_out => transition_607_symbol_out,
      symbol_in  => true);

  transition_608_preds(0) <= place_1353_token;
  LambdaOut(162) <= transition_608_symbol_out;
  transition_608 : transition
    port map(
      preds      => transition_608_preds,
      symbol_out => transition_608_symbol_out,
      symbol_in  => true);

  transition_609_preds(0) <= place_612_token;
  transition_609 : transition
    port map(
      preds      => transition_609_preds,
      symbol_out => transition_609_symbol_out,
      symbol_in  => LambdaIn(162));

  transition_610_preds(0) <= place_613_token;
  LambdaOut(163) <= transition_610_symbol_out;
  transition_610 : transition
    port map(
      preds      => transition_610_preds,
      symbol_out => transition_610_symbol_out,
      symbol_in  => true);

  transition_611_preds(0) <= place_614_token;
  transition_611 : transition
    port map(
      preds      => transition_611_preds,
      symbol_out => transition_611_symbol_out,
      symbol_in  => LambdaIn(163));

  transition_616_preds(0) <= place_615_token;
  transition_616 : transition
    port map(
      preds      => transition_616_preds,
      symbol_out => transition_616_symbol_out,
      symbol_in  => LambdaIn(164));

  transition_617_preds(0) <= place_1355_token;
  LambdaOut(164) <= transition_617_symbol_out;
  transition_617 : transition
    port map(
      preds      => transition_617_preds,
      symbol_out => transition_617_symbol_out,
      symbol_in  => true);

  transition_618_preds(0) <= place_1337_token;
  transition_618_preds(1) <= place_1343_token;
  transition_618_preds(2) <= place_1354_token;
  transition_618 : transition
    port map(
      preds      => transition_618_preds,
      symbol_out => transition_618_symbol_out,
      symbol_in  => true);

  transition_619_preds(0) <= place_1359_token;
  LambdaOut(165) <= transition_619_symbol_out;
  transition_619 : transition
    port map(
      preds      => transition_619_preds,
      symbol_out => transition_619_symbol_out,
      symbol_in  => true);

  transition_620_preds(0) <= place_623_token;
  transition_620 : transition
    port map(
      preds      => transition_620_preds,
      symbol_out => transition_620_symbol_out,
      symbol_in  => LambdaIn(165));

  transition_621_preds(0) <= place_624_token;
  LambdaOut(166) <= transition_621_symbol_out;
  transition_621 : transition
    port map(
      preds      => transition_621_preds,
      symbol_out => transition_621_symbol_out,
      symbol_in  => true);

  transition_622_preds(0) <= place_625_token;
  transition_622 : transition
    port map(
      preds      => transition_622_preds,
      symbol_out => transition_622_symbol_out,
      symbol_in  => LambdaIn(166));

  transition_626_preds(0) <= place_1361_token;
  transition_626_preds(1) <= place_1362_token;
  transition_626 : transition
    port map(
      preds      => transition_626_preds,
      symbol_out => transition_626_symbol_out,
      symbol_in  => true);

  transition_627_preds(0) <= place_1360_token;
  LambdaOut(167) <= transition_627_symbol_out;
  transition_627 : transition
    port map(
      preds      => transition_627_preds,
      symbol_out => transition_627_symbol_out,
      symbol_in  => true);

  transition_628_preds(0) <= place_631_token;
  transition_628 : transition
    port map(
      preds      => transition_628_preds,
      symbol_out => transition_628_symbol_out,
      symbol_in  => LambdaIn(167));

  transition_629_preds(0) <= place_632_token;
  LambdaOut(168) <= transition_629_symbol_out;
  transition_629 : transition
    port map(
      preds      => transition_629_preds,
      symbol_out => transition_629_symbol_out,
      symbol_in  => true);

  transition_630_preds(0) <= place_633_token;
  transition_630 : transition
    port map(
      preds      => transition_630_preds,
      symbol_out => transition_630_symbol_out,
      symbol_in  => LambdaIn(168));

  transition_634_preds(0) <= place_1365_token;
  LambdaOut(169) <= transition_634_symbol_out;
  transition_634 : transition
    port map(
      preds      => transition_634_preds,
      symbol_out => transition_634_symbol_out,
      symbol_in  => true);

  transition_635_preds(0) <= place_638_token;
  transition_635 : transition
    port map(
      preds      => transition_635_preds,
      symbol_out => transition_635_symbol_out,
      symbol_in  => LambdaIn(169));

  transition_636_preds(0) <= place_639_token;
  LambdaOut(170) <= transition_636_symbol_out;
  transition_636 : transition
    port map(
      preds      => transition_636_preds,
      symbol_out => transition_636_symbol_out,
      symbol_in  => true);

  transition_637_preds(0) <= place_640_token;
  transition_637 : transition
    port map(
      preds      => transition_637_preds,
      symbol_out => transition_637_symbol_out,
      symbol_in  => LambdaIn(170));

  transition_641_preds(0) <= place_1367_token;
  LambdaOut(171) <= transition_641_symbol_out;
  transition_641 : transition
    port map(
      preds      => transition_641_preds,
      symbol_out => transition_641_symbol_out,
      symbol_in  => true);

  transition_642_preds(0) <= place_645_token;
  transition_642 : transition
    port map(
      preds      => transition_642_preds,
      symbol_out => transition_642_symbol_out,
      symbol_in  => LambdaIn(171));

  transition_643_preds(0) <= place_646_token;
  LambdaOut(172) <= transition_643_symbol_out;
  transition_643 : transition
    port map(
      preds      => transition_643_preds,
      symbol_out => transition_643_symbol_out,
      symbol_in  => true);

  transition_644_preds(0) <= place_647_token;
  transition_644 : transition
    port map(
      preds      => transition_644_preds,
      symbol_out => transition_644_symbol_out,
      symbol_in  => LambdaIn(172));

  transition_648_preds(0) <= place_1368_token;
  LambdaOut(173) <= transition_648_symbol_out;
  transition_648 : transition
    port map(
      preds      => transition_648_preds,
      symbol_out => transition_648_symbol_out,
      symbol_in  => true);

  transition_649_preds(0) <= place_652_token;
  transition_649 : transition
    port map(
      preds      => transition_649_preds,
      symbol_out => transition_649_symbol_out,
      symbol_in  => LambdaIn(173));

  transition_650_preds(0) <= place_653_token;
  LambdaOut(174) <= transition_650_symbol_out;
  transition_650 : transition
    port map(
      preds      => transition_650_preds,
      symbol_out => transition_650_symbol_out,
      symbol_in  => true);

  transition_651_preds(0) <= place_654_token;
  transition_651 : transition
    port map(
      preds      => transition_651_preds,
      symbol_out => transition_651_symbol_out,
      symbol_in  => LambdaIn(174));

  transition_655_preds(0) <= place_1366_token;
  transition_655_preds(1) <= place_1364_token;
  transition_655 : transition
    port map(
      preds      => transition_655_preds,
      symbol_out => transition_655_symbol_out,
      symbol_in  => true);

  transition_656_preds(0) <= place_1372_token;
  LambdaOut(175) <= transition_656_symbol_out;
  transition_656 : transition
    port map(
      preds      => transition_656_preds,
      symbol_out => transition_656_symbol_out,
      symbol_in  => true);

  transition_657_preds(0) <= place_660_token;
  transition_657 : transition
    port map(
      preds      => transition_657_preds,
      symbol_out => transition_657_symbol_out,
      symbol_in  => LambdaIn(175));

  transition_658_preds(0) <= place_661_token;
  LambdaOut(176) <= transition_658_symbol_out;
  transition_658 : transition
    port map(
      preds      => transition_658_preds,
      symbol_out => transition_658_symbol_out,
      symbol_in  => true);

  transition_659_preds(0) <= place_662_token;
  transition_659 : transition
    port map(
      preds      => transition_659_preds,
      symbol_out => transition_659_symbol_out,
      symbol_in  => LambdaIn(176));

  transition_663_preds(0) <= place_1373_token;
  LambdaOut(177) <= transition_663_symbol_out;
  transition_663 : transition
    port map(
      preds      => transition_663_preds,
      symbol_out => transition_663_symbol_out,
      symbol_in  => true);

  transition_664_preds(0) <= place_667_token;
  transition_664 : transition
    port map(
      preds      => transition_664_preds,
      symbol_out => transition_664_symbol_out,
      symbol_in  => LambdaIn(177));

  transition_665_preds(0) <= place_668_token;
  LambdaOut(178) <= transition_665_symbol_out;
  transition_665 : transition
    port map(
      preds      => transition_665_preds,
      symbol_out => transition_665_symbol_out,
      symbol_in  => true);

  transition_666_preds(0) <= place_669_token;
  transition_666 : transition
    port map(
      preds      => transition_666_preds,
      symbol_out => transition_666_symbol_out,
      symbol_in  => LambdaIn(178));

  transition_670_preds(0) <= place_1370_token;
  transition_670_preds(1) <= place_1371_token;
  transition_670 : transition
    port map(
      preds      => transition_670_preds,
      symbol_out => transition_670_symbol_out,
      symbol_in  => true);

  transition_671_preds(0) <= place_1374_token;
  LambdaOut(179) <= transition_671_symbol_out;
  transition_671 : transition
    port map(
      preds      => transition_671_preds,
      symbol_out => transition_671_symbol_out,
      symbol_in  => true);

  transition_672_preds(0) <= place_675_token;
  transition_672 : transition
    port map(
      preds      => transition_672_preds,
      symbol_out => transition_672_symbol_out,
      symbol_in  => LambdaIn(179));

  transition_673_preds(0) <= place_676_token;
  LambdaOut(180) <= transition_673_symbol_out;
  transition_673 : transition
    port map(
      preds      => transition_673_preds,
      symbol_out => transition_673_symbol_out,
      symbol_in  => true);

  transition_674_preds(0) <= place_677_token;
  transition_674 : transition
    port map(
      preds      => transition_674_preds,
      symbol_out => transition_674_symbol_out,
      symbol_in  => LambdaIn(180));

  transition_679_preds(0) <= place_678_token;
  transition_679 : transition
    port map(
      preds      => transition_679_preds,
      symbol_out => transition_679_symbol_out,
      symbol_in  => LambdaIn(181));

  transition_680_preds(0) <= place_1376_token;
  LambdaOut(181) <= transition_680_symbol_out;
  transition_680 : transition
    port map(
      preds      => transition_680_preds,
      symbol_out => transition_680_symbol_out,
      symbol_in  => true);

  transition_681_preds(0) <= place_1356_token;
  transition_681_preds(1) <= place_1363_token;
  transition_681_preds(2) <= place_1375_token;
  transition_681 : transition
    port map(
      preds      => transition_681_preds,
      symbol_out => transition_681_symbol_out,
      symbol_in  => true);

  transition_682_preds(0) <= place_1377_token;
  transition_682 : transition
    port map(
      preds      => transition_682_preds,
      symbol_out => transition_682_symbol_out,
      symbol_in  => true);

  transition_683_preds(0) <= place_1379_token;
  LambdaOut(182) <= transition_683_symbol_out;
  transition_683 : transition
    port map(
      preds      => transition_683_preds,
      symbol_out => transition_683_symbol_out,
      symbol_in  => true);

  transition_684_preds(0) <= place_687_token;
  transition_684 : transition
    port map(
      preds      => transition_684_preds,
      symbol_out => transition_684_symbol_out,
      symbol_in  => LambdaIn(182));

  transition_685_preds(0) <= place_688_token;
  LambdaOut(183) <= transition_685_symbol_out;
  transition_685 : transition
    port map(
      preds      => transition_685_preds,
      symbol_out => transition_685_symbol_out,
      symbol_in  => true);

  transition_686_preds(0) <= place_689_token;
  transition_686 : transition
    port map(
      preds      => transition_686_preds,
      symbol_out => transition_686_symbol_out,
      symbol_in  => LambdaIn(183));

  transition_690_preds(0) <= place_1381_token;
  LambdaOut(184) <= transition_690_symbol_out;
  transition_690 : transition
    port map(
      preds      => transition_690_preds,
      symbol_out => transition_690_symbol_out,
      symbol_in  => true);

  transition_691_preds(0) <= place_694_token;
  transition_691 : transition
    port map(
      preds      => transition_691_preds,
      symbol_out => transition_691_symbol_out,
      symbol_in  => LambdaIn(184));

  transition_692_preds(0) <= place_695_token;
  LambdaOut(185) <= transition_692_symbol_out;
  transition_692 : transition
    port map(
      preds      => transition_692_preds,
      symbol_out => transition_692_symbol_out,
      symbol_in  => true);

  transition_693_preds(0) <= place_696_token;
  transition_693 : transition
    port map(
      preds      => transition_693_preds,
      symbol_out => transition_693_symbol_out,
      symbol_in  => LambdaIn(185));

  transition_697_preds(0) <= place_1383_token;
  LambdaOut(186) <= transition_697_symbol_out;
  transition_697 : transition
    port map(
      preds      => transition_697_preds,
      symbol_out => transition_697_symbol_out,
      symbol_in  => true);

  transition_698_preds(0) <= place_701_token;
  transition_698 : transition
    port map(
      preds      => transition_698_preds,
      symbol_out => transition_698_symbol_out,
      symbol_in  => LambdaIn(186));

  transition_699_preds(0) <= place_702_token;
  LambdaOut(187) <= transition_699_symbol_out;
  transition_699 : transition
    port map(
      preds      => transition_699_preds,
      symbol_out => transition_699_symbol_out,
      symbol_in  => true);

  transition_700_preds(0) <= place_703_token;
  transition_700 : transition
    port map(
      preds      => transition_700_preds,
      symbol_out => transition_700_symbol_out,
      symbol_in  => LambdaIn(187));

  transition_704_preds(0) <= place_1380_token;
  transition_704_preds(1) <= place_1378_token;
  transition_704 : transition
    port map(
      preds      => transition_704_preds,
      symbol_out => transition_704_symbol_out,
      symbol_in  => true);

  transition_705_preds(0) <= place_1386_token;
  LambdaOut(188) <= transition_705_symbol_out;
  transition_705 : transition
    port map(
      preds      => transition_705_preds,
      symbol_out => transition_705_symbol_out,
      symbol_in  => true);

  transition_706_preds(0) <= place_709_token;
  transition_706 : transition
    port map(
      preds      => transition_706_preds,
      symbol_out => transition_706_symbol_out,
      symbol_in  => LambdaIn(188));

  transition_707_preds(0) <= place_710_token;
  LambdaOut(189) <= transition_707_symbol_out;
  transition_707 : transition
    port map(
      preds      => transition_707_preds,
      symbol_out => transition_707_symbol_out,
      symbol_in  => true);

  transition_708_preds(0) <= place_711_token;
  transition_708 : transition
    port map(
      preds      => transition_708_preds,
      symbol_out => transition_708_symbol_out,
      symbol_in  => LambdaIn(189));

  transition_712_preds(0) <= place_1387_token;
  LambdaOut(190) <= transition_712_symbol_out;
  transition_712 : transition
    port map(
      preds      => transition_712_preds,
      symbol_out => transition_712_symbol_out,
      symbol_in  => true);

  transition_713_preds(0) <= place_716_token;
  transition_713 : transition
    port map(
      preds      => transition_713_preds,
      symbol_out => transition_713_symbol_out,
      symbol_in  => LambdaIn(190));

  transition_714_preds(0) <= place_717_token;
  LambdaOut(191) <= transition_714_symbol_out;
  transition_714 : transition
    port map(
      preds      => transition_714_preds,
      symbol_out => transition_714_symbol_out,
      symbol_in  => true);

  transition_715_preds(0) <= place_718_token;
  transition_715 : transition
    port map(
      preds      => transition_715_preds,
      symbol_out => transition_715_symbol_out,
      symbol_in  => LambdaIn(191));

  transition_719_preds(0) <= place_1384_token;
  transition_719_preds(1) <= place_1385_token;
  transition_719 : transition
    port map(
      preds      => transition_719_preds,
      symbol_out => transition_719_symbol_out,
      symbol_in  => true);

  transition_720_preds(0) <= place_1388_token;
  LambdaOut(192) <= transition_720_symbol_out;
  transition_720 : transition
    port map(
      preds      => transition_720_preds,
      symbol_out => transition_720_symbol_out,
      symbol_in  => true);

  transition_721_preds(0) <= place_724_token;
  transition_721 : transition
    port map(
      preds      => transition_721_preds,
      symbol_out => transition_721_symbol_out,
      symbol_in  => LambdaIn(192));

  transition_722_preds(0) <= place_725_token;
  LambdaOut(193) <= transition_722_symbol_out;
  transition_722 : transition
    port map(
      preds      => transition_722_preds,
      symbol_out => transition_722_symbol_out,
      symbol_in  => true);

  transition_723_preds(0) <= place_726_token;
  transition_723 : transition
    port map(
      preds      => transition_723_preds,
      symbol_out => transition_723_symbol_out,
      symbol_in  => LambdaIn(193));

  transition_728_preds(0) <= place_727_token;
  transition_728 : transition
    port map(
      preds      => transition_728_preds,
      symbol_out => transition_728_symbol_out,
      symbol_in  => LambdaIn(194));

  transition_729_preds(0) <= place_1390_token;
  LambdaOut(194) <= transition_729_symbol_out;
  transition_729 : transition
    port map(
      preds      => transition_729_preds,
      symbol_out => transition_729_symbol_out,
      symbol_in  => true);

  transition_730_preds(0) <= place_1389_token;
  transition_730_preds(1) <= place_1394_token;
  transition_730 : transition
    port map(
      preds      => transition_730_preds,
      symbol_out => transition_730_symbol_out,
      symbol_in  => true);

  transition_732_preds(0) <= place_731_token;
  transition_732 : transition
    port map(
      preds      => transition_732_preds,
      symbol_out => transition_732_symbol_out,
      symbol_in  => LambdaIn(195));

  transition_733_preds(0) <= place_1392_token;
  LambdaOut(195) <= transition_733_symbol_out;
  transition_733 : transition
    port map(
      preds      => transition_733_preds,
      symbol_out => transition_733_symbol_out,
      symbol_in  => true);

  transition_734_preds(0) <= place_1396_token;
  LambdaOut(196) <= transition_734_symbol_out;
  transition_734 : transition
    port map(
      preds      => transition_734_preds,
      symbol_out => transition_734_symbol_out,
      symbol_in  => true);

  transition_735_preds(0) <= place_738_token;
  transition_735 : transition
    port map(
      preds      => transition_735_preds,
      symbol_out => transition_735_symbol_out,
      symbol_in  => LambdaIn(196));

  transition_736_preds(0) <= place_739_token;
  LambdaOut(197) <= transition_736_symbol_out;
  transition_736 : transition
    port map(
      preds      => transition_736_preds,
      symbol_out => transition_736_symbol_out,
      symbol_in  => true);

  transition_737_preds(0) <= place_740_token;
  transition_737 : transition
    port map(
      preds      => transition_737_preds,
      symbol_out => transition_737_symbol_out,
      symbol_in  => LambdaIn(197));

  transition_741_preds(0) <= place_1398_token;
  LambdaOut(198) <= transition_741_symbol_out;
  transition_741 : transition
    port map(
      preds      => transition_741_preds,
      symbol_out => transition_741_symbol_out,
      symbol_in  => true);

  transition_742_preds(0) <= place_745_token;
  transition_742 : transition
    port map(
      preds      => transition_742_preds,
      symbol_out => transition_742_symbol_out,
      symbol_in  => LambdaIn(198));

  transition_743_preds(0) <= place_746_token;
  LambdaOut(199) <= transition_743_symbol_out;
  transition_743 : transition
    port map(
      preds      => transition_743_preds,
      symbol_out => transition_743_symbol_out,
      symbol_in  => true);

  transition_744_preds(0) <= place_747_token;
  transition_744 : transition
    port map(
      preds      => transition_744_preds,
      symbol_out => transition_744_symbol_out,
      symbol_in  => LambdaIn(199));

  transition_748_preds(0) <= place_1399_token;
  LambdaOut(200) <= transition_748_symbol_out;
  transition_748 : transition
    port map(
      preds      => transition_748_preds,
      symbol_out => transition_748_symbol_out,
      symbol_in  => true);

  transition_749_preds(0) <= place_752_token;
  transition_749 : transition
    port map(
      preds      => transition_749_preds,
      symbol_out => transition_749_symbol_out,
      symbol_in  => LambdaIn(200));

  transition_750_preds(0) <= place_753_token;
  LambdaOut(201) <= transition_750_symbol_out;
  transition_750 : transition
    port map(
      preds      => transition_750_preds,
      symbol_out => transition_750_symbol_out,
      symbol_in  => true);

  transition_751_preds(0) <= place_754_token;
  transition_751 : transition
    port map(
      preds      => transition_751_preds,
      symbol_out => transition_751_symbol_out,
      symbol_in  => LambdaIn(201));

  transition_755_preds(0) <= place_1395_token;
  transition_755_preds(1) <= place_1397_token;
  transition_755 : transition
    port map(
      preds      => transition_755_preds,
      symbol_out => transition_755_symbol_out,
      symbol_in  => true);

  transition_756_preds(0) <= place_1403_token;
  LambdaOut(202) <= transition_756_symbol_out;
  transition_756 : transition
    port map(
      preds      => transition_756_preds,
      symbol_out => transition_756_symbol_out,
      symbol_in  => true);

  transition_757_preds(0) <= place_760_token;
  transition_757 : transition
    port map(
      preds      => transition_757_preds,
      symbol_out => transition_757_symbol_out,
      symbol_in  => LambdaIn(202));

  transition_758_preds(0) <= place_761_token;
  LambdaOut(203) <= transition_758_symbol_out;
  transition_758 : transition
    port map(
      preds      => transition_758_preds,
      symbol_out => transition_758_symbol_out,
      symbol_in  => true);

  transition_759_preds(0) <= place_762_token;
  transition_759 : transition
    port map(
      preds      => transition_759_preds,
      symbol_out => transition_759_symbol_out,
      symbol_in  => LambdaIn(203));

  transition_763_preds(0) <= place_1404_token;
  LambdaOut(204) <= transition_763_symbol_out;
  transition_763 : transition
    port map(
      preds      => transition_763_preds,
      symbol_out => transition_763_symbol_out,
      symbol_in  => true);

  transition_764_preds(0) <= place_767_token;
  transition_764 : transition
    port map(
      preds      => transition_764_preds,
      symbol_out => transition_764_symbol_out,
      symbol_in  => LambdaIn(204));

  transition_765_preds(0) <= place_768_token;
  LambdaOut(205) <= transition_765_symbol_out;
  transition_765 : transition
    port map(
      preds      => transition_765_preds,
      symbol_out => transition_765_symbol_out,
      symbol_in  => true);

  transition_766_preds(0) <= place_769_token;
  transition_766 : transition
    port map(
      preds      => transition_766_preds,
      symbol_out => transition_766_symbol_out,
      symbol_in  => LambdaIn(205));

  transition_770_preds(0) <= place_1402_token;
  transition_770_preds(1) <= place_1400_token;
  transition_770 : transition
    port map(
      preds      => transition_770_preds,
      symbol_out => transition_770_symbol_out,
      symbol_in  => true);

  transition_771_preds(0) <= place_1405_token;
  LambdaOut(206) <= transition_771_symbol_out;
  transition_771 : transition
    port map(
      preds      => transition_771_preds,
      symbol_out => transition_771_symbol_out,
      symbol_in  => true);

  transition_772_preds(0) <= place_775_token;
  transition_772 : transition
    port map(
      preds      => transition_772_preds,
      symbol_out => transition_772_symbol_out,
      symbol_in  => LambdaIn(206));

  transition_773_preds(0) <= place_776_token;
  LambdaOut(207) <= transition_773_symbol_out;
  transition_773 : transition
    port map(
      preds      => transition_773_preds,
      symbol_out => transition_773_symbol_out,
      symbol_in  => true);

  transition_774_preds(0) <= place_777_token;
  transition_774 : transition
    port map(
      preds      => transition_774_preds,
      symbol_out => transition_774_symbol_out,
      symbol_in  => LambdaIn(207));

  transition_779_preds(0) <= place_778_token;
  transition_779 : transition
    port map(
      preds      => transition_779_preds,
      symbol_out => transition_779_symbol_out,
      symbol_in  => LambdaIn(208));

  transition_780_preds(0) <= place_1408_token;
  LambdaOut(208) <= transition_780_symbol_out;
  transition_780 : transition
    port map(
      preds      => transition_780_preds,
      symbol_out => transition_780_symbol_out,
      symbol_in  => true);

  transition_781_preds(0) <= place_1407_token;
  transition_781_preds(1) <= place_1412_token;
  transition_781 : transition
    port map(
      preds      => transition_781_preds,
      symbol_out => transition_781_symbol_out,
      symbol_in  => true);

  transition_783_preds(0) <= place_782_token;
  transition_783 : transition
    port map(
      preds      => transition_783_preds,
      symbol_out => transition_783_symbol_out,
      symbol_in  => LambdaIn(209));

  transition_784_preds(0) <= place_1409_token;
  LambdaOut(209) <= transition_784_symbol_out;
  transition_784 : transition
    port map(
      preds      => transition_784_preds,
      symbol_out => transition_784_symbol_out,
      symbol_in  => true);

  transition_785_preds(0) <= place_1413_token;
  LambdaOut(210) <= transition_785_symbol_out;
  transition_785 : transition
    port map(
      preds      => transition_785_preds,
      symbol_out => transition_785_symbol_out,
      symbol_in  => true);

  transition_786_preds(0) <= place_789_token;
  transition_786 : transition
    port map(
      preds      => transition_786_preds,
      symbol_out => transition_786_symbol_out,
      symbol_in  => LambdaIn(210));

  transition_787_preds(0) <= place_790_token;
  LambdaOut(211) <= transition_787_symbol_out;
  transition_787 : transition
    port map(
      preds      => transition_787_preds,
      symbol_out => transition_787_symbol_out,
      symbol_in  => true);

  transition_788_preds(0) <= place_791_token;
  transition_788 : transition
    port map(
      preds      => transition_788_preds,
      symbol_out => transition_788_symbol_out,
      symbol_in  => LambdaIn(211));

  transition_792_preds(0) <= place_1393_token;
  transition_792_preds(1) <= place_1410_token;
  transition_792 : transition
    port map(
      preds      => transition_792_preds,
      symbol_out => transition_792_symbol_out,
      symbol_in  => true);

  transition_793_preds(0) <= place_1414_token;
  LambdaOut(212) <= transition_793_symbol_out;
  transition_793 : transition
    port map(
      preds      => transition_793_preds,
      symbol_out => transition_793_symbol_out,
      symbol_in  => true);

  transition_794_preds(0) <= place_797_token;
  transition_794 : transition
    port map(
      preds      => transition_794_preds,
      symbol_out => transition_794_symbol_out,
      symbol_in  => LambdaIn(212));

  transition_795_preds(0) <= place_798_token;
  LambdaOut(213) <= transition_795_symbol_out;
  transition_795 : transition
    port map(
      preds      => transition_795_preds,
      symbol_out => transition_795_symbol_out,
      symbol_in  => true);

  transition_796_preds(0) <= place_799_token;
  transition_796 : transition
    port map(
      preds      => transition_796_preds,
      symbol_out => transition_796_symbol_out,
      symbol_in  => LambdaIn(213));

  transition_800_preds(0) <= place_1417_token;
  LambdaOut(214) <= transition_800_symbol_out;
  transition_800 : transition
    port map(
      preds      => transition_800_preds,
      symbol_out => transition_800_symbol_out,
      symbol_in  => true);

  transition_801_preds(0) <= place_804_token;
  transition_801 : transition
    port map(
      preds      => transition_801_preds,
      symbol_out => transition_801_symbol_out,
      symbol_in  => LambdaIn(214));

  transition_802_preds(0) <= place_805_token;
  LambdaOut(215) <= transition_802_symbol_out;
  transition_802 : transition
    port map(
      preds      => transition_802_preds,
      symbol_out => transition_802_symbol_out,
      symbol_in  => true);

  transition_803_preds(0) <= place_806_token;
  transition_803 : transition
    port map(
      preds      => transition_803_preds,
      symbol_out => transition_803_symbol_out,
      symbol_in  => LambdaIn(215));

  transition_807_preds(0) <= place_1419_token;
  LambdaOut(216) <= transition_807_symbol_out;
  transition_807 : transition
    port map(
      preds      => transition_807_preds,
      symbol_out => transition_807_symbol_out,
      symbol_in  => true);

  transition_808_preds(0) <= place_811_token;
  transition_808 : transition
    port map(
      preds      => transition_808_preds,
      symbol_out => transition_808_symbol_out,
      symbol_in  => LambdaIn(216));

  transition_809_preds(0) <= place_812_token;
  LambdaOut(217) <= transition_809_symbol_out;
  transition_809 : transition
    port map(
      preds      => transition_809_preds,
      symbol_out => transition_809_symbol_out,
      symbol_in  => true);

  transition_810_preds(0) <= place_813_token;
  transition_810 : transition
    port map(
      preds      => transition_810_preds,
      symbol_out => transition_810_symbol_out,
      symbol_in  => LambdaIn(217));

  transition_814_preds(0) <= place_1420_token;
  LambdaOut(218) <= transition_814_symbol_out;
  transition_814 : transition
    port map(
      preds      => transition_814_preds,
      symbol_out => transition_814_symbol_out,
      symbol_in  => true);

  transition_815_preds(0) <= place_818_token;
  transition_815 : transition
    port map(
      preds      => transition_815_preds,
      symbol_out => transition_815_symbol_out,
      symbol_in  => LambdaIn(218));

  transition_816_preds(0) <= place_819_token;
  LambdaOut(219) <= transition_816_symbol_out;
  transition_816 : transition
    port map(
      preds      => transition_816_preds,
      symbol_out => transition_816_symbol_out,
      symbol_in  => true);

  transition_817_preds(0) <= place_820_token;
  transition_817 : transition
    port map(
      preds      => transition_817_preds,
      symbol_out => transition_817_symbol_out,
      symbol_in  => LambdaIn(219));

  transition_821_preds(0) <= place_1416_token;
  transition_821_preds(1) <= place_1418_token;
  transition_821 : transition
    port map(
      preds      => transition_821_preds,
      symbol_out => transition_821_symbol_out,
      symbol_in  => true);

  transition_822_preds(0) <= place_1423_token;
  LambdaOut(220) <= transition_822_symbol_out;
  transition_822 : transition
    port map(
      preds      => transition_822_preds,
      symbol_out => transition_822_symbol_out,
      symbol_in  => true);

  transition_823_preds(0) <= place_826_token;
  transition_823 : transition
    port map(
      preds      => transition_823_preds,
      symbol_out => transition_823_symbol_out,
      symbol_in  => LambdaIn(220));

  transition_824_preds(0) <= place_827_token;
  LambdaOut(221) <= transition_824_symbol_out;
  transition_824 : transition
    port map(
      preds      => transition_824_preds,
      symbol_out => transition_824_symbol_out,
      symbol_in  => true);

  transition_825_preds(0) <= place_828_token;
  transition_825 : transition
    port map(
      preds      => transition_825_preds,
      symbol_out => transition_825_symbol_out,
      symbol_in  => LambdaIn(221));

  transition_829_preds(0) <= place_1424_token;
  LambdaOut(222) <= transition_829_symbol_out;
  transition_829 : transition
    port map(
      preds      => transition_829_preds,
      symbol_out => transition_829_symbol_out,
      symbol_in  => true);

  transition_830_preds(0) <= place_833_token;
  transition_830 : transition
    port map(
      preds      => transition_830_preds,
      symbol_out => transition_830_symbol_out,
      symbol_in  => LambdaIn(222));

  transition_831_preds(0) <= place_834_token;
  LambdaOut(223) <= transition_831_symbol_out;
  transition_831 : transition
    port map(
      preds      => transition_831_preds,
      symbol_out => transition_831_symbol_out,
      symbol_in  => true);

  transition_832_preds(0) <= place_835_token;
  transition_832 : transition
    port map(
      preds      => transition_832_preds,
      symbol_out => transition_832_symbol_out,
      symbol_in  => LambdaIn(223));

  transition_836_preds(0) <= place_1421_token;
  transition_836_preds(1) <= place_1422_token;
  transition_836 : transition
    port map(
      preds      => transition_836_preds,
      symbol_out => transition_836_symbol_out,
      symbol_in  => true);

  transition_837_preds(0) <= place_1425_token;
  LambdaOut(224) <= transition_837_symbol_out;
  transition_837 : transition
    port map(
      preds      => transition_837_preds,
      symbol_out => transition_837_symbol_out,
      symbol_in  => true);

  transition_838_preds(0) <= place_841_token;
  transition_838 : transition
    port map(
      preds      => transition_838_preds,
      symbol_out => transition_838_symbol_out,
      symbol_in  => LambdaIn(224));

  transition_839_preds(0) <= place_842_token;
  LambdaOut(225) <= transition_839_symbol_out;
  transition_839 : transition
    port map(
      preds      => transition_839_preds,
      symbol_out => transition_839_symbol_out,
      symbol_in  => true);

  transition_840_preds(0) <= place_843_token;
  transition_840 : transition
    port map(
      preds      => transition_840_preds,
      symbol_out => transition_840_symbol_out,
      symbol_in  => LambdaIn(225));

  transition_845_preds(0) <= place_844_token;
  transition_845 : transition
    port map(
      preds      => transition_845_preds,
      symbol_out => transition_845_symbol_out,
      symbol_in  => LambdaIn(226));

  transition_846_preds(0) <= place_1427_token;
  LambdaOut(226) <= transition_846_symbol_out;
  transition_846 : transition
    port map(
      preds      => transition_846_preds,
      symbol_out => transition_846_symbol_out,
      symbol_in  => true);

  transition_847_preds(0) <= place_1415_token;
  transition_847_preds(1) <= place_1426_token;
  transition_847 : transition
    port map(
      preds      => transition_847_preds,
      symbol_out => transition_847_symbol_out,
      symbol_in  => true);

  transition_848_preds(0) <= place_1428_token;
  transition_848 : transition
    port map(
      preds      => transition_848_preds,
      symbol_out => transition_848_symbol_out,
      symbol_in  => true);

  transition_849_preds(0) <= place_1430_token;
  LambdaOut(227) <= transition_849_symbol_out;
  transition_849 : transition
    port map(
      preds      => transition_849_preds,
      symbol_out => transition_849_symbol_out,
      symbol_in  => true);

  transition_850_preds(0) <= place_853_token;
  transition_850 : transition
    port map(
      preds      => transition_850_preds,
      symbol_out => transition_850_symbol_out,
      symbol_in  => LambdaIn(227));

  transition_851_preds(0) <= place_854_token;
  LambdaOut(228) <= transition_851_symbol_out;
  transition_851 : transition
    port map(
      preds      => transition_851_preds,
      symbol_out => transition_851_symbol_out,
      symbol_in  => true);

  transition_852_preds(0) <= place_855_token;
  transition_852 : transition
    port map(
      preds      => transition_852_preds,
      symbol_out => transition_852_symbol_out,
      symbol_in  => LambdaIn(228));

  transition_856_preds(0) <= place_1432_token;
  LambdaOut(229) <= transition_856_symbol_out;
  transition_856 : transition
    port map(
      preds      => transition_856_preds,
      symbol_out => transition_856_symbol_out,
      symbol_in  => true);

  transition_857_preds(0) <= place_860_token;
  transition_857 : transition
    port map(
      preds      => transition_857_preds,
      symbol_out => transition_857_symbol_out,
      symbol_in  => LambdaIn(229));

  transition_858_preds(0) <= place_861_token;
  LambdaOut(230) <= transition_858_symbol_out;
  transition_858 : transition
    port map(
      preds      => transition_858_preds,
      symbol_out => transition_858_symbol_out,
      symbol_in  => true);

  transition_859_preds(0) <= place_862_token;
  transition_859 : transition
    port map(
      preds      => transition_859_preds,
      symbol_out => transition_859_symbol_out,
      symbol_in  => LambdaIn(230));

  transition_863_preds(0) <= place_1433_token;
  LambdaOut(231) <= transition_863_symbol_out;
  transition_863 : transition
    port map(
      preds      => transition_863_preds,
      symbol_out => transition_863_symbol_out,
      symbol_in  => true);

  transition_864_preds(0) <= place_867_token;
  transition_864 : transition
    port map(
      preds      => transition_864_preds,
      symbol_out => transition_864_symbol_out,
      symbol_in  => LambdaIn(231));

  transition_865_preds(0) <= place_868_token;
  LambdaOut(232) <= transition_865_symbol_out;
  transition_865 : transition
    port map(
      preds      => transition_865_preds,
      symbol_out => transition_865_symbol_out,
      symbol_in  => true);

  transition_866_preds(0) <= place_869_token;
  transition_866 : transition
    port map(
      preds      => transition_866_preds,
      symbol_out => transition_866_symbol_out,
      symbol_in  => LambdaIn(232));

  transition_870_preds(0) <= place_1429_token;
  transition_870_preds(1) <= place_1431_token;
  transition_870 : transition
    port map(
      preds      => transition_870_preds,
      symbol_out => transition_870_symbol_out,
      symbol_in  => true);

  transition_871_preds(0) <= place_1437_token;
  LambdaOut(233) <= transition_871_symbol_out;
  transition_871 : transition
    port map(
      preds      => transition_871_preds,
      symbol_out => transition_871_symbol_out,
      symbol_in  => true);

  transition_872_preds(0) <= place_875_token;
  transition_872 : transition
    port map(
      preds      => transition_872_preds,
      symbol_out => transition_872_symbol_out,
      symbol_in  => LambdaIn(233));

  transition_873_preds(0) <= place_876_token;
  LambdaOut(234) <= transition_873_symbol_out;
  transition_873 : transition
    port map(
      preds      => transition_873_preds,
      symbol_out => transition_873_symbol_out,
      symbol_in  => true);

  transition_874_preds(0) <= place_877_token;
  transition_874 : transition
    port map(
      preds      => transition_874_preds,
      symbol_out => transition_874_symbol_out,
      symbol_in  => LambdaIn(234));

  transition_878_preds(0) <= place_1438_token;
  LambdaOut(235) <= transition_878_symbol_out;
  transition_878 : transition
    port map(
      preds      => transition_878_preds,
      symbol_out => transition_878_symbol_out,
      symbol_in  => true);

  transition_879_preds(0) <= place_882_token;
  transition_879 : transition
    port map(
      preds      => transition_879_preds,
      symbol_out => transition_879_symbol_out,
      symbol_in  => LambdaIn(235));

  transition_880_preds(0) <= place_883_token;
  LambdaOut(236) <= transition_880_symbol_out;
  transition_880 : transition
    port map(
      preds      => transition_880_preds,
      symbol_out => transition_880_symbol_out,
      symbol_in  => true);

  transition_881_preds(0) <= place_884_token;
  transition_881 : transition
    port map(
      preds      => transition_881_preds,
      symbol_out => transition_881_symbol_out,
      symbol_in  => LambdaIn(236));

  transition_885_preds(0) <= place_1436_token;
  transition_885_preds(1) <= place_1434_token;
  transition_885 : transition
    port map(
      preds      => transition_885_preds,
      symbol_out => transition_885_symbol_out,
      symbol_in  => true);

  transition_886_preds(0) <= place_1439_token;
  LambdaOut(237) <= transition_886_symbol_out;
  transition_886 : transition
    port map(
      preds      => transition_886_preds,
      symbol_out => transition_886_symbol_out,
      symbol_in  => true);

  transition_887_preds(0) <= place_890_token;
  transition_887 : transition
    port map(
      preds      => transition_887_preds,
      symbol_out => transition_887_symbol_out,
      symbol_in  => LambdaIn(237));

  transition_888_preds(0) <= place_891_token;
  LambdaOut(238) <= transition_888_symbol_out;
  transition_888 : transition
    port map(
      preds      => transition_888_preds,
      symbol_out => transition_888_symbol_out,
      symbol_in  => true);

  transition_889_preds(0) <= place_892_token;
  transition_889 : transition
    port map(
      preds      => transition_889_preds,
      symbol_out => transition_889_symbol_out,
      symbol_in  => LambdaIn(238));

  transition_894_preds(0) <= place_893_token;
  transition_894 : transition
    port map(
      preds      => transition_894_preds,
      symbol_out => transition_894_symbol_out,
      symbol_in  => LambdaIn(239));

  transition_895_preds(0) <= place_1441_token;
  LambdaOut(239) <= transition_895_symbol_out;
  transition_895 : transition
    port map(
      preds      => transition_895_preds,
      symbol_out => transition_895_symbol_out,
      symbol_in  => true);

  transition_896_preds(0) <= place_1440_token;
  transition_896_preds(1) <= place_1445_token;
  transition_896 : transition
    port map(
      preds      => transition_896_preds,
      symbol_out => transition_896_symbol_out,
      symbol_in  => true);

  transition_898_preds(0) <= place_897_token;
  transition_898 : transition
    port map(
      preds      => transition_898_preds,
      symbol_out => transition_898_symbol_out,
      symbol_in  => LambdaIn(240));

  transition_899_preds(0) <= place_1442_token;
  LambdaOut(240) <= transition_899_symbol_out;
  transition_899 : transition
    port map(
      preds      => transition_899_preds,
      symbol_out => transition_899_symbol_out,
      symbol_in  => true);

  transition_900_preds(0) <= place_1447_token;
  LambdaOut(241) <= transition_900_symbol_out;
  transition_900 : transition
    port map(
      preds      => transition_900_preds,
      symbol_out => transition_900_symbol_out,
      symbol_in  => true);

  transition_901_preds(0) <= place_904_token;
  transition_901 : transition
    port map(
      preds      => transition_901_preds,
      symbol_out => transition_901_symbol_out,
      symbol_in  => LambdaIn(241));

  transition_902_preds(0) <= place_905_token;
  LambdaOut(242) <= transition_902_symbol_out;
  transition_902 : transition
    port map(
      preds      => transition_902_preds,
      symbol_out => transition_902_symbol_out,
      symbol_in  => true);

  transition_903_preds(0) <= place_906_token;
  transition_903 : transition
    port map(
      preds      => transition_903_preds,
      symbol_out => transition_903_symbol_out,
      symbol_in  => LambdaIn(242));

  transition_907_preds(0) <= place_1450_token;
  LambdaOut(243) <= transition_907_symbol_out;
  transition_907 : transition
    port map(
      preds      => transition_907_preds,
      symbol_out => transition_907_symbol_out,
      symbol_in  => true);

  transition_908_preds(0) <= place_911_token;
  transition_908 : transition
    port map(
      preds      => transition_908_preds,
      symbol_out => transition_908_symbol_out,
      symbol_in  => LambdaIn(243));

  transition_909_preds(0) <= place_912_token;
  LambdaOut(244) <= transition_909_symbol_out;
  transition_909 : transition
    port map(
      preds      => transition_909_preds,
      symbol_out => transition_909_symbol_out,
      symbol_in  => true);

  transition_910_preds(0) <= place_913_token;
  transition_910 : transition
    port map(
      preds      => transition_910_preds,
      symbol_out => transition_910_symbol_out,
      symbol_in  => LambdaIn(244));

  transition_914_preds(0) <= place_1451_token;
  LambdaOut(245) <= transition_914_symbol_out;
  transition_914 : transition
    port map(
      preds      => transition_914_preds,
      symbol_out => transition_914_symbol_out,
      symbol_in  => true);

  transition_915_preds(0) <= place_918_token;
  transition_915 : transition
    port map(
      preds      => transition_915_preds,
      symbol_out => transition_915_symbol_out,
      symbol_in  => LambdaIn(245));

  transition_916_preds(0) <= place_919_token;
  LambdaOut(246) <= transition_916_symbol_out;
  transition_916 : transition
    port map(
      preds      => transition_916_preds,
      symbol_out => transition_916_symbol_out,
      symbol_in  => true);

  transition_917_preds(0) <= place_920_token;
  transition_917 : transition
    port map(
      preds      => transition_917_preds,
      symbol_out => transition_917_symbol_out,
      symbol_in  => LambdaIn(246));

  transition_921_preds(0) <= place_1448_token;
  transition_921_preds(1) <= place_1446_token;
  transition_921 : transition
    port map(
      preds      => transition_921_preds,
      symbol_out => transition_921_symbol_out,
      symbol_in  => true);

  transition_922_preds(0) <= place_1455_token;
  LambdaOut(247) <= transition_922_symbol_out;
  transition_922 : transition
    port map(
      preds      => transition_922_preds,
      symbol_out => transition_922_symbol_out,
      symbol_in  => true);

  transition_923_preds(0) <= place_926_token;
  transition_923 : transition
    port map(
      preds      => transition_923_preds,
      symbol_out => transition_923_symbol_out,
      symbol_in  => LambdaIn(247));

  transition_924_preds(0) <= place_927_token;
  LambdaOut(248) <= transition_924_symbol_out;
  transition_924 : transition
    port map(
      preds      => transition_924_preds,
      symbol_out => transition_924_symbol_out,
      symbol_in  => true);

  transition_925_preds(0) <= place_928_token;
  transition_925 : transition
    port map(
      preds      => transition_925_preds,
      symbol_out => transition_925_symbol_out,
      symbol_in  => LambdaIn(248));

  transition_929_preds(0) <= place_1456_token;
  LambdaOut(249) <= transition_929_symbol_out;
  transition_929 : transition
    port map(
      preds      => transition_929_preds,
      symbol_out => transition_929_symbol_out,
      symbol_in  => true);

  transition_930_preds(0) <= place_933_token;
  transition_930 : transition
    port map(
      preds      => transition_930_preds,
      symbol_out => transition_930_symbol_out,
      symbol_in  => LambdaIn(249));

  transition_931_preds(0) <= place_934_token;
  LambdaOut(250) <= transition_931_symbol_out;
  transition_931 : transition
    port map(
      preds      => transition_931_preds,
      symbol_out => transition_931_symbol_out,
      symbol_in  => true);

  transition_932_preds(0) <= place_935_token;
  transition_932 : transition
    port map(
      preds      => transition_932_preds,
      symbol_out => transition_932_symbol_out,
      symbol_in  => LambdaIn(250));

  transition_936_preds(0) <= place_1452_token;
  transition_936_preds(1) <= place_1453_token;
  transition_936 : transition
    port map(
      preds      => transition_936_preds,
      symbol_out => transition_936_symbol_out,
      symbol_in  => true);

  transition_937_preds(0) <= place_1457_token;
  LambdaOut(251) <= transition_937_symbol_out;
  transition_937 : transition
    port map(
      preds      => transition_937_preds,
      symbol_out => transition_937_symbol_out,
      symbol_in  => true);

  transition_938_preds(0) <= place_941_token;
  transition_938 : transition
    port map(
      preds      => transition_938_preds,
      symbol_out => transition_938_symbol_out,
      symbol_in  => LambdaIn(251));

  transition_939_preds(0) <= place_942_token;
  LambdaOut(252) <= transition_939_symbol_out;
  transition_939 : transition
    port map(
      preds      => transition_939_preds,
      symbol_out => transition_939_symbol_out,
      symbol_in  => true);

  transition_940_preds(0) <= place_943_token;
  transition_940 : transition
    port map(
      preds      => transition_940_preds,
      symbol_out => transition_940_symbol_out,
      symbol_in  => LambdaIn(252));

  transition_945_preds(0) <= place_944_token;
  transition_945 : transition
    port map(
      preds      => transition_945_preds,
      symbol_out => transition_945_symbol_out,
      symbol_in  => LambdaIn(253));

  transition_946_preds(0) <= place_1459_token;
  LambdaOut(253) <= transition_946_symbol_out;
  transition_946 : transition
    port map(
      preds      => transition_946_preds,
      symbol_out => transition_946_symbol_out,
      symbol_in  => true);

  transition_947_preds(0) <= place_1458_token;
  transition_947_preds(1) <= place_1462_token;
  transition_947 : transition
    port map(
      preds      => transition_947_preds,
      symbol_out => transition_947_symbol_out,
      symbol_in  => true);

  transition_949_preds(0) <= place_948_token;
  transition_949 : transition
    port map(
      preds      => transition_949_preds,
      symbol_out => transition_949_symbol_out,
      symbol_in  => LambdaIn(254));

  transition_950_preds(0) <= place_1460_token;
  LambdaOut(254) <= transition_950_symbol_out;
  transition_950 : transition
    port map(
      preds      => transition_950_preds,
      symbol_out => transition_950_symbol_out,
      symbol_in  => true);

  transition_951_preds(0) <= place_1463_token;
  LambdaOut(255) <= transition_951_symbol_out;
  transition_951 : transition
    port map(
      preds      => transition_951_preds,
      symbol_out => transition_951_symbol_out,
      symbol_in  => true);

  transition_952_preds(0) <= place_955_token;
  transition_952 : transition
    port map(
      preds      => transition_952_preds,
      symbol_out => transition_952_symbol_out,
      symbol_in  => LambdaIn(255));

  transition_953_preds(0) <= place_956_token;
  LambdaOut(256) <= transition_953_symbol_out;
  transition_953 : transition
    port map(
      preds      => transition_953_preds,
      symbol_out => transition_953_symbol_out,
      symbol_in  => true);

  transition_954_preds(0) <= place_957_token;
  transition_954 : transition
    port map(
      preds      => transition_954_preds,
      symbol_out => transition_954_symbol_out,
      symbol_in  => LambdaIn(256));

  transition_958_preds(0) <= place_1443_token;
  transition_958_preds(1) <= place_1461_token;
  transition_958 : transition
    port map(
      preds      => transition_958_preds,
      symbol_out => transition_958_symbol_out,
      symbol_in  => true);

  transition_959_preds(0) <= place_1464_token;
  LambdaOut(257) <= transition_959_symbol_out;
  transition_959 : transition
    port map(
      preds      => transition_959_preds,
      symbol_out => transition_959_symbol_out,
      symbol_in  => true);

  transition_960_preds(0) <= place_963_token;
  transition_960 : transition
    port map(
      preds      => transition_960_preds,
      symbol_out => transition_960_symbol_out,
      symbol_in  => LambdaIn(257));

  transition_961_preds(0) <= place_964_token;
  LambdaOut(258) <= transition_961_symbol_out;
  transition_961 : transition
    port map(
      preds      => transition_961_preds,
      symbol_out => transition_961_symbol_out,
      symbol_in  => true);

  transition_962_preds(0) <= place_965_token;
  transition_962 : transition
    port map(
      preds      => transition_962_preds,
      symbol_out => transition_962_symbol_out,
      symbol_in  => LambdaIn(258));

  transition_966_preds(0) <= place_1467_token;
  LambdaOut(259) <= transition_966_symbol_out;
  transition_966 : transition
    port map(
      preds      => transition_966_preds,
      symbol_out => transition_966_symbol_out,
      symbol_in  => true);

  transition_967_preds(0) <= place_970_token;
  transition_967 : transition
    port map(
      preds      => transition_967_preds,
      symbol_out => transition_967_symbol_out,
      symbol_in  => LambdaIn(259));

  transition_968_preds(0) <= place_971_token;
  LambdaOut(260) <= transition_968_symbol_out;
  transition_968 : transition
    port map(
      preds      => transition_968_preds,
      symbol_out => transition_968_symbol_out,
      symbol_in  => true);

  transition_969_preds(0) <= place_972_token;
  transition_969 : transition
    port map(
      preds      => transition_969_preds,
      symbol_out => transition_969_symbol_out,
      symbol_in  => LambdaIn(260));

  transition_973_preds(0) <= place_1469_token;
  LambdaOut(261) <= transition_973_symbol_out;
  transition_973 : transition
    port map(
      preds      => transition_973_preds,
      symbol_out => transition_973_symbol_out,
      symbol_in  => true);

  transition_974_preds(0) <= place_977_token;
  transition_974 : transition
    port map(
      preds      => transition_974_preds,
      symbol_out => transition_974_symbol_out,
      symbol_in  => LambdaIn(261));

  transition_975_preds(0) <= place_978_token;
  LambdaOut(262) <= transition_975_symbol_out;
  transition_975 : transition
    port map(
      preds      => transition_975_preds,
      symbol_out => transition_975_symbol_out,
      symbol_in  => true);

  transition_976_preds(0) <= place_979_token;
  transition_976 : transition
    port map(
      preds      => transition_976_preds,
      symbol_out => transition_976_symbol_out,
      symbol_in  => LambdaIn(262));

  transition_980_preds(0) <= place_1470_token;
  LambdaOut(263) <= transition_980_symbol_out;
  transition_980 : transition
    port map(
      preds      => transition_980_preds,
      symbol_out => transition_980_symbol_out,
      symbol_in  => true);

  transition_981_preds(0) <= place_984_token;
  transition_981 : transition
    port map(
      preds      => transition_981_preds,
      symbol_out => transition_981_symbol_out,
      symbol_in  => LambdaIn(263));

  transition_982_preds(0) <= place_985_token;
  LambdaOut(264) <= transition_982_symbol_out;
  transition_982 : transition
    port map(
      preds      => transition_982_preds,
      symbol_out => transition_982_symbol_out,
      symbol_in  => true);

  transition_983_preds(0) <= place_986_token;
  transition_983 : transition
    port map(
      preds      => transition_983_preds,
      symbol_out => transition_983_symbol_out,
      symbol_in  => LambdaIn(264));

  transition_987_preds(0) <= place_1466_token;
  transition_987_preds(1) <= place_1468_token;
  transition_987 : transition
    port map(
      preds      => transition_987_preds,
      symbol_out => transition_987_symbol_out,
      symbol_in  => true);

  transition_988_preds(0) <= place_1473_token;
  LambdaOut(265) <= transition_988_symbol_out;
  transition_988 : transition
    port map(
      preds      => transition_988_preds,
      symbol_out => transition_988_symbol_out,
      symbol_in  => true);

  transition_989_preds(0) <= place_992_token;
  transition_989 : transition
    port map(
      preds      => transition_989_preds,
      symbol_out => transition_989_symbol_out,
      symbol_in  => LambdaIn(265));

  transition_990_preds(0) <= place_993_token;
  LambdaOut(266) <= transition_990_symbol_out;
  transition_990 : transition
    port map(
      preds      => transition_990_preds,
      symbol_out => transition_990_symbol_out,
      symbol_in  => true);

  transition_991_preds(0) <= place_994_token;
  transition_991 : transition
    port map(
      preds      => transition_991_preds,
      symbol_out => transition_991_symbol_out,
      symbol_in  => LambdaIn(266));

  transition_995_preds(0) <= place_1474_token;
  LambdaOut(267) <= transition_995_symbol_out;
  transition_995 : transition
    port map(
      preds      => transition_995_preds,
      symbol_out => transition_995_symbol_out,
      symbol_in  => true);

  transition_996_preds(0) <= place_999_token;
  transition_996 : transition
    port map(
      preds      => transition_996_preds,
      symbol_out => transition_996_symbol_out,
      symbol_in  => LambdaIn(267));

  transition_997_preds(0) <= place_1000_token;
  LambdaOut(268) <= transition_997_symbol_out;
  transition_997 : transition
    port map(
      preds      => transition_997_preds,
      symbol_out => transition_997_symbol_out,
      symbol_in  => true);

  transition_998_preds(0) <= place_1001_token;
  transition_998 : transition
    port map(
      preds      => transition_998_preds,
      symbol_out => transition_998_symbol_out,
      symbol_in  => LambdaIn(268));

  transition_1002_preds(0) <= place_1471_token;
  transition_1002_preds(1) <= place_1472_token;
  transition_1002 : transition
    port map(
      preds      => transition_1002_preds,
      symbol_out => transition_1002_symbol_out,
      symbol_in  => true);

  transition_1003_preds(0) <= place_1475_token;
  LambdaOut(269) <= transition_1003_symbol_out;
  transition_1003 : transition
    port map(
      preds      => transition_1003_preds,
      symbol_out => transition_1003_symbol_out,
      symbol_in  => true);

  transition_1004_preds(0) <= place_1007_token;
  transition_1004 : transition
    port map(
      preds      => transition_1004_preds,
      symbol_out => transition_1004_symbol_out,
      symbol_in  => LambdaIn(269));

  transition_1005_preds(0) <= place_1008_token;
  LambdaOut(270) <= transition_1005_symbol_out;
  transition_1005 : transition
    port map(
      preds      => transition_1005_preds,
      symbol_out => transition_1005_symbol_out,
      symbol_in  => true);

  transition_1006_preds(0) <= place_1009_token;
  transition_1006 : transition
    port map(
      preds      => transition_1006_preds,
      symbol_out => transition_1006_symbol_out,
      symbol_in  => LambdaIn(270));

  transition_1011_preds(0) <= place_1010_token;
  transition_1011 : transition
    port map(
      preds      => transition_1011_preds,
      symbol_out => transition_1011_symbol_out,
      symbol_in  => LambdaIn(271));

  transition_1012_preds(0) <= place_1478_token;
  LambdaOut(271) <= transition_1012_symbol_out;
  transition_1012 : transition
    port map(
      preds      => transition_1012_preds,
      symbol_out => transition_1012_symbol_out,
      symbol_in  => true);

  transition_1013_preds(0) <= place_1465_token;
  transition_1013_preds(1) <= place_1477_token;
  transition_1013 : transition
    port map(
      preds      => transition_1013_preds,
      symbol_out => transition_1013_symbol_out,
      symbol_in  => true);

  transition_1014_preds(0) <= place_1479_token;
  transition_1014 : transition
    port map(
      preds      => transition_1014_preds,
      symbol_out => transition_1014_symbol_out,
      symbol_in  => true);

  transition_1015_preds(0) <= place_1481_token;
  LambdaOut(272) <= transition_1015_symbol_out;
  transition_1015 : transition
    port map(
      preds      => transition_1015_preds,
      symbol_out => transition_1015_symbol_out,
      symbol_in  => true);

  transition_1016_preds(0) <= place_1019_token;
  transition_1016 : transition
    port map(
      preds      => transition_1016_preds,
      symbol_out => transition_1016_symbol_out,
      symbol_in  => LambdaIn(272));

  transition_1017_preds(0) <= place_1020_token;
  LambdaOut(273) <= transition_1017_symbol_out;
  transition_1017 : transition
    port map(
      preds      => transition_1017_preds,
      symbol_out => transition_1017_symbol_out,
      symbol_in  => true);

  transition_1018_preds(0) <= place_1021_token;
  transition_1018 : transition
    port map(
      preds      => transition_1018_preds,
      symbol_out => transition_1018_symbol_out,
      symbol_in  => LambdaIn(273));

  transition_1022_preds(0) <= place_1483_token;
  LambdaOut(274) <= transition_1022_symbol_out;
  transition_1022 : transition
    port map(
      preds      => transition_1022_preds,
      symbol_out => transition_1022_symbol_out,
      symbol_in  => true);

  transition_1023_preds(0) <= place_1026_token;
  transition_1023 : transition
    port map(
      preds      => transition_1023_preds,
      symbol_out => transition_1023_symbol_out,
      symbol_in  => LambdaIn(274));

  transition_1024_preds(0) <= place_1027_token;
  LambdaOut(275) <= transition_1024_symbol_out;
  transition_1024 : transition
    port map(
      preds      => transition_1024_preds,
      symbol_out => transition_1024_symbol_out,
      symbol_in  => true);

  transition_1025_preds(0) <= place_1028_token;
  transition_1025 : transition
    port map(
      preds      => transition_1025_preds,
      symbol_out => transition_1025_symbol_out,
      symbol_in  => LambdaIn(275));

  transition_1029_preds(0) <= place_1484_token;
  LambdaOut(276) <= transition_1029_symbol_out;
  transition_1029 : transition
    port map(
      preds      => transition_1029_preds,
      symbol_out => transition_1029_symbol_out,
      symbol_in  => true);

  transition_1030_preds(0) <= place_1033_token;
  transition_1030 : transition
    port map(
      preds      => transition_1030_preds,
      symbol_out => transition_1030_symbol_out,
      symbol_in  => LambdaIn(276));

  transition_1031_preds(0) <= place_1034_token;
  LambdaOut(277) <= transition_1031_symbol_out;
  transition_1031 : transition
    port map(
      preds      => transition_1031_preds,
      symbol_out => transition_1031_symbol_out,
      symbol_in  => true);

  transition_1032_preds(0) <= place_1035_token;
  transition_1032 : transition
    port map(
      preds      => transition_1032_preds,
      symbol_out => transition_1032_symbol_out,
      symbol_in  => LambdaIn(277));

  transition_1036_preds(0) <= place_1480_token;
  transition_1036_preds(1) <= place_1482_token;
  transition_1036 : transition
    port map(
      preds      => transition_1036_preds,
      symbol_out => transition_1036_symbol_out,
      symbol_in  => true);

  transition_1037_preds(0) <= place_1487_token;
  LambdaOut(278) <= transition_1037_symbol_out;
  transition_1037 : transition
    port map(
      preds      => transition_1037_preds,
      symbol_out => transition_1037_symbol_out,
      symbol_in  => true);

  transition_1038_preds(0) <= place_1041_token;
  transition_1038 : transition
    port map(
      preds      => transition_1038_preds,
      symbol_out => transition_1038_symbol_out,
      symbol_in  => LambdaIn(278));

  transition_1039_preds(0) <= place_1042_token;
  LambdaOut(279) <= transition_1039_symbol_out;
  transition_1039 : transition
    port map(
      preds      => transition_1039_preds,
      symbol_out => transition_1039_symbol_out,
      symbol_in  => true);

  transition_1040_preds(0) <= place_1043_token;
  transition_1040 : transition
    port map(
      preds      => transition_1040_preds,
      symbol_out => transition_1040_symbol_out,
      symbol_in  => LambdaIn(279));

  transition_1044_preds(0) <= place_1488_token;
  LambdaOut(280) <= transition_1044_symbol_out;
  transition_1044 : transition
    port map(
      preds      => transition_1044_preds,
      symbol_out => transition_1044_symbol_out,
      symbol_in  => true);

  transition_1045_preds(0) <= place_1048_token;
  transition_1045 : transition
    port map(
      preds      => transition_1045_preds,
      symbol_out => transition_1045_symbol_out,
      symbol_in  => LambdaIn(280));

  transition_1046_preds(0) <= place_1049_token;
  LambdaOut(281) <= transition_1046_symbol_out;
  transition_1046 : transition
    port map(
      preds      => transition_1046_preds,
      symbol_out => transition_1046_symbol_out,
      symbol_in  => true);

  transition_1047_preds(0) <= place_1050_token;
  transition_1047 : transition
    port map(
      preds      => transition_1047_preds,
      symbol_out => transition_1047_symbol_out,
      symbol_in  => LambdaIn(281));

  transition_1051_preds(0) <= place_1485_token;
  transition_1051_preds(1) <= place_1486_token;
  transition_1051 : transition
    port map(
      preds      => transition_1051_preds,
      symbol_out => transition_1051_symbol_out,
      symbol_in  => true);

  transition_1052_preds(0) <= place_1489_token;
  LambdaOut(282) <= transition_1052_symbol_out;
  transition_1052 : transition
    port map(
      preds      => transition_1052_preds,
      symbol_out => transition_1052_symbol_out,
      symbol_in  => true);

  transition_1053_preds(0) <= place_1056_token;
  transition_1053 : transition
    port map(
      preds      => transition_1053_preds,
      symbol_out => transition_1053_symbol_out,
      symbol_in  => LambdaIn(282));

  transition_1054_preds(0) <= place_1057_token;
  LambdaOut(283) <= transition_1054_symbol_out;
  transition_1054 : transition
    port map(
      preds      => transition_1054_preds,
      symbol_out => transition_1054_symbol_out,
      symbol_in  => true);

  transition_1055_preds(0) <= place_1058_token;
  transition_1055 : transition
    port map(
      preds      => transition_1055_preds,
      symbol_out => transition_1055_symbol_out,
      symbol_in  => LambdaIn(283));

  transition_1060_preds(0) <= place_1059_token;
  transition_1060 : transition
    port map(
      preds      => transition_1060_preds,
      symbol_out => transition_1060_symbol_out,
      symbol_in  => LambdaIn(284));

  transition_1061_preds(0) <= place_1492_token;
  LambdaOut(284) <= transition_1061_symbol_out;
  transition_1061 : transition
    port map(
      preds      => transition_1061_preds,
      symbol_out => transition_1061_symbol_out,
      symbol_in  => true);

  transition_1062_preds(0) <= place_1491_token;
  transition_1062_preds(1) <= place_1496_token;
  transition_1062 : transition
    port map(
      preds      => transition_1062_preds,
      symbol_out => transition_1062_symbol_out,
      symbol_in  => true);

  transition_1064_preds(0) <= place_1063_token;
  transition_1064 : transition
    port map(
      preds      => transition_1064_preds,
      symbol_out => transition_1064_symbol_out,
      symbol_in  => LambdaIn(285));

  transition_1065_preds(0) <= place_1493_token;
  LambdaOut(285) <= transition_1065_symbol_out;
  transition_1065 : transition
    port map(
      preds      => transition_1065_preds,
      symbol_out => transition_1065_symbol_out,
      symbol_in  => true);

  transition_1066_preds(0) <= place_1498_token;
  LambdaOut(286) <= transition_1066_symbol_out;
  transition_1066 : transition
    port map(
      preds      => transition_1066_preds,
      symbol_out => transition_1066_symbol_out,
      symbol_in  => true);

  transition_1067_preds(0) <= place_1070_token;
  transition_1067 : transition
    port map(
      preds      => transition_1067_preds,
      symbol_out => transition_1067_symbol_out,
      symbol_in  => LambdaIn(286));

  transition_1068_preds(0) <= place_1071_token;
  LambdaOut(287) <= transition_1068_symbol_out;
  transition_1068 : transition
    port map(
      preds      => transition_1068_preds,
      symbol_out => transition_1068_symbol_out,
      symbol_in  => true);

  transition_1069_preds(0) <= place_1072_token;
  transition_1069 : transition
    port map(
      preds      => transition_1069_preds,
      symbol_out => transition_1069_symbol_out,
      symbol_in  => LambdaIn(287));

  transition_1073_preds(0) <= place_1500_token;
  LambdaOut(288) <= transition_1073_symbol_out;
  transition_1073 : transition
    port map(
      preds      => transition_1073_preds,
      symbol_out => transition_1073_symbol_out,
      symbol_in  => true);

  transition_1074_preds(0) <= place_1077_token;
  transition_1074 : transition
    port map(
      preds      => transition_1074_preds,
      symbol_out => transition_1074_symbol_out,
      symbol_in  => LambdaIn(288));

  transition_1075_preds(0) <= place_1078_token;
  LambdaOut(289) <= transition_1075_symbol_out;
  transition_1075 : transition
    port map(
      preds      => transition_1075_preds,
      symbol_out => transition_1075_symbol_out,
      symbol_in  => true);

  transition_1076_preds(0) <= place_1079_token;
  transition_1076 : transition
    port map(
      preds      => transition_1076_preds,
      symbol_out => transition_1076_symbol_out,
      symbol_in  => LambdaIn(289));

  transition_1080_preds(0) <= place_1502_token;
  LambdaOut(290) <= transition_1080_symbol_out;
  transition_1080 : transition
    port map(
      preds      => transition_1080_preds,
      symbol_out => transition_1080_symbol_out,
      symbol_in  => true);

  transition_1081_preds(0) <= place_1084_token;
  transition_1081 : transition
    port map(
      preds      => transition_1081_preds,
      symbol_out => transition_1081_symbol_out,
      symbol_in  => LambdaIn(290));

  transition_1082_preds(0) <= place_1085_token;
  LambdaOut(291) <= transition_1082_symbol_out;
  transition_1082 : transition
    port map(
      preds      => transition_1082_preds,
      symbol_out => transition_1082_symbol_out,
      symbol_in  => true);

  transition_1083_preds(0) <= place_1086_token;
  transition_1083 : transition
    port map(
      preds      => transition_1083_preds,
      symbol_out => transition_1083_symbol_out,
      symbol_in  => LambdaIn(291));

  transition_1087_preds(0) <= place_1497_token;
  transition_1087_preds(1) <= place_1499_token;
  transition_1087 : transition
    port map(
      preds      => transition_1087_preds,
      symbol_out => transition_1087_symbol_out,
      symbol_in  => true);

  transition_1088_preds(0) <= place_1505_token;
  LambdaOut(292) <= transition_1088_symbol_out;
  transition_1088 : transition
    port map(
      preds      => transition_1088_preds,
      symbol_out => transition_1088_symbol_out,
      symbol_in  => true);

  transition_1089_preds(0) <= place_1092_token;
  transition_1089 : transition
    port map(
      preds      => transition_1089_preds,
      symbol_out => transition_1089_symbol_out,
      symbol_in  => LambdaIn(292));

  transition_1090_preds(0) <= place_1093_token;
  LambdaOut(293) <= transition_1090_symbol_out;
  transition_1090 : transition
    port map(
      preds      => transition_1090_preds,
      symbol_out => transition_1090_symbol_out,
      symbol_in  => true);

  transition_1091_preds(0) <= place_1094_token;
  transition_1091 : transition
    port map(
      preds      => transition_1091_preds,
      symbol_out => transition_1091_symbol_out,
      symbol_in  => LambdaIn(293));

  transition_1095_preds(0) <= place_1506_token;
  LambdaOut(294) <= transition_1095_symbol_out;
  transition_1095 : transition
    port map(
      preds      => transition_1095_preds,
      symbol_out => transition_1095_symbol_out,
      symbol_in  => true);

  transition_1096_preds(0) <= place_1099_token;
  transition_1096 : transition
    port map(
      preds      => transition_1096_preds,
      symbol_out => transition_1096_symbol_out,
      symbol_in  => LambdaIn(294));

  transition_1097_preds(0) <= place_1100_token;
  LambdaOut(295) <= transition_1097_symbol_out;
  transition_1097 : transition
    port map(
      preds      => transition_1097_preds,
      symbol_out => transition_1097_symbol_out,
      symbol_in  => true);

  transition_1098_preds(0) <= place_1101_token;
  transition_1098 : transition
    port map(
      preds      => transition_1098_preds,
      symbol_out => transition_1098_symbol_out,
      symbol_in  => LambdaIn(295));

  transition_1102_preds(0) <= place_1503_token;
  transition_1102_preds(1) <= place_1504_token;
  transition_1102 : transition
    port map(
      preds      => transition_1102_preds,
      symbol_out => transition_1102_symbol_out,
      symbol_in  => true);

  transition_1103_preds(0) <= place_1508_token;
  LambdaOut(296) <= transition_1103_symbol_out;
  transition_1103 : transition
    port map(
      preds      => transition_1103_preds,
      symbol_out => transition_1103_symbol_out,
      symbol_in  => true);

  transition_1104_preds(0) <= place_1107_token;
  transition_1104 : transition
    port map(
      preds      => transition_1104_preds,
      symbol_out => transition_1104_symbol_out,
      symbol_in  => LambdaIn(296));

  transition_1105_preds(0) <= place_1108_token;
  LambdaOut(297) <= transition_1105_symbol_out;
  transition_1105 : transition
    port map(
      preds      => transition_1105_preds,
      symbol_out => transition_1105_symbol_out,
      symbol_in  => true);

  transition_1106_preds(0) <= place_1109_token;
  transition_1106 : transition
    port map(
      preds      => transition_1106_preds,
      symbol_out => transition_1106_symbol_out,
      symbol_in  => LambdaIn(297));

  transition_1111_preds(0) <= place_1110_token;
  transition_1111 : transition
    port map(
      preds      => transition_1111_preds,
      symbol_out => transition_1111_symbol_out,
      symbol_in  => LambdaIn(298));

  transition_1112_preds(0) <= place_1510_token;
  LambdaOut(298) <= transition_1112_symbol_out;
  transition_1112 : transition
    port map(
      preds      => transition_1112_preds,
      symbol_out => transition_1112_symbol_out,
      symbol_in  => true);

  transition_1113_preds(0) <= place_1509_token;
  transition_1113_preds(1) <= place_1513_token;
  transition_1113 : transition
    port map(
      preds      => transition_1113_preds,
      symbol_out => transition_1113_symbol_out,
      symbol_in  => true);

  transition_1115_preds(0) <= place_1114_token;
  transition_1115 : transition
    port map(
      preds      => transition_1115_preds,
      symbol_out => transition_1115_symbol_out,
      symbol_in  => LambdaIn(299));

  transition_1116_preds(0) <= place_1511_token;
  LambdaOut(299) <= transition_1116_symbol_out;
  transition_1116 : transition
    port map(
      preds      => transition_1116_preds,
      symbol_out => transition_1116_symbol_out,
      symbol_in  => true);

  transition_1117_preds(0) <= place_1514_token;
  LambdaOut(300) <= transition_1117_symbol_out;
  transition_1117 : transition
    port map(
      preds      => transition_1117_preds,
      symbol_out => transition_1117_symbol_out,
      symbol_in  => true);

  transition_1118_preds(0) <= place_1121_token;
  transition_1118 : transition
    port map(
      preds      => transition_1118_preds,
      symbol_out => transition_1118_symbol_out,
      symbol_in  => LambdaIn(300));

  transition_1119_preds(0) <= place_1122_token;
  LambdaOut(301) <= transition_1119_symbol_out;
  transition_1119 : transition
    port map(
      preds      => transition_1119_preds,
      symbol_out => transition_1119_symbol_out,
      symbol_in  => true);

  transition_1120_preds(0) <= place_1123_token;
  transition_1120 : transition
    port map(
      preds      => transition_1120_preds,
      symbol_out => transition_1120_symbol_out,
      symbol_in  => LambdaIn(301));

  transition_1124_preds(0) <= place_1494_token;
  transition_1124_preds(1) <= place_1512_token;
  transition_1124 : transition
    port map(
      preds      => transition_1124_preds,
      symbol_out => transition_1124_symbol_out,
      symbol_in  => true);

  transition_1125_preds(0) <= place_1515_token;
  LambdaOut(302) <= transition_1125_symbol_out;
  transition_1125 : transition
    port map(
      preds      => transition_1125_preds,
      symbol_out => transition_1125_symbol_out,
      symbol_in  => true);

  transition_1126_preds(0) <= place_1129_token;
  transition_1126 : transition
    port map(
      preds      => transition_1126_preds,
      symbol_out => transition_1126_symbol_out,
      symbol_in  => LambdaIn(302));

  transition_1127_preds(0) <= place_1130_token;
  LambdaOut(303) <= transition_1127_symbol_out;
  transition_1127 : transition
    port map(
      preds      => transition_1127_preds,
      symbol_out => transition_1127_symbol_out,
      symbol_in  => true);

  transition_1128_preds(0) <= place_1131_token;
  transition_1128 : transition
    port map(
      preds      => transition_1128_preds,
      symbol_out => transition_1128_symbol_out,
      symbol_in  => LambdaIn(303));

  transition_1132_preds(0) <= place_1518_token;
  LambdaOut(304) <= transition_1132_symbol_out;
  transition_1132 : transition
    port map(
      preds      => transition_1132_preds,
      symbol_out => transition_1132_symbol_out,
      symbol_in  => true);

  transition_1133_preds(0) <= place_1136_token;
  transition_1133 : transition
    port map(
      preds      => transition_1133_preds,
      symbol_out => transition_1133_symbol_out,
      symbol_in  => LambdaIn(304));

  transition_1134_preds(0) <= place_1137_token;
  LambdaOut(305) <= transition_1134_symbol_out;
  transition_1134 : transition
    port map(
      preds      => transition_1134_preds,
      symbol_out => transition_1134_symbol_out,
      symbol_in  => true);

  transition_1135_preds(0) <= place_1138_token;
  transition_1135 : transition
    port map(
      preds      => transition_1135_preds,
      symbol_out => transition_1135_symbol_out,
      symbol_in  => LambdaIn(305));

  transition_1139_preds(0) <= place_1520_token;
  LambdaOut(306) <= transition_1139_symbol_out;
  transition_1139 : transition
    port map(
      preds      => transition_1139_preds,
      symbol_out => transition_1139_symbol_out,
      symbol_in  => true);

  transition_1140_preds(0) <= place_1143_token;
  transition_1140 : transition
    port map(
      preds      => transition_1140_preds,
      symbol_out => transition_1140_symbol_out,
      symbol_in  => LambdaIn(306));

  transition_1141_preds(0) <= place_1144_token;
  LambdaOut(307) <= transition_1141_symbol_out;
  transition_1141 : transition
    port map(
      preds      => transition_1141_preds,
      symbol_out => transition_1141_symbol_out,
      symbol_in  => true);

  transition_1142_preds(0) <= place_1145_token;
  transition_1142 : transition
    port map(
      preds      => transition_1142_preds,
      symbol_out => transition_1142_symbol_out,
      symbol_in  => LambdaIn(307));

  transition_1146_preds(0) <= place_1521_token;
  LambdaOut(308) <= transition_1146_symbol_out;
  transition_1146 : transition
    port map(
      preds      => transition_1146_preds,
      symbol_out => transition_1146_symbol_out,
      symbol_in  => true);

  transition_1147_preds(0) <= place_1150_token;
  transition_1147 : transition
    port map(
      preds      => transition_1147_preds,
      symbol_out => transition_1147_symbol_out,
      symbol_in  => LambdaIn(308));

  transition_1148_preds(0) <= place_1151_token;
  LambdaOut(309) <= transition_1148_symbol_out;
  transition_1148 : transition
    port map(
      preds      => transition_1148_preds,
      symbol_out => transition_1148_symbol_out,
      symbol_in  => true);

  transition_1149_preds(0) <= place_1152_token;
  transition_1149 : transition
    port map(
      preds      => transition_1149_preds,
      symbol_out => transition_1149_symbol_out,
      symbol_in  => LambdaIn(309));

  transition_1153_preds(0) <= place_1519_token;
  transition_1153_preds(1) <= place_1517_token;
  transition_1153 : transition
    port map(
      preds      => transition_1153_preds,
      symbol_out => transition_1153_symbol_out,
      symbol_in  => true);

  transition_1154_preds(0) <= place_1525_token;
  LambdaOut(310) <= transition_1154_symbol_out;
  transition_1154 : transition
    port map(
      preds      => transition_1154_preds,
      symbol_out => transition_1154_symbol_out,
      symbol_in  => true);

  transition_1155_preds(0) <= place_1158_token;
  transition_1155 : transition
    port map(
      preds      => transition_1155_preds,
      symbol_out => transition_1155_symbol_out,
      symbol_in  => LambdaIn(310));

  transition_1156_preds(0) <= place_1159_token;
  LambdaOut(311) <= transition_1156_symbol_out;
  transition_1156 : transition
    port map(
      preds      => transition_1156_preds,
      symbol_out => transition_1156_symbol_out,
      symbol_in  => true);

  transition_1157_preds(0) <= place_1160_token;
  transition_1157 : transition
    port map(
      preds      => transition_1157_preds,
      symbol_out => transition_1157_symbol_out,
      symbol_in  => LambdaIn(311));

  transition_1161_preds(0) <= place_1526_token;
  LambdaOut(312) <= transition_1161_symbol_out;
  transition_1161 : transition
    port map(
      preds      => transition_1161_preds,
      symbol_out => transition_1161_symbol_out,
      symbol_in  => true);

  transition_1162_preds(0) <= place_1165_token;
  transition_1162 : transition
    port map(
      preds      => transition_1162_preds,
      symbol_out => transition_1162_symbol_out,
      symbol_in  => LambdaIn(312));

  transition_1163_preds(0) <= place_1166_token;
  LambdaOut(313) <= transition_1163_symbol_out;
  transition_1163 : transition
    port map(
      preds      => transition_1163_preds,
      symbol_out => transition_1163_symbol_out,
      symbol_in  => true);

  transition_1164_preds(0) <= place_1167_token;
  transition_1164 : transition
    port map(
      preds      => transition_1164_preds,
      symbol_out => transition_1164_symbol_out,
      symbol_in  => LambdaIn(313));

  transition_1168_preds(0) <= place_1522_token;
  transition_1168_preds(1) <= place_1523_token;
  transition_1168 : transition
    port map(
      preds      => transition_1168_preds,
      symbol_out => transition_1168_symbol_out,
      symbol_in  => true);

  transition_1169_preds(0) <= place_1527_token;
  LambdaOut(314) <= transition_1169_symbol_out;
  transition_1169 : transition
    port map(
      preds      => transition_1169_preds,
      symbol_out => transition_1169_symbol_out,
      symbol_in  => true);

  transition_1170_preds(0) <= place_1173_token;
  transition_1170 : transition
    port map(
      preds      => transition_1170_preds,
      symbol_out => transition_1170_symbol_out,
      symbol_in  => LambdaIn(314));

  transition_1171_preds(0) <= place_1174_token;
  LambdaOut(315) <= transition_1171_symbol_out;
  transition_1171 : transition
    port map(
      preds      => transition_1171_preds,
      symbol_out => transition_1171_symbol_out,
      symbol_in  => true);

  transition_1172_preds(0) <= place_1175_token;
  transition_1172 : transition
    port map(
      preds      => transition_1172_preds,
      symbol_out => transition_1172_symbol_out,
      symbol_in  => LambdaIn(315));

  transition_1177_preds(0) <= place_1176_token;
  transition_1177 : transition
    port map(
      preds      => transition_1177_preds,
      symbol_out => transition_1177_symbol_out,
      symbol_in  => LambdaIn(316));

  transition_1178_preds(0) <= place_1530_token;
  LambdaOut(316) <= transition_1178_symbol_out;
  transition_1178 : transition
    port map(
      preds      => transition_1178_preds,
      symbol_out => transition_1178_symbol_out,
      symbol_in  => true);

  transition_1179_preds(0) <= place_1516_token;
  transition_1179_preds(1) <= place_1528_token;
  transition_1179 : transition
    port map(
      preds      => transition_1179_preds,
      symbol_out => transition_1179_symbol_out,
      symbol_in  => true);

  transition_1180_preds(0) <= place_1532_token;
  LambdaOut(317) <= transition_1180_symbol_out;
  transition_1180 : transition
    port map(
      preds      => transition_1180_preds,
      symbol_out => transition_1180_symbol_out,
      symbol_in  => true);

  transition_1181_preds(0) <= place_1184_token;
  transition_1181 : transition
    port map(
      preds      => transition_1181_preds,
      symbol_out => transition_1181_symbol_out,
      symbol_in  => LambdaIn(317));

  transition_1182_preds(0) <= place_1185_token;
  LambdaOut(318) <= transition_1182_symbol_out;
  transition_1182 : transition
    port map(
      preds      => transition_1182_preds,
      symbol_out => transition_1182_symbol_out,
      symbol_in  => true);

  transition_1183_preds(0) <= place_1186_token;
  transition_1183 : transition
    port map(
      preds      => transition_1183_preds,
      symbol_out => transition_1183_symbol_out,
      symbol_in  => LambdaIn(318));

  transition_1187_preds(0) <= place_1534_token;
  transition_1187_preds(1) <= place_1535_token;
  transition_1187 : transition
    port map(
      preds      => transition_1187_preds,
      symbol_out => transition_1187_symbol_out,
      symbol_in  => true);

  transition_1188_preds(0) <= place_1537_token;
  LambdaOut(319) <= transition_1188_symbol_out;
  transition_1188 : transition
    port map(
      preds      => transition_1188_preds,
      symbol_out => transition_1188_symbol_out,
      symbol_in  => true);

  transition_1189_preds(0) <= place_1192_token;
  transition_1189 : transition
    port map(
      preds      => transition_1189_preds,
      symbol_out => transition_1189_symbol_out,
      symbol_in  => LambdaIn(319));

  transition_1190_preds(0) <= place_1193_token;
  LambdaOut(320) <= transition_1190_symbol_out;
  transition_1190 : transition
    port map(
      preds      => transition_1190_preds,
      symbol_out => transition_1190_symbol_out,
      symbol_in  => true);

  transition_1191_preds(0) <= place_1194_token;
  transition_1191 : transition
    port map(
      preds      => transition_1191_preds,
      symbol_out => transition_1191_symbol_out,
      symbol_in  => LambdaIn(320));

  transition_1195_preds(0) <= place_1533_token;
  transition_1195_preds(1) <= place_1539_token;
  transition_1195 : transition
    port map(
      preds      => transition_1195_preds,
      symbol_out => transition_1195_symbol_out,
      symbol_in  => true);

  transition_1196_preds(0) <= place_1538_token;
  LambdaOut(321) <= transition_1196_symbol_out;
  transition_1196 : transition
    port map(
      preds      => transition_1196_preds,
      symbol_out => transition_1196_symbol_out,
      symbol_in  => true);

  transition_1197_preds(0) <= place_1200_token;
  transition_1197 : transition
    port map(
      preds      => transition_1197_preds,
      symbol_out => transition_1197_symbol_out,
      symbol_in  => LambdaIn(321));

  transition_1198_preds(0) <= place_1201_token;
  LambdaOut(322) <= transition_1198_symbol_out;
  transition_1198 : transition
    port map(
      preds      => transition_1198_preds,
      symbol_out => transition_1198_symbol_out,
      symbol_in  => true);

  transition_1199_preds(0) <= place_1202_token;
  transition_1199 : transition
    port map(
      preds      => transition_1199_preds,
      symbol_out => transition_1199_symbol_out,
      symbol_in  => LambdaIn(322));

  transition_1204_preds(0) <= place_1203_token;
  transition_1204 : transition
    port map(
      preds      => transition_1204_preds,
      symbol_out => transition_1204_symbol_out,
      symbol_in  => LambdaIn(323));

  transition_1205_preds(0) <= place_1541_token;
  LambdaOut(323) <= transition_1205_symbol_out;
  transition_1205 : transition
    port map(
      preds      => transition_1205_preds,
      symbol_out => transition_1205_symbol_out,
      symbol_in  => true);

end architecture default_arch;