-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant GV_15_base_address : std_logic_vector(8 downto 0) := "000000000";
  constant GV_16_base_address : std_logic_vector(4 downto 0) := "00000";
  constant ahir_heap_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant click_bc_iNtErNal_x_ZZN14LinearIPLookup4pushEiP6PacketE10complained_base_address : std_logic_vector(0 downto 0) := "0";
  constant free_queue_ram_base_address : std_logic_vector(15 downto 0) := "0000000000000000";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity GV_15_initializer_in_click_bc is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity GV_15_initializer_in_click_bc;
architecture Default of GV_15_initializer_in_click_bc is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal GV_15_initializer_in_click_bc_CP_0_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_176_gather_scatter_req_0 : boolean;
  signal array_obj_ref_176_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_241_store_0_ack_0 : boolean;
  signal array_obj_ref_241_store_0_req_1 : boolean;
  signal array_obj_ref_241_store_0_ack_1 : boolean;
  signal array_obj_ref_176_store_0_req_0 : boolean;
  signal array_obj_ref_176_store_0_ack_0 : boolean;
  signal array_obj_ref_176_store_0_req_1 : boolean;
  signal array_obj_ref_176_store_0_ack_1 : boolean;
  signal array_obj_ref_185_gather_scatter_req_0 : boolean;
  signal array_obj_ref_185_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_185_store_0_req_0 : boolean;
  signal array_obj_ref_185_store_0_ack_0 : boolean;
  signal array_obj_ref_185_store_0_req_1 : boolean;
  signal array_obj_ref_185_store_0_ack_1 : boolean;
  signal array_obj_ref_192_gather_scatter_req_0 : boolean;
  signal array_obj_ref_192_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_192_store_0_req_0 : boolean;
  signal array_obj_ref_192_store_0_ack_0 : boolean;
  signal array_obj_ref_192_store_0_req_1 : boolean;
  signal array_obj_ref_192_store_0_ack_1 : boolean;
  signal array_obj_ref_199_gather_scatter_req_0 : boolean;
  signal array_obj_ref_199_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_199_store_0_req_0 : boolean;
  signal array_obj_ref_199_store_0_ack_0 : boolean;
  signal array_obj_ref_199_store_0_req_1 : boolean;
  signal array_obj_ref_199_store_0_ack_1 : boolean;
  signal array_obj_ref_206_gather_scatter_req_0 : boolean;
  signal array_obj_ref_206_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_206_store_0_req_0 : boolean;
  signal array_obj_ref_206_store_0_ack_0 : boolean;
  signal array_obj_ref_206_store_0_req_1 : boolean;
  signal array_obj_ref_206_store_0_ack_1 : boolean;
  signal array_obj_ref_213_gather_scatter_req_0 : boolean;
  signal array_obj_ref_213_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_213_store_0_req_0 : boolean;
  signal array_obj_ref_213_store_0_ack_0 : boolean;
  signal array_obj_ref_213_store_0_req_1 : boolean;
  signal array_obj_ref_213_store_0_ack_1 : boolean;
  signal array_obj_ref_220_gather_scatter_req_0 : boolean;
  signal array_obj_ref_220_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_220_store_0_req_0 : boolean;
  signal array_obj_ref_220_store_0_ack_0 : boolean;
  signal array_obj_ref_220_store_0_req_1 : boolean;
  signal array_obj_ref_220_store_0_ack_1 : boolean;
  signal array_obj_ref_227_gather_scatter_req_0 : boolean;
  signal array_obj_ref_227_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_227_store_0_req_0 : boolean;
  signal array_obj_ref_227_store_0_ack_0 : boolean;
  signal array_obj_ref_227_store_0_req_1 : boolean;
  signal array_obj_ref_227_store_0_ack_1 : boolean;
  signal array_obj_ref_234_gather_scatter_req_0 : boolean;
  signal array_obj_ref_234_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_234_store_0_req_0 : boolean;
  signal array_obj_ref_234_store_0_ack_0 : boolean;
  signal array_obj_ref_234_store_0_req_1 : boolean;
  signal array_obj_ref_234_store_0_ack_1 : boolean;
  signal array_obj_ref_241_gather_scatter_req_0 : boolean;
  signal array_obj_ref_241_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_241_store_0_req_0 : boolean;
  signal array_obj_ref_248_gather_scatter_req_0 : boolean;
  signal array_obj_ref_248_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_248_store_0_req_0 : boolean;
  signal array_obj_ref_248_store_0_ack_0 : boolean;
  signal array_obj_ref_248_store_0_req_1 : boolean;
  signal array_obj_ref_248_store_0_ack_1 : boolean;
  signal array_obj_ref_255_gather_scatter_req_0 : boolean;
  signal array_obj_ref_255_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_255_store_0_req_0 : boolean;
  signal array_obj_ref_255_store_0_ack_0 : boolean;
  signal array_obj_ref_255_store_0_req_1 : boolean;
  signal array_obj_ref_255_store_0_ack_1 : boolean;
  signal array_obj_ref_262_gather_scatter_req_0 : boolean;
  signal array_obj_ref_262_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_262_store_0_req_0 : boolean;
  signal array_obj_ref_262_store_0_ack_0 : boolean;
  signal array_obj_ref_262_store_0_req_1 : boolean;
  signal array_obj_ref_262_store_0_ack_1 : boolean;
  signal array_obj_ref_269_gather_scatter_req_0 : boolean;
  signal array_obj_ref_269_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_269_store_0_req_0 : boolean;
  signal array_obj_ref_269_store_0_ack_0 : boolean;
  signal array_obj_ref_269_store_0_req_1 : boolean;
  signal array_obj_ref_269_store_0_ack_1 : boolean;
  signal array_obj_ref_276_gather_scatter_req_0 : boolean;
  signal array_obj_ref_276_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_0 : boolean;
  signal array_obj_ref_276_store_0_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_1 : boolean;
  signal array_obj_ref_276_store_0_ack_1 : boolean;
  signal array_obj_ref_283_gather_scatter_req_0 : boolean;
  signal array_obj_ref_283_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_283_store_0_req_0 : boolean;
  signal array_obj_ref_283_store_0_ack_0 : boolean;
  signal array_obj_ref_283_store_0_req_1 : boolean;
  signal array_obj_ref_283_store_0_ack_1 : boolean;
  signal array_obj_ref_290_gather_scatter_req_0 : boolean;
  signal array_obj_ref_290_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_290_store_0_req_0 : boolean;
  signal array_obj_ref_290_store_0_ack_0 : boolean;
  signal array_obj_ref_290_store_0_req_1 : boolean;
  signal array_obj_ref_290_store_0_ack_1 : boolean;
  signal array_obj_ref_297_gather_scatter_req_0 : boolean;
  signal array_obj_ref_297_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_297_store_0_req_0 : boolean;
  signal array_obj_ref_297_store_0_ack_0 : boolean;
  signal array_obj_ref_297_store_0_req_1 : boolean;
  signal array_obj_ref_297_store_0_ack_1 : boolean;
  signal array_obj_ref_304_gather_scatter_req_0 : boolean;
  signal array_obj_ref_304_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_304_store_0_req_0 : boolean;
  signal array_obj_ref_304_store_0_ack_0 : boolean;
  signal array_obj_ref_304_store_0_req_1 : boolean;
  signal array_obj_ref_304_store_0_ack_1 : boolean;
  signal array_obj_ref_311_gather_scatter_req_0 : boolean;
  signal array_obj_ref_311_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_311_store_0_req_0 : boolean;
  signal array_obj_ref_311_store_0_ack_0 : boolean;
  signal array_obj_ref_311_store_0_req_1 : boolean;
  signal array_obj_ref_311_store_0_ack_1 : boolean;
  signal array_obj_ref_318_gather_scatter_req_0 : boolean;
  signal array_obj_ref_318_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_0 : boolean;
  signal array_obj_ref_318_store_0_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_1 : boolean;
  signal array_obj_ref_318_store_0_ack_1 : boolean;
  signal array_obj_ref_325_gather_scatter_req_0 : boolean;
  signal array_obj_ref_325_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_325_store_0_req_0 : boolean;
  signal array_obj_ref_325_store_0_ack_0 : boolean;
  signal array_obj_ref_325_store_0_req_1 : boolean;
  signal array_obj_ref_325_store_0_ack_1 : boolean;
  signal array_obj_ref_332_gather_scatter_req_0 : boolean;
  signal array_obj_ref_332_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_332_store_0_req_0 : boolean;
  signal array_obj_ref_332_store_0_ack_0 : boolean;
  signal array_obj_ref_332_store_0_req_1 : boolean;
  signal array_obj_ref_332_store_0_ack_1 : boolean;
  signal array_obj_ref_339_gather_scatter_req_0 : boolean;
  signal array_obj_ref_339_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_339_store_0_req_0 : boolean;
  signal array_obj_ref_339_store_0_ack_0 : boolean;
  signal array_obj_ref_339_store_0_req_1 : boolean;
  signal array_obj_ref_339_store_0_ack_1 : boolean;
  signal array_obj_ref_346_gather_scatter_req_0 : boolean;
  signal array_obj_ref_346_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_0 : boolean;
  signal array_obj_ref_346_store_0_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_1 : boolean;
  signal array_obj_ref_346_store_0_ack_1 : boolean;
  signal array_obj_ref_353_gather_scatter_req_0 : boolean;
  signal array_obj_ref_353_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_353_store_0_req_0 : boolean;
  signal array_obj_ref_353_store_0_ack_0 : boolean;
  signal array_obj_ref_353_store_0_req_1 : boolean;
  signal array_obj_ref_353_store_0_ack_1 : boolean;
  signal array_obj_ref_360_gather_scatter_req_0 : boolean;
  signal array_obj_ref_360_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_360_store_0_req_0 : boolean;
  signal array_obj_ref_360_store_0_ack_0 : boolean;
  signal array_obj_ref_360_store_0_req_1 : boolean;
  signal array_obj_ref_360_store_0_ack_1 : boolean;
  signal array_obj_ref_367_gather_scatter_req_0 : boolean;
  signal array_obj_ref_367_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_367_store_0_req_0 : boolean;
  signal array_obj_ref_367_store_0_ack_0 : boolean;
  signal array_obj_ref_367_store_0_req_1 : boolean;
  signal array_obj_ref_367_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  GV_15_initializer_in_click_bc_CP_0: Block -- control-path 
    signal cp_elements: BooleanArray(84 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(84);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(84), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    split_req_12_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => array_obj_ref_176_gather_scatter_req_0); -- 
    split_ack_13_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_176_gather_scatter_ack_0, ack => cp_elements(1)); -- 
    rr_20_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => array_obj_ref_176_store_0_req_0); -- 
    ra_21_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_176_store_0_ack_0, ack => cp_elements(2)); -- 
    cr_22_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => array_obj_ref_176_store_0_req_1); -- 
    ca_23_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_176_store_0_ack_1, ack => cp_elements(3)); -- 
    split_req_33_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => array_obj_ref_185_gather_scatter_req_0); -- 
    split_ack_34_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_gather_scatter_ack_0, ack => cp_elements(4)); -- 
    rr_41_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => array_obj_ref_185_store_0_req_0); -- 
    ra_42_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_store_0_ack_0, ack => cp_elements(5)); -- 
    cr_43_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => array_obj_ref_185_store_0_req_1); -- 
    ca_44_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_store_0_ack_1, ack => cp_elements(6)); -- 
    split_req_54_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => array_obj_ref_192_gather_scatter_req_0); -- 
    split_ack_55_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_192_gather_scatter_ack_0, ack => cp_elements(7)); -- 
    rr_62_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => array_obj_ref_192_store_0_req_0); -- 
    ra_63_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_192_store_0_ack_0, ack => cp_elements(8)); -- 
    cr_64_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => array_obj_ref_192_store_0_req_1); -- 
    ca_65_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_192_store_0_ack_1, ack => cp_elements(9)); -- 
    split_req_75_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => array_obj_ref_199_gather_scatter_req_0); -- 
    split_ack_76_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_199_gather_scatter_ack_0, ack => cp_elements(10)); -- 
    rr_83_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => array_obj_ref_199_store_0_req_0); -- 
    ra_84_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_199_store_0_ack_0, ack => cp_elements(11)); -- 
    cr_85_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => array_obj_ref_199_store_0_req_1); -- 
    ca_86_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_199_store_0_ack_1, ack => cp_elements(12)); -- 
    split_req_96_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => array_obj_ref_206_gather_scatter_req_0); -- 
    split_ack_97_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_gather_scatter_ack_0, ack => cp_elements(13)); -- 
    rr_104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => array_obj_ref_206_store_0_req_0); -- 
    ra_105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_store_0_ack_0, ack => cp_elements(14)); -- 
    cr_106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => array_obj_ref_206_store_0_req_1); -- 
    ca_107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_store_0_ack_1, ack => cp_elements(15)); -- 
    split_req_117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => array_obj_ref_213_gather_scatter_req_0); -- 
    split_ack_118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_gather_scatter_ack_0, ack => cp_elements(16)); -- 
    rr_125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_213_store_0_req_0); -- 
    ra_126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_store_0_ack_0, ack => cp_elements(17)); -- 
    cr_127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => array_obj_ref_213_store_0_req_1); -- 
    ca_128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_store_0_ack_1, ack => cp_elements(18)); -- 
    split_req_138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => array_obj_ref_220_gather_scatter_req_0); -- 
    split_ack_139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_220_gather_scatter_ack_0, ack => cp_elements(19)); -- 
    rr_146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => array_obj_ref_220_store_0_req_0); -- 
    ra_147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_220_store_0_ack_0, ack => cp_elements(20)); -- 
    cr_148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => array_obj_ref_220_store_0_req_1); -- 
    ca_149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_220_store_0_ack_1, ack => cp_elements(21)); -- 
    split_req_159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_227_gather_scatter_req_0); -- 
    split_ack_160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_227_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    rr_167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_227_store_0_req_0); -- 
    ra_168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_227_store_0_ack_0, ack => cp_elements(23)); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => array_obj_ref_227_store_0_req_1); -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_227_store_0_ack_1, ack => cp_elements(24)); -- 
    split_req_180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => array_obj_ref_234_gather_scatter_req_0); -- 
    split_ack_181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_234_gather_scatter_ack_0, ack => cp_elements(25)); -- 
    rr_188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => array_obj_ref_234_store_0_req_0); -- 
    ra_189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_234_store_0_ack_0, ack => cp_elements(26)); -- 
    cr_190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => array_obj_ref_234_store_0_req_1); -- 
    ca_191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_234_store_0_ack_1, ack => cp_elements(27)); -- 
    split_req_201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => array_obj_ref_241_gather_scatter_req_0); -- 
    split_ack_202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_241_gather_scatter_ack_0, ack => cp_elements(28)); -- 
    rr_209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => array_obj_ref_241_store_0_req_0); -- 
    ra_210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_241_store_0_ack_0, ack => cp_elements(29)); -- 
    cr_211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => array_obj_ref_241_store_0_req_1); -- 
    ca_212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_241_store_0_ack_1, ack => cp_elements(30)); -- 
    split_req_222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => array_obj_ref_248_gather_scatter_req_0); -- 
    split_ack_223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_248_gather_scatter_ack_0, ack => cp_elements(31)); -- 
    rr_230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_248_store_0_req_0); -- 
    ra_231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_248_store_0_ack_0, ack => cp_elements(32)); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_248_store_0_req_1); -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_248_store_0_ack_1, ack => cp_elements(33)); -- 
    split_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_255_gather_scatter_req_0); -- 
    split_ack_244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_255_gather_scatter_ack_0, ack => cp_elements(34)); -- 
    rr_251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_255_store_0_req_0); -- 
    ra_252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_255_store_0_ack_0, ack => cp_elements(35)); -- 
    cr_253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => array_obj_ref_255_store_0_req_1); -- 
    ca_254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_255_store_0_ack_1, ack => cp_elements(36)); -- 
    split_req_264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_262_gather_scatter_req_0); -- 
    split_ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_262_gather_scatter_ack_0, ack => cp_elements(37)); -- 
    rr_272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_262_store_0_req_0); -- 
    ra_273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_262_store_0_ack_0, ack => cp_elements(38)); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_262_store_0_req_1); -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_262_store_0_ack_1, ack => cp_elements(39)); -- 
    split_req_285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => array_obj_ref_269_gather_scatter_req_0); -- 
    split_ack_286_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_gather_scatter_ack_0, ack => cp_elements(40)); -- 
    rr_293_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => array_obj_ref_269_store_0_req_0); -- 
    ra_294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_store_0_ack_0, ack => cp_elements(41)); -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => array_obj_ref_269_store_0_req_1); -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_store_0_ack_1, ack => cp_elements(42)); -- 
    split_req_306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => array_obj_ref_276_gather_scatter_req_0); -- 
    split_ack_307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_gather_scatter_ack_0, ack => cp_elements(43)); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => array_obj_ref_276_store_0_req_0); -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_store_0_ack_0, ack => cp_elements(44)); -- 
    cr_316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => array_obj_ref_276_store_0_req_1); -- 
    ca_317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_store_0_ack_1, ack => cp_elements(45)); -- 
    split_req_327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => array_obj_ref_283_gather_scatter_req_0); -- 
    split_ack_328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_gather_scatter_ack_0, ack => cp_elements(46)); -- 
    rr_335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => array_obj_ref_283_store_0_req_0); -- 
    ra_336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_store_0_ack_0, ack => cp_elements(47)); -- 
    cr_337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => array_obj_ref_283_store_0_req_1); -- 
    ca_338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_store_0_ack_1, ack => cp_elements(48)); -- 
    split_req_348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => array_obj_ref_290_gather_scatter_req_0); -- 
    split_ack_349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_290_gather_scatter_ack_0, ack => cp_elements(49)); -- 
    rr_356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => array_obj_ref_290_store_0_req_0); -- 
    ra_357_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_290_store_0_ack_0, ack => cp_elements(50)); -- 
    cr_358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => array_obj_ref_290_store_0_req_1); -- 
    ca_359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_290_store_0_ack_1, ack => cp_elements(51)); -- 
    split_req_369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_297_gather_scatter_req_0); -- 
    split_ack_370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_gather_scatter_ack_0, ack => cp_elements(52)); -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => array_obj_ref_297_store_0_req_0); -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_store_0_ack_0, ack => cp_elements(53)); -- 
    cr_379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_297_store_0_req_1); -- 
    ca_380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_store_0_ack_1, ack => cp_elements(54)); -- 
    split_req_390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => array_obj_ref_304_gather_scatter_req_0); -- 
    split_ack_391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_gather_scatter_ack_0, ack => cp_elements(55)); -- 
    rr_398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => array_obj_ref_304_store_0_req_0); -- 
    ra_399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_store_0_ack_0, ack => cp_elements(56)); -- 
    cr_400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => array_obj_ref_304_store_0_req_1); -- 
    ca_401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_store_0_ack_1, ack => cp_elements(57)); -- 
    split_req_411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => array_obj_ref_311_gather_scatter_req_0); -- 
    split_ack_412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_gather_scatter_ack_0, ack => cp_elements(58)); -- 
    rr_419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => array_obj_ref_311_store_0_req_0); -- 
    ra_420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_store_0_ack_0, ack => cp_elements(59)); -- 
    cr_421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => array_obj_ref_311_store_0_req_1); -- 
    ca_422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_store_0_ack_1, ack => cp_elements(60)); -- 
    split_req_432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => array_obj_ref_318_gather_scatter_req_0); -- 
    split_ack_433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_318_gather_scatter_ack_0, ack => cp_elements(61)); -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => array_obj_ref_318_store_0_req_0); -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_318_store_0_ack_0, ack => cp_elements(62)); -- 
    cr_442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => array_obj_ref_318_store_0_req_1); -- 
    ca_443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_318_store_0_ack_1, ack => cp_elements(63)); -- 
    split_req_453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => array_obj_ref_325_gather_scatter_req_0); -- 
    split_ack_454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_325_gather_scatter_ack_0, ack => cp_elements(64)); -- 
    rr_461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => array_obj_ref_325_store_0_req_0); -- 
    ra_462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_325_store_0_ack_0, ack => cp_elements(65)); -- 
    cr_463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => array_obj_ref_325_store_0_req_1); -- 
    ca_464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_325_store_0_ack_1, ack => cp_elements(66)); -- 
    split_req_474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => array_obj_ref_332_gather_scatter_req_0); -- 
    split_ack_475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_gather_scatter_ack_0, ack => cp_elements(67)); -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => array_obj_ref_332_store_0_req_0); -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_store_0_ack_0, ack => cp_elements(68)); -- 
    cr_484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => array_obj_ref_332_store_0_req_1); -- 
    ca_485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_store_0_ack_1, ack => cp_elements(69)); -- 
    split_req_495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_339_gather_scatter_req_0); -- 
    split_ack_496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_339_gather_scatter_ack_0, ack => cp_elements(70)); -- 
    rr_503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_339_store_0_req_0); -- 
    ra_504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_339_store_0_ack_0, ack => cp_elements(71)); -- 
    cr_505_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_339_store_0_req_1); -- 
    ca_506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_339_store_0_ack_1, ack => cp_elements(72)); -- 
    split_req_516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_346_gather_scatter_req_0); -- 
    split_ack_517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_346_gather_scatter_ack_0, ack => cp_elements(73)); -- 
    rr_524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_346_store_0_req_0); -- 
    ra_525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_346_store_0_ack_0, ack => cp_elements(74)); -- 
    cr_526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_346_store_0_req_1); -- 
    ca_527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_346_store_0_ack_1, ack => cp_elements(75)); -- 
    split_req_537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_353_gather_scatter_req_0); -- 
    split_ack_538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_353_gather_scatter_ack_0, ack => cp_elements(76)); -- 
    rr_545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => array_obj_ref_353_store_0_req_0); -- 
    ra_546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_353_store_0_ack_0, ack => cp_elements(77)); -- 
    cr_547_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => array_obj_ref_353_store_0_req_1); -- 
    ca_548_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_353_store_0_ack_1, ack => cp_elements(78)); -- 
    split_req_558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => array_obj_ref_360_gather_scatter_req_0); -- 
    split_ack_559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_360_gather_scatter_ack_0, ack => cp_elements(79)); -- 
    rr_566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => array_obj_ref_360_store_0_req_0); -- 
    ra_567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_360_store_0_ack_0, ack => cp_elements(80)); -- 
    cr_568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => array_obj_ref_360_store_0_req_1); -- 
    ca_569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_360_store_0_ack_1, ack => cp_elements(81)); -- 
    split_req_579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_367_gather_scatter_req_0); -- 
    split_ack_580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_367_gather_scatter_ack_0, ack => cp_elements(82)); -- 
    rr_587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_367_store_0_req_0); -- 
    ra_588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_367_store_0_ack_0, ack => cp_elements(83)); -- 
    cr_589_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => array_obj_ref_367_store_0_req_1); -- 
    ca_590_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_367_store_0_ack_1, ack => cp_elements(84)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_176_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_176_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_185_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_185_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_192_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_192_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_199_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_199_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_206_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_206_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_213_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_213_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_220_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_220_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_227_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_227_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_234_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_234_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_241_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_241_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_248_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_248_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_255_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_255_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_262_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_262_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_269_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_269_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_276_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_283_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_283_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_290_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_290_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_297_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_297_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_304_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_304_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_311_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_311_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_318_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_318_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_325_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_325_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_332_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_332_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_339_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_339_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_346_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_346_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_353_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_353_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_360_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_360_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_367_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_367_word_address_0 : std_logic_vector(8 downto 0);
    signal expr_177_wire_constant : std_logic_vector(7 downto 0);
    signal expr_186_wire_constant : std_logic_vector(7 downto 0);
    signal expr_193_wire_constant : std_logic_vector(7 downto 0);
    signal expr_200_wire_constant : std_logic_vector(7 downto 0);
    signal expr_207_wire_constant : std_logic_vector(7 downto 0);
    signal expr_214_wire_constant : std_logic_vector(7 downto 0);
    signal expr_221_wire_constant : std_logic_vector(7 downto 0);
    signal expr_228_wire_constant : std_logic_vector(7 downto 0);
    signal expr_235_wire_constant : std_logic_vector(7 downto 0);
    signal expr_242_wire_constant : std_logic_vector(7 downto 0);
    signal expr_249_wire_constant : std_logic_vector(7 downto 0);
    signal expr_256_wire_constant : std_logic_vector(7 downto 0);
    signal expr_263_wire_constant : std_logic_vector(7 downto 0);
    signal expr_270_wire_constant : std_logic_vector(7 downto 0);
    signal expr_277_wire_constant : std_logic_vector(7 downto 0);
    signal expr_284_wire_constant : std_logic_vector(7 downto 0);
    signal expr_291_wire_constant : std_logic_vector(7 downto 0);
    signal expr_298_wire_constant : std_logic_vector(7 downto 0);
    signal expr_305_wire_constant : std_logic_vector(7 downto 0);
    signal expr_312_wire_constant : std_logic_vector(7 downto 0);
    signal expr_319_wire_constant : std_logic_vector(7 downto 0);
    signal expr_326_wire_constant : std_logic_vector(7 downto 0);
    signal expr_333_wire_constant : std_logic_vector(7 downto 0);
    signal expr_340_wire_constant : std_logic_vector(7 downto 0);
    signal expr_347_wire_constant : std_logic_vector(7 downto 0);
    signal expr_354_wire_constant : std_logic_vector(7 downto 0);
    signal expr_361_wire_constant : std_logic_vector(7 downto 0);
    signal expr_368_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_176_word_address_0 <= "000000000";
    array_obj_ref_185_word_address_0 <= "000000001";
    array_obj_ref_192_word_address_0 <= "000000010";
    array_obj_ref_199_word_address_0 <= "000000011";
    array_obj_ref_206_word_address_0 <= "000000100";
    array_obj_ref_213_word_address_0 <= "000000101";
    array_obj_ref_220_word_address_0 <= "000000110";
    array_obj_ref_227_word_address_0 <= "001001000";
    array_obj_ref_234_word_address_0 <= "001001001";
    array_obj_ref_241_word_address_0 <= "001001010";
    array_obj_ref_248_word_address_0 <= "001001011";
    array_obj_ref_255_word_address_0 <= "001001100";
    array_obj_ref_262_word_address_0 <= "001001101";
    array_obj_ref_269_word_address_0 <= "001001110";
    array_obj_ref_276_word_address_0 <= "010010000";
    array_obj_ref_283_word_address_0 <= "010010001";
    array_obj_ref_290_word_address_0 <= "010010010";
    array_obj_ref_297_word_address_0 <= "010010011";
    array_obj_ref_304_word_address_0 <= "010010100";
    array_obj_ref_311_word_address_0 <= "010010101";
    array_obj_ref_318_word_address_0 <= "010010110";
    array_obj_ref_325_word_address_0 <= "011011000";
    array_obj_ref_332_word_address_0 <= "011011001";
    array_obj_ref_339_word_address_0 <= "011011010";
    array_obj_ref_346_word_address_0 <= "011011011";
    array_obj_ref_353_word_address_0 <= "011011100";
    array_obj_ref_360_word_address_0 <= "011011101";
    array_obj_ref_367_word_address_0 <= "011011110";
    expr_177_wire_constant <= "01110100";
    expr_186_wire_constant <= "01101111";
    expr_193_wire_constant <= "00110000";
    expr_200_wire_constant <= "01011111";
    expr_207_wire_constant <= "01101001";
    expr_214_wire_constant <= "01101110";
    expr_221_wire_constant <= "00110000";
    expr_228_wire_constant <= "01110100";
    expr_235_wire_constant <= "01101111";
    expr_242_wire_constant <= "00110001";
    expr_249_wire_constant <= "01011111";
    expr_256_wire_constant <= "01101001";
    expr_263_wire_constant <= "01101110";
    expr_270_wire_constant <= "00110000";
    expr_277_wire_constant <= "01110100";
    expr_284_wire_constant <= "01101111";
    expr_291_wire_constant <= "00110010";
    expr_298_wire_constant <= "01011111";
    expr_305_wire_constant <= "01101001";
    expr_312_wire_constant <= "01101110";
    expr_319_wire_constant <= "00110000";
    expr_326_wire_constant <= "01110100";
    expr_333_wire_constant <= "01101111";
    expr_340_wire_constant <= "00110011";
    expr_347_wire_constant <= "01011111";
    expr_354_wire_constant <= "01101001";
    expr_361_wire_constant <= "01101110";
    expr_368_wire_constant <= "00110000";
    array_obj_ref_176_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_176_gather_scatter_ack_0 <= array_obj_ref_176_gather_scatter_req_0;
      aggregated_sig <= expr_177_wire_constant;
      array_obj_ref_176_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_185_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_185_gather_scatter_ack_0 <= array_obj_ref_185_gather_scatter_req_0;
      aggregated_sig <= expr_186_wire_constant;
      array_obj_ref_185_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_192_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_192_gather_scatter_ack_0 <= array_obj_ref_192_gather_scatter_req_0;
      aggregated_sig <= expr_193_wire_constant;
      array_obj_ref_192_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_199_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_199_gather_scatter_ack_0 <= array_obj_ref_199_gather_scatter_req_0;
      aggregated_sig <= expr_200_wire_constant;
      array_obj_ref_199_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_206_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_206_gather_scatter_ack_0 <= array_obj_ref_206_gather_scatter_req_0;
      aggregated_sig <= expr_207_wire_constant;
      array_obj_ref_206_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_213_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_213_gather_scatter_ack_0 <= array_obj_ref_213_gather_scatter_req_0;
      aggregated_sig <= expr_214_wire_constant;
      array_obj_ref_213_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_220_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_220_gather_scatter_ack_0 <= array_obj_ref_220_gather_scatter_req_0;
      aggregated_sig <= expr_221_wire_constant;
      array_obj_ref_220_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_227_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_227_gather_scatter_ack_0 <= array_obj_ref_227_gather_scatter_req_0;
      aggregated_sig <= expr_228_wire_constant;
      array_obj_ref_227_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_234_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_234_gather_scatter_ack_0 <= array_obj_ref_234_gather_scatter_req_0;
      aggregated_sig <= expr_235_wire_constant;
      array_obj_ref_234_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_241_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_241_gather_scatter_ack_0 <= array_obj_ref_241_gather_scatter_req_0;
      aggregated_sig <= expr_242_wire_constant;
      array_obj_ref_241_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_248_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_248_gather_scatter_ack_0 <= array_obj_ref_248_gather_scatter_req_0;
      aggregated_sig <= expr_249_wire_constant;
      array_obj_ref_248_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_255_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_255_gather_scatter_ack_0 <= array_obj_ref_255_gather_scatter_req_0;
      aggregated_sig <= expr_256_wire_constant;
      array_obj_ref_255_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_262_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_262_gather_scatter_ack_0 <= array_obj_ref_262_gather_scatter_req_0;
      aggregated_sig <= expr_263_wire_constant;
      array_obj_ref_262_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_269_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_269_gather_scatter_ack_0 <= array_obj_ref_269_gather_scatter_req_0;
      aggregated_sig <= expr_270_wire_constant;
      array_obj_ref_269_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_276_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_276_gather_scatter_ack_0 <= array_obj_ref_276_gather_scatter_req_0;
      aggregated_sig <= expr_277_wire_constant;
      array_obj_ref_276_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_283_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_283_gather_scatter_ack_0 <= array_obj_ref_283_gather_scatter_req_0;
      aggregated_sig <= expr_284_wire_constant;
      array_obj_ref_283_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_290_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_290_gather_scatter_ack_0 <= array_obj_ref_290_gather_scatter_req_0;
      aggregated_sig <= expr_291_wire_constant;
      array_obj_ref_290_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_297_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_297_gather_scatter_ack_0 <= array_obj_ref_297_gather_scatter_req_0;
      aggregated_sig <= expr_298_wire_constant;
      array_obj_ref_297_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_304_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_304_gather_scatter_ack_0 <= array_obj_ref_304_gather_scatter_req_0;
      aggregated_sig <= expr_305_wire_constant;
      array_obj_ref_304_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_311_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_311_gather_scatter_ack_0 <= array_obj_ref_311_gather_scatter_req_0;
      aggregated_sig <= expr_312_wire_constant;
      array_obj_ref_311_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_318_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_318_gather_scatter_ack_0 <= array_obj_ref_318_gather_scatter_req_0;
      aggregated_sig <= expr_319_wire_constant;
      array_obj_ref_318_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_325_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_325_gather_scatter_ack_0 <= array_obj_ref_325_gather_scatter_req_0;
      aggregated_sig <= expr_326_wire_constant;
      array_obj_ref_325_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_332_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_332_gather_scatter_ack_0 <= array_obj_ref_332_gather_scatter_req_0;
      aggregated_sig <= expr_333_wire_constant;
      array_obj_ref_332_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_339_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_339_gather_scatter_ack_0 <= array_obj_ref_339_gather_scatter_req_0;
      aggregated_sig <= expr_340_wire_constant;
      array_obj_ref_339_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_346_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_346_gather_scatter_ack_0 <= array_obj_ref_346_gather_scatter_req_0;
      aggregated_sig <= expr_347_wire_constant;
      array_obj_ref_346_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_353_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_353_gather_scatter_ack_0 <= array_obj_ref_353_gather_scatter_req_0;
      aggregated_sig <= expr_354_wire_constant;
      array_obj_ref_353_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_360_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_360_gather_scatter_ack_0 <= array_obj_ref_360_gather_scatter_req_0;
      aggregated_sig <= expr_361_wire_constant;
      array_obj_ref_360_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_367_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_367_gather_scatter_ack_0 <= array_obj_ref_367_gather_scatter_req_0;
      aggregated_sig <= expr_368_wire_constant;
      array_obj_ref_367_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if array_obj_ref_176_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_176_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_176_word_address_0) &  " data array_obj_ref_176_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_176_data_0) severity note; --
        end if;
        if array_obj_ref_185_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_185_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_185_word_address_0) &  " data array_obj_ref_185_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_185_data_0) severity note; --
        end if;
        if array_obj_ref_192_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_192_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_192_word_address_0) &  " data array_obj_ref_192_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_192_data_0) severity note; --
        end if;
        if array_obj_ref_199_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_199_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_199_word_address_0) &  " data array_obj_ref_199_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_199_data_0) severity note; --
        end if;
        if array_obj_ref_206_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_206_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_206_word_address_0) &  " data array_obj_ref_206_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_206_data_0) severity note; --
        end if;
        if array_obj_ref_213_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_213_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_213_word_address_0) &  " data array_obj_ref_213_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_213_data_0) severity note; --
        end if;
        if array_obj_ref_220_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_220_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_220_word_address_0) &  " data array_obj_ref_220_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_220_data_0) severity note; --
        end if;
        if array_obj_ref_227_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_227_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_227_word_address_0) &  " data array_obj_ref_227_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_227_data_0) severity note; --
        end if;
        if array_obj_ref_234_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_234_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_234_word_address_0) &  " data array_obj_ref_234_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_234_data_0) severity note; --
        end if;
        if array_obj_ref_241_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_241_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_241_word_address_0) &  " data array_obj_ref_241_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_241_data_0) severity note; --
        end if;
        if array_obj_ref_248_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_248_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_248_word_address_0) &  " data array_obj_ref_248_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_248_data_0) severity note; --
        end if;
        if array_obj_ref_255_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_255_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_255_word_address_0) &  " data array_obj_ref_255_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_255_data_0) severity note; --
        end if;
        if array_obj_ref_262_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_262_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_262_word_address_0) &  " data array_obj_ref_262_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_262_data_0) severity note; --
        end if;
        if array_obj_ref_269_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_269_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_269_word_address_0) &  " data array_obj_ref_269_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_269_data_0) severity note; --
        end if;
        if array_obj_ref_276_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_276_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_276_word_address_0) &  " data array_obj_ref_276_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_276_data_0) severity note; --
        end if;
        if array_obj_ref_283_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_283_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_283_word_address_0) &  " data array_obj_ref_283_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_283_data_0) severity note; --
        end if;
        if array_obj_ref_290_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_290_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_290_word_address_0) &  " data array_obj_ref_290_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_290_data_0) severity note; --
        end if;
        if array_obj_ref_297_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_297_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_297_word_address_0) &  " data array_obj_ref_297_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_297_data_0) severity note; --
        end if;
        if array_obj_ref_304_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_304_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_304_word_address_0) &  " data array_obj_ref_304_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_304_data_0) severity note; --
        end if;
        if array_obj_ref_311_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_311_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_311_word_address_0) &  " data array_obj_ref_311_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_311_data_0) severity note; --
        end if;
        if array_obj_ref_318_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_318_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_318_word_address_0) &  " data array_obj_ref_318_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_318_data_0) severity note; --
        end if;
        if array_obj_ref_325_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_325_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_325_word_address_0) &  " data array_obj_ref_325_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_325_data_0) severity note; --
        end if;
        if array_obj_ref_332_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_332_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_332_word_address_0) &  " data array_obj_ref_332_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_332_data_0) severity note; --
        end if;
        if array_obj_ref_339_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_339_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_339_word_address_0) &  " data array_obj_ref_339_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_339_data_0) severity note; --
        end if;
        if array_obj_ref_346_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_346_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_346_word_address_0) &  " data array_obj_ref_346_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_346_data_0) severity note; --
        end if;
        if array_obj_ref_353_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_353_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_353_word_address_0) &  " data array_obj_ref_353_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_353_data_0) severity note; --
        end if;
        if array_obj_ref_360_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_360_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_360_word_address_0) &  " data array_obj_ref_360_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_360_data_0) severity note; --
        end if;
        if array_obj_ref_367_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_367_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_367_word_address_0) &  " data array_obj_ref_367_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_367_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : array_obj_ref_176_store_0 array_obj_ref_185_store_0 array_obj_ref_192_store_0 array_obj_ref_199_store_0 array_obj_ref_206_store_0 array_obj_ref_213_store_0 array_obj_ref_220_store_0 array_obj_ref_227_store_0 array_obj_ref_234_store_0 array_obj_ref_241_store_0 array_obj_ref_248_store_0 array_obj_ref_255_store_0 array_obj_ref_262_store_0 array_obj_ref_269_store_0 array_obj_ref_276_store_0 array_obj_ref_283_store_0 array_obj_ref_290_store_0 array_obj_ref_297_store_0 array_obj_ref_304_store_0 array_obj_ref_311_store_0 array_obj_ref_318_store_0 array_obj_ref_325_store_0 array_obj_ref_332_store_0 array_obj_ref_339_store_0 array_obj_ref_346_store_0 array_obj_ref_353_store_0 array_obj_ref_360_store_0 array_obj_ref_367_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(251 downto 0);
      signal data_in: std_logic_vector(223 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 27 downto 0);
      -- 
    begin -- 
      reqL(27) <= array_obj_ref_176_store_0_req_0;
      reqL(26) <= array_obj_ref_185_store_0_req_0;
      reqL(25) <= array_obj_ref_192_store_0_req_0;
      reqL(24) <= array_obj_ref_199_store_0_req_0;
      reqL(23) <= array_obj_ref_206_store_0_req_0;
      reqL(22) <= array_obj_ref_213_store_0_req_0;
      reqL(21) <= array_obj_ref_220_store_0_req_0;
      reqL(20) <= array_obj_ref_227_store_0_req_0;
      reqL(19) <= array_obj_ref_234_store_0_req_0;
      reqL(18) <= array_obj_ref_241_store_0_req_0;
      reqL(17) <= array_obj_ref_248_store_0_req_0;
      reqL(16) <= array_obj_ref_255_store_0_req_0;
      reqL(15) <= array_obj_ref_262_store_0_req_0;
      reqL(14) <= array_obj_ref_269_store_0_req_0;
      reqL(13) <= array_obj_ref_276_store_0_req_0;
      reqL(12) <= array_obj_ref_283_store_0_req_0;
      reqL(11) <= array_obj_ref_290_store_0_req_0;
      reqL(10) <= array_obj_ref_297_store_0_req_0;
      reqL(9) <= array_obj_ref_304_store_0_req_0;
      reqL(8) <= array_obj_ref_311_store_0_req_0;
      reqL(7) <= array_obj_ref_318_store_0_req_0;
      reqL(6) <= array_obj_ref_325_store_0_req_0;
      reqL(5) <= array_obj_ref_332_store_0_req_0;
      reqL(4) <= array_obj_ref_339_store_0_req_0;
      reqL(3) <= array_obj_ref_346_store_0_req_0;
      reqL(2) <= array_obj_ref_353_store_0_req_0;
      reqL(1) <= array_obj_ref_360_store_0_req_0;
      reqL(0) <= array_obj_ref_367_store_0_req_0;
      array_obj_ref_176_store_0_ack_0 <= ackL(27);
      array_obj_ref_185_store_0_ack_0 <= ackL(26);
      array_obj_ref_192_store_0_ack_0 <= ackL(25);
      array_obj_ref_199_store_0_ack_0 <= ackL(24);
      array_obj_ref_206_store_0_ack_0 <= ackL(23);
      array_obj_ref_213_store_0_ack_0 <= ackL(22);
      array_obj_ref_220_store_0_ack_0 <= ackL(21);
      array_obj_ref_227_store_0_ack_0 <= ackL(20);
      array_obj_ref_234_store_0_ack_0 <= ackL(19);
      array_obj_ref_241_store_0_ack_0 <= ackL(18);
      array_obj_ref_248_store_0_ack_0 <= ackL(17);
      array_obj_ref_255_store_0_ack_0 <= ackL(16);
      array_obj_ref_262_store_0_ack_0 <= ackL(15);
      array_obj_ref_269_store_0_ack_0 <= ackL(14);
      array_obj_ref_276_store_0_ack_0 <= ackL(13);
      array_obj_ref_283_store_0_ack_0 <= ackL(12);
      array_obj_ref_290_store_0_ack_0 <= ackL(11);
      array_obj_ref_297_store_0_ack_0 <= ackL(10);
      array_obj_ref_304_store_0_ack_0 <= ackL(9);
      array_obj_ref_311_store_0_ack_0 <= ackL(8);
      array_obj_ref_318_store_0_ack_0 <= ackL(7);
      array_obj_ref_325_store_0_ack_0 <= ackL(6);
      array_obj_ref_332_store_0_ack_0 <= ackL(5);
      array_obj_ref_339_store_0_ack_0 <= ackL(4);
      array_obj_ref_346_store_0_ack_0 <= ackL(3);
      array_obj_ref_353_store_0_ack_0 <= ackL(2);
      array_obj_ref_360_store_0_ack_0 <= ackL(1);
      array_obj_ref_367_store_0_ack_0 <= ackL(0);
      reqR(27) <= array_obj_ref_176_store_0_req_1;
      reqR(26) <= array_obj_ref_185_store_0_req_1;
      reqR(25) <= array_obj_ref_192_store_0_req_1;
      reqR(24) <= array_obj_ref_199_store_0_req_1;
      reqR(23) <= array_obj_ref_206_store_0_req_1;
      reqR(22) <= array_obj_ref_213_store_0_req_1;
      reqR(21) <= array_obj_ref_220_store_0_req_1;
      reqR(20) <= array_obj_ref_227_store_0_req_1;
      reqR(19) <= array_obj_ref_234_store_0_req_1;
      reqR(18) <= array_obj_ref_241_store_0_req_1;
      reqR(17) <= array_obj_ref_248_store_0_req_1;
      reqR(16) <= array_obj_ref_255_store_0_req_1;
      reqR(15) <= array_obj_ref_262_store_0_req_1;
      reqR(14) <= array_obj_ref_269_store_0_req_1;
      reqR(13) <= array_obj_ref_276_store_0_req_1;
      reqR(12) <= array_obj_ref_283_store_0_req_1;
      reqR(11) <= array_obj_ref_290_store_0_req_1;
      reqR(10) <= array_obj_ref_297_store_0_req_1;
      reqR(9) <= array_obj_ref_304_store_0_req_1;
      reqR(8) <= array_obj_ref_311_store_0_req_1;
      reqR(7) <= array_obj_ref_318_store_0_req_1;
      reqR(6) <= array_obj_ref_325_store_0_req_1;
      reqR(5) <= array_obj_ref_332_store_0_req_1;
      reqR(4) <= array_obj_ref_339_store_0_req_1;
      reqR(3) <= array_obj_ref_346_store_0_req_1;
      reqR(2) <= array_obj_ref_353_store_0_req_1;
      reqR(1) <= array_obj_ref_360_store_0_req_1;
      reqR(0) <= array_obj_ref_367_store_0_req_1;
      array_obj_ref_176_store_0_ack_1 <= ackR(27);
      array_obj_ref_185_store_0_ack_1 <= ackR(26);
      array_obj_ref_192_store_0_ack_1 <= ackR(25);
      array_obj_ref_199_store_0_ack_1 <= ackR(24);
      array_obj_ref_206_store_0_ack_1 <= ackR(23);
      array_obj_ref_213_store_0_ack_1 <= ackR(22);
      array_obj_ref_220_store_0_ack_1 <= ackR(21);
      array_obj_ref_227_store_0_ack_1 <= ackR(20);
      array_obj_ref_234_store_0_ack_1 <= ackR(19);
      array_obj_ref_241_store_0_ack_1 <= ackR(18);
      array_obj_ref_248_store_0_ack_1 <= ackR(17);
      array_obj_ref_255_store_0_ack_1 <= ackR(16);
      array_obj_ref_262_store_0_ack_1 <= ackR(15);
      array_obj_ref_269_store_0_ack_1 <= ackR(14);
      array_obj_ref_276_store_0_ack_1 <= ackR(13);
      array_obj_ref_283_store_0_ack_1 <= ackR(12);
      array_obj_ref_290_store_0_ack_1 <= ackR(11);
      array_obj_ref_297_store_0_ack_1 <= ackR(10);
      array_obj_ref_304_store_0_ack_1 <= ackR(9);
      array_obj_ref_311_store_0_ack_1 <= ackR(8);
      array_obj_ref_318_store_0_ack_1 <= ackR(7);
      array_obj_ref_325_store_0_ack_1 <= ackR(6);
      array_obj_ref_332_store_0_ack_1 <= ackR(5);
      array_obj_ref_339_store_0_ack_1 <= ackR(4);
      array_obj_ref_346_store_0_ack_1 <= ackR(3);
      array_obj_ref_353_store_0_ack_1 <= ackR(2);
      array_obj_ref_360_store_0_ack_1 <= ackR(1);
      array_obj_ref_367_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_176_word_address_0 & array_obj_ref_185_word_address_0 & array_obj_ref_192_word_address_0 & array_obj_ref_199_word_address_0 & array_obj_ref_206_word_address_0 & array_obj_ref_213_word_address_0 & array_obj_ref_220_word_address_0 & array_obj_ref_227_word_address_0 & array_obj_ref_234_word_address_0 & array_obj_ref_241_word_address_0 & array_obj_ref_248_word_address_0 & array_obj_ref_255_word_address_0 & array_obj_ref_262_word_address_0 & array_obj_ref_269_word_address_0 & array_obj_ref_276_word_address_0 & array_obj_ref_283_word_address_0 & array_obj_ref_290_word_address_0 & array_obj_ref_297_word_address_0 & array_obj_ref_304_word_address_0 & array_obj_ref_311_word_address_0 & array_obj_ref_318_word_address_0 & array_obj_ref_325_word_address_0 & array_obj_ref_332_word_address_0 & array_obj_ref_339_word_address_0 & array_obj_ref_346_word_address_0 & array_obj_ref_353_word_address_0 & array_obj_ref_360_word_address_0 & array_obj_ref_367_word_address_0;
      data_in <= array_obj_ref_176_data_0 & array_obj_ref_185_data_0 & array_obj_ref_192_data_0 & array_obj_ref_199_data_0 & array_obj_ref_206_data_0 & array_obj_ref_213_data_0 & array_obj_ref_220_data_0 & array_obj_ref_227_data_0 & array_obj_ref_234_data_0 & array_obj_ref_241_data_0 & array_obj_ref_248_data_0 & array_obj_ref_255_data_0 & array_obj_ref_262_data_0 & array_obj_ref_269_data_0 & array_obj_ref_276_data_0 & array_obj_ref_283_data_0 & array_obj_ref_290_data_0 & array_obj_ref_297_data_0 & array_obj_ref_304_data_0 & array_obj_ref_311_data_0 & array_obj_ref_318_data_0 & array_obj_ref_325_data_0 & array_obj_ref_332_data_0 & array_obj_ref_339_data_0 & array_obj_ref_346_data_0 & array_obj_ref_353_data_0 & array_obj_ref_360_data_0 & array_obj_ref_367_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 9,
        data_width => 8,
        num_reqs => 28,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(8 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 28,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity GV_16_initializer_in_click_bc is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity GV_16_initializer_in_click_bc;
architecture Default of GV_16_initializer_in_click_bc is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal GV_16_initializer_in_click_bc_CP_591_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_376_gather_scatter_req_0 : boolean;
  signal array_obj_ref_376_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_376_store_0_req_0 : boolean;
  signal array_obj_ref_376_store_0_ack_0 : boolean;
  signal array_obj_ref_376_store_0_req_1 : boolean;
  signal array_obj_ref_376_store_0_ack_1 : boolean;
  signal array_obj_ref_388_gather_scatter_req_0 : boolean;
  signal array_obj_ref_388_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_388_store_0_req_0 : boolean;
  signal array_obj_ref_388_store_0_ack_0 : boolean;
  signal array_obj_ref_388_store_0_req_1 : boolean;
  signal array_obj_ref_388_store_0_ack_1 : boolean;
  signal array_obj_ref_395_gather_scatter_req_0 : boolean;
  signal array_obj_ref_395_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_395_store_0_req_0 : boolean;
  signal array_obj_ref_395_store_0_ack_0 : boolean;
  signal array_obj_ref_395_store_0_req_1 : boolean;
  signal array_obj_ref_395_store_0_ack_1 : boolean;
  signal array_obj_ref_402_gather_scatter_req_0 : boolean;
  signal array_obj_ref_402_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_402_store_0_req_0 : boolean;
  signal array_obj_ref_402_store_0_ack_0 : boolean;
  signal array_obj_ref_402_store_0_req_1 : boolean;
  signal array_obj_ref_402_store_0_ack_1 : boolean;
  signal array_obj_ref_410_gather_scatter_req_0 : boolean;
  signal array_obj_ref_410_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_410_store_0_req_0 : boolean;
  signal array_obj_ref_410_store_0_ack_0 : boolean;
  signal array_obj_ref_410_store_0_req_1 : boolean;
  signal array_obj_ref_410_store_0_ack_1 : boolean;
  signal array_obj_ref_417_gather_scatter_req_0 : boolean;
  signal array_obj_ref_417_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_417_store_0_req_0 : boolean;
  signal array_obj_ref_417_store_0_ack_0 : boolean;
  signal array_obj_ref_417_store_0_req_1 : boolean;
  signal array_obj_ref_417_store_0_ack_1 : boolean;
  signal array_obj_ref_423_gather_scatter_req_0 : boolean;
  signal array_obj_ref_423_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_423_store_0_req_0 : boolean;
  signal array_obj_ref_423_store_0_ack_0 : boolean;
  signal array_obj_ref_423_store_0_req_1 : boolean;
  signal array_obj_ref_423_store_0_ack_1 : boolean;
  signal array_obj_ref_430_gather_scatter_req_0 : boolean;
  signal array_obj_ref_430_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_430_store_0_req_0 : boolean;
  signal array_obj_ref_430_store_0_ack_0 : boolean;
  signal array_obj_ref_430_store_0_req_1 : boolean;
  signal array_obj_ref_430_store_0_ack_1 : boolean;
  signal array_obj_ref_438_gather_scatter_req_0 : boolean;
  signal array_obj_ref_438_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_0 : boolean;
  signal array_obj_ref_438_store_0_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_1 : boolean;
  signal array_obj_ref_438_store_0_ack_1 : boolean;
  signal array_obj_ref_445_gather_scatter_req_0 : boolean;
  signal array_obj_ref_445_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_445_store_0_req_0 : boolean;
  signal array_obj_ref_445_store_0_ack_0 : boolean;
  signal array_obj_ref_445_store_0_req_1 : boolean;
  signal array_obj_ref_445_store_0_ack_1 : boolean;
  signal array_obj_ref_451_gather_scatter_req_0 : boolean;
  signal array_obj_ref_451_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_451_store_0_req_0 : boolean;
  signal array_obj_ref_451_store_0_ack_0 : boolean;
  signal array_obj_ref_451_store_0_req_1 : boolean;
  signal array_obj_ref_451_store_0_ack_1 : boolean;
  signal array_obj_ref_458_gather_scatter_req_0 : boolean;
  signal array_obj_ref_458_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_0 : boolean;
  signal array_obj_ref_458_store_0_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_1 : boolean;
  signal array_obj_ref_458_store_0_ack_1 : boolean;
  signal array_obj_ref_466_gather_scatter_req_0 : boolean;
  signal array_obj_ref_466_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_0 : boolean;
  signal array_obj_ref_466_store_0_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_1 : boolean;
  signal array_obj_ref_466_store_0_ack_1 : boolean;
  signal array_obj_ref_473_gather_scatter_req_0 : boolean;
  signal array_obj_ref_473_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_473_store_0_req_0 : boolean;
  signal array_obj_ref_473_store_0_ack_0 : boolean;
  signal array_obj_ref_473_store_0_req_1 : boolean;
  signal array_obj_ref_473_store_0_ack_1 : boolean;
  signal array_obj_ref_479_gather_scatter_req_0 : boolean;
  signal array_obj_ref_479_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_479_store_0_req_0 : boolean;
  signal array_obj_ref_479_store_0_ack_0 : boolean;
  signal array_obj_ref_479_store_0_req_1 : boolean;
  signal array_obj_ref_479_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  GV_16_initializer_in_click_bc_CP_591: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    split_req_603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => array_obj_ref_376_gather_scatter_req_0); -- 
    split_ack_604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_376_gather_scatter_ack_0, ack => cp_elements(1)); -- 
    rr_611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => array_obj_ref_376_store_0_req_0); -- 
    ra_612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_376_store_0_ack_0, ack => cp_elements(2)); -- 
    cr_613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => array_obj_ref_376_store_0_req_1); -- 
    ca_614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_376_store_0_ack_1, ack => cp_elements(3)); -- 
    split_req_624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => array_obj_ref_388_gather_scatter_req_0); -- 
    split_ack_625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_388_gather_scatter_ack_0, ack => cp_elements(4)); -- 
    rr_632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => array_obj_ref_388_store_0_req_0); -- 
    ra_633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_388_store_0_ack_0, ack => cp_elements(5)); -- 
    cr_634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => array_obj_ref_388_store_0_req_1); -- 
    ca_635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_388_store_0_ack_1, ack => cp_elements(6)); -- 
    split_req_645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => array_obj_ref_395_gather_scatter_req_0); -- 
    split_ack_646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_395_gather_scatter_ack_0, ack => cp_elements(7)); -- 
    rr_653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => array_obj_ref_395_store_0_req_0); -- 
    ra_654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_395_store_0_ack_0, ack => cp_elements(8)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => array_obj_ref_395_store_0_req_1); -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_395_store_0_ack_1, ack => cp_elements(9)); -- 
    split_req_666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => array_obj_ref_402_gather_scatter_req_0); -- 
    split_ack_667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_gather_scatter_ack_0, ack => cp_elements(10)); -- 
    rr_674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => array_obj_ref_402_store_0_req_0); -- 
    ra_675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_store_0_ack_0, ack => cp_elements(11)); -- 
    cr_676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => array_obj_ref_402_store_0_req_1); -- 
    ca_677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_store_0_ack_1, ack => cp_elements(12)); -- 
    split_req_687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => array_obj_ref_410_gather_scatter_req_0); -- 
    split_ack_688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_gather_scatter_ack_0, ack => cp_elements(13)); -- 
    rr_695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => array_obj_ref_410_store_0_req_0); -- 
    ra_696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_store_0_ack_0, ack => cp_elements(14)); -- 
    cr_697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => array_obj_ref_410_store_0_req_1); -- 
    ca_698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_store_0_ack_1, ack => cp_elements(15)); -- 
    split_req_708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => array_obj_ref_417_gather_scatter_req_0); -- 
    split_ack_709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_417_gather_scatter_ack_0, ack => cp_elements(16)); -- 
    rr_716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_417_store_0_req_0); -- 
    ra_717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_417_store_0_ack_0, ack => cp_elements(17)); -- 
    cr_718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => array_obj_ref_417_store_0_req_1); -- 
    ca_719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_417_store_0_ack_1, ack => cp_elements(18)); -- 
    split_req_729_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => array_obj_ref_423_gather_scatter_req_0); -- 
    split_ack_730_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_gather_scatter_ack_0, ack => cp_elements(19)); -- 
    rr_737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => array_obj_ref_423_store_0_req_0); -- 
    ra_738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_store_0_ack_0, ack => cp_elements(20)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => array_obj_ref_423_store_0_req_1); -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_store_0_ack_1, ack => cp_elements(21)); -- 
    split_req_750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_430_gather_scatter_req_0); -- 
    split_ack_751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_430_store_0_req_0); -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_store_0_ack_0, ack => cp_elements(23)); -- 
    cr_760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => array_obj_ref_430_store_0_req_1); -- 
    ca_761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_store_0_ack_1, ack => cp_elements(24)); -- 
    split_req_771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => array_obj_ref_438_gather_scatter_req_0); -- 
    split_ack_772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_gather_scatter_ack_0, ack => cp_elements(25)); -- 
    rr_779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => array_obj_ref_438_store_0_req_0); -- 
    ra_780_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_store_0_ack_0, ack => cp_elements(26)); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => array_obj_ref_438_store_0_req_1); -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_store_0_ack_1, ack => cp_elements(27)); -- 
    split_req_792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => array_obj_ref_445_gather_scatter_req_0); -- 
    split_ack_793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_445_gather_scatter_ack_0, ack => cp_elements(28)); -- 
    rr_800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => array_obj_ref_445_store_0_req_0); -- 
    ra_801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_445_store_0_ack_0, ack => cp_elements(29)); -- 
    cr_802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => array_obj_ref_445_store_0_req_1); -- 
    ca_803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_445_store_0_ack_1, ack => cp_elements(30)); -- 
    split_req_813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => array_obj_ref_451_gather_scatter_req_0); -- 
    split_ack_814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_gather_scatter_ack_0, ack => cp_elements(31)); -- 
    rr_821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_451_store_0_req_0); -- 
    ra_822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_store_0_ack_0, ack => cp_elements(32)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_451_store_0_req_1); -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_store_0_ack_1, ack => cp_elements(33)); -- 
    split_req_834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_458_gather_scatter_req_0); -- 
    split_ack_835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_gather_scatter_ack_0, ack => cp_elements(34)); -- 
    rr_842_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_458_store_0_req_0); -- 
    ra_843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_store_0_ack_0, ack => cp_elements(35)); -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => array_obj_ref_458_store_0_req_1); -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_store_0_ack_1, ack => cp_elements(36)); -- 
    split_req_855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_466_gather_scatter_req_0); -- 
    split_ack_856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_466_gather_scatter_ack_0, ack => cp_elements(37)); -- 
    rr_863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_466_store_0_req_0); -- 
    ra_864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_466_store_0_ack_0, ack => cp_elements(38)); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_466_store_0_req_1); -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_466_store_0_ack_1, ack => cp_elements(39)); -- 
    split_req_876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => array_obj_ref_473_gather_scatter_req_0); -- 
    split_ack_877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_gather_scatter_ack_0, ack => cp_elements(40)); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => array_obj_ref_473_store_0_req_0); -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_store_0_ack_0, ack => cp_elements(41)); -- 
    cr_886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => array_obj_ref_473_store_0_req_1); -- 
    ca_887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_store_0_ack_1, ack => cp_elements(42)); -- 
    split_req_897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => array_obj_ref_479_gather_scatter_req_0); -- 
    split_ack_898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_479_gather_scatter_ack_0, ack => cp_elements(43)); -- 
    rr_905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => array_obj_ref_479_store_0_req_0); -- 
    ra_906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_479_store_0_ack_0, ack => cp_elements(44)); -- 
    cr_907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => array_obj_ref_479_store_0_req_1); -- 
    ca_908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_479_store_0_ack_1, ack => cp_elements(45)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_376_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_376_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_388_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_388_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_395_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_395_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_402_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_402_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_410_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_410_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_417_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_417_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_423_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_423_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_430_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_430_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_438_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_438_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_445_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_445_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_451_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_451_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_458_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_458_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_466_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_466_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_473_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_473_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_479_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_479_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_377_wire_constant : std_logic_vector(31 downto 0);
    signal expr_389_wire_constant : std_logic_vector(31 downto 0);
    signal expr_396_wire_constant : std_logic_vector(31 downto 0);
    signal expr_403_wire_constant : std_logic_vector(31 downto 0);
    signal expr_411_wire_constant : std_logic_vector(31 downto 0);
    signal expr_418_wire_constant : std_logic_vector(31 downto 0);
    signal expr_424_wire_constant : std_logic_vector(31 downto 0);
    signal expr_431_wire_constant : std_logic_vector(31 downto 0);
    signal expr_439_wire_constant : std_logic_vector(31 downto 0);
    signal expr_446_wire_constant : std_logic_vector(31 downto 0);
    signal expr_452_wire_constant : std_logic_vector(31 downto 0);
    signal expr_459_wire_constant : std_logic_vector(31 downto 0);
    signal expr_467_wire_constant : std_logic_vector(31 downto 0);
    signal expr_474_wire_constant : std_logic_vector(31 downto 0);
    signal expr_480_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_376_word_address_0 <= "00000";
    array_obj_ref_388_word_address_0 <= "00001";
    array_obj_ref_395_word_address_0 <= "00100";
    array_obj_ref_402_word_address_0 <= "00101";
    array_obj_ref_410_word_address_0 <= "00110";
    array_obj_ref_417_word_address_0 <= "01000";
    array_obj_ref_423_word_address_0 <= "01001";
    array_obj_ref_430_word_address_0 <= "01010";
    array_obj_ref_438_word_address_0 <= "01011";
    array_obj_ref_445_word_address_0 <= "01101";
    array_obj_ref_451_word_address_0 <= "01110";
    array_obj_ref_458_word_address_0 <= "01111";
    array_obj_ref_466_word_address_0 <= "10000";
    array_obj_ref_473_word_address_0 <= "10010";
    array_obj_ref_479_word_address_0 <= "10011";
    expr_377_wire_constant <= "00000000000000000001000010101100";
    expr_389_wire_constant <= "00000000111111111111111111111111";
    expr_396_wire_constant <= "01111111111111111111111111111111";
    expr_403_wire_constant <= "00000000000000010001000010101100";
    expr_411_wire_constant <= "00000000111111111111111111111111";
    expr_418_wire_constant <= "00000000000000000000000000000001";
    expr_424_wire_constant <= "01111111111111111111111111111111";
    expr_431_wire_constant <= "00000000000000100001000010101100";
    expr_439_wire_constant <= "00000000111111111111111111111111";
    expr_446_wire_constant <= "00000000000000000000000000000010";
    expr_452_wire_constant <= "01111111111111111111111111111111";
    expr_459_wire_constant <= "00000000000000110001000010101100";
    expr_467_wire_constant <= "00000000111111111111111111111111";
    expr_474_wire_constant <= "00000000000000000000000000000011";
    expr_480_wire_constant <= "01111111111111111111111111111111";
    array_obj_ref_376_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_376_gather_scatter_ack_0 <= array_obj_ref_376_gather_scatter_req_0;
      aggregated_sig <= expr_377_wire_constant;
      array_obj_ref_376_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_388_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_388_gather_scatter_ack_0 <= array_obj_ref_388_gather_scatter_req_0;
      aggregated_sig <= expr_389_wire_constant;
      array_obj_ref_388_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_395_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_395_gather_scatter_ack_0 <= array_obj_ref_395_gather_scatter_req_0;
      aggregated_sig <= expr_396_wire_constant;
      array_obj_ref_395_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_402_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_402_gather_scatter_ack_0 <= array_obj_ref_402_gather_scatter_req_0;
      aggregated_sig <= expr_403_wire_constant;
      array_obj_ref_402_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_410_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_410_gather_scatter_ack_0 <= array_obj_ref_410_gather_scatter_req_0;
      aggregated_sig <= expr_411_wire_constant;
      array_obj_ref_410_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_417_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_417_gather_scatter_ack_0 <= array_obj_ref_417_gather_scatter_req_0;
      aggregated_sig <= expr_418_wire_constant;
      array_obj_ref_417_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_423_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_423_gather_scatter_ack_0 <= array_obj_ref_423_gather_scatter_req_0;
      aggregated_sig <= expr_424_wire_constant;
      array_obj_ref_423_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_430_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_430_gather_scatter_ack_0 <= array_obj_ref_430_gather_scatter_req_0;
      aggregated_sig <= expr_431_wire_constant;
      array_obj_ref_430_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_438_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_438_gather_scatter_ack_0 <= array_obj_ref_438_gather_scatter_req_0;
      aggregated_sig <= expr_439_wire_constant;
      array_obj_ref_438_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_445_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_445_gather_scatter_ack_0 <= array_obj_ref_445_gather_scatter_req_0;
      aggregated_sig <= expr_446_wire_constant;
      array_obj_ref_445_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_451_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_451_gather_scatter_ack_0 <= array_obj_ref_451_gather_scatter_req_0;
      aggregated_sig <= expr_452_wire_constant;
      array_obj_ref_451_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_458_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_458_gather_scatter_ack_0 <= array_obj_ref_458_gather_scatter_req_0;
      aggregated_sig <= expr_459_wire_constant;
      array_obj_ref_458_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_466_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_466_gather_scatter_ack_0 <= array_obj_ref_466_gather_scatter_req_0;
      aggregated_sig <= expr_467_wire_constant;
      array_obj_ref_466_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_473_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_473_gather_scatter_ack_0 <= array_obj_ref_473_gather_scatter_req_0;
      aggregated_sig <= expr_474_wire_constant;
      array_obj_ref_473_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_479_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_479_gather_scatter_ack_0 <= array_obj_ref_479_gather_scatter_req_0;
      aggregated_sig <= expr_480_wire_constant;
      array_obj_ref_479_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if array_obj_ref_417_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_417_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_417_word_address_0) &  " data array_obj_ref_417_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_417_data_0) severity note; --
        end if;
        if array_obj_ref_466_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_466_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_466_word_address_0) &  " data array_obj_ref_466_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_466_data_0) severity note; --
        end if;
        if array_obj_ref_410_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_410_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_410_word_address_0) &  " data array_obj_ref_410_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_410_data_0) severity note; --
        end if;
        if array_obj_ref_458_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_458_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_458_word_address_0) &  " data array_obj_ref_458_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_458_data_0) severity note; --
        end if;
        if array_obj_ref_402_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_402_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_402_word_address_0) &  " data array_obj_ref_402_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_402_data_0) severity note; --
        end if;
        if array_obj_ref_451_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_451_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_451_word_address_0) &  " data array_obj_ref_451_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_451_data_0) severity note; --
        end if;
        if array_obj_ref_445_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_445_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_445_word_address_0) &  " data array_obj_ref_445_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_445_data_0) severity note; --
        end if;
        if array_obj_ref_395_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_395_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_395_word_address_0) &  " data array_obj_ref_395_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_395_data_0) severity note; --
        end if;
        if array_obj_ref_479_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_479_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_479_word_address_0) &  " data array_obj_ref_479_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_479_data_0) severity note; --
        end if;
        if array_obj_ref_438_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_438_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_438_word_address_0) &  " data array_obj_ref_438_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_438_data_0) severity note; --
        end if;
        if array_obj_ref_388_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_388_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_388_word_address_0) &  " data array_obj_ref_388_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_388_data_0) severity note; --
        end if;
        if array_obj_ref_430_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_430_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_430_word_address_0) &  " data array_obj_ref_430_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_430_data_0) severity note; --
        end if;
        if array_obj_ref_376_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_376_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_376_word_address_0) &  " data array_obj_ref_376_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_376_data_0) severity note; --
        end if;
        if array_obj_ref_423_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_423_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_423_word_address_0) &  " data array_obj_ref_423_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_423_data_0) severity note; --
        end if;
        if array_obj_ref_473_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_473_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_473_word_address_0) &  " data array_obj_ref_473_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_473_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : array_obj_ref_417_store_0 array_obj_ref_466_store_0 array_obj_ref_410_store_0 array_obj_ref_458_store_0 array_obj_ref_402_store_0 array_obj_ref_451_store_0 array_obj_ref_445_store_0 array_obj_ref_395_store_0 array_obj_ref_479_store_0 array_obj_ref_438_store_0 array_obj_ref_388_store_0 array_obj_ref_430_store_0 array_obj_ref_376_store_0 array_obj_ref_423_store_0 array_obj_ref_473_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(74 downto 0);
      signal data_in: std_logic_vector(479 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_417_store_0_req_0;
      reqL(13) <= array_obj_ref_466_store_0_req_0;
      reqL(12) <= array_obj_ref_410_store_0_req_0;
      reqL(11) <= array_obj_ref_458_store_0_req_0;
      reqL(10) <= array_obj_ref_402_store_0_req_0;
      reqL(9) <= array_obj_ref_451_store_0_req_0;
      reqL(8) <= array_obj_ref_445_store_0_req_0;
      reqL(7) <= array_obj_ref_395_store_0_req_0;
      reqL(6) <= array_obj_ref_479_store_0_req_0;
      reqL(5) <= array_obj_ref_438_store_0_req_0;
      reqL(4) <= array_obj_ref_388_store_0_req_0;
      reqL(3) <= array_obj_ref_430_store_0_req_0;
      reqL(2) <= array_obj_ref_376_store_0_req_0;
      reqL(1) <= array_obj_ref_423_store_0_req_0;
      reqL(0) <= array_obj_ref_473_store_0_req_0;
      array_obj_ref_417_store_0_ack_0 <= ackL(14);
      array_obj_ref_466_store_0_ack_0 <= ackL(13);
      array_obj_ref_410_store_0_ack_0 <= ackL(12);
      array_obj_ref_458_store_0_ack_0 <= ackL(11);
      array_obj_ref_402_store_0_ack_0 <= ackL(10);
      array_obj_ref_451_store_0_ack_0 <= ackL(9);
      array_obj_ref_445_store_0_ack_0 <= ackL(8);
      array_obj_ref_395_store_0_ack_0 <= ackL(7);
      array_obj_ref_479_store_0_ack_0 <= ackL(6);
      array_obj_ref_438_store_0_ack_0 <= ackL(5);
      array_obj_ref_388_store_0_ack_0 <= ackL(4);
      array_obj_ref_430_store_0_ack_0 <= ackL(3);
      array_obj_ref_376_store_0_ack_0 <= ackL(2);
      array_obj_ref_423_store_0_ack_0 <= ackL(1);
      array_obj_ref_473_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_417_store_0_req_1;
      reqR(13) <= array_obj_ref_466_store_0_req_1;
      reqR(12) <= array_obj_ref_410_store_0_req_1;
      reqR(11) <= array_obj_ref_458_store_0_req_1;
      reqR(10) <= array_obj_ref_402_store_0_req_1;
      reqR(9) <= array_obj_ref_451_store_0_req_1;
      reqR(8) <= array_obj_ref_445_store_0_req_1;
      reqR(7) <= array_obj_ref_395_store_0_req_1;
      reqR(6) <= array_obj_ref_479_store_0_req_1;
      reqR(5) <= array_obj_ref_438_store_0_req_1;
      reqR(4) <= array_obj_ref_388_store_0_req_1;
      reqR(3) <= array_obj_ref_430_store_0_req_1;
      reqR(2) <= array_obj_ref_376_store_0_req_1;
      reqR(1) <= array_obj_ref_423_store_0_req_1;
      reqR(0) <= array_obj_ref_473_store_0_req_1;
      array_obj_ref_417_store_0_ack_1 <= ackR(14);
      array_obj_ref_466_store_0_ack_1 <= ackR(13);
      array_obj_ref_410_store_0_ack_1 <= ackR(12);
      array_obj_ref_458_store_0_ack_1 <= ackR(11);
      array_obj_ref_402_store_0_ack_1 <= ackR(10);
      array_obj_ref_451_store_0_ack_1 <= ackR(9);
      array_obj_ref_445_store_0_ack_1 <= ackR(8);
      array_obj_ref_395_store_0_ack_1 <= ackR(7);
      array_obj_ref_479_store_0_ack_1 <= ackR(6);
      array_obj_ref_438_store_0_ack_1 <= ackR(5);
      array_obj_ref_388_store_0_ack_1 <= ackR(4);
      array_obj_ref_430_store_0_ack_1 <= ackR(3);
      array_obj_ref_376_store_0_ack_1 <= ackR(2);
      array_obj_ref_423_store_0_ack_1 <= ackR(1);
      array_obj_ref_473_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_417_word_address_0 & array_obj_ref_466_word_address_0 & array_obj_ref_410_word_address_0 & array_obj_ref_458_word_address_0 & array_obj_ref_402_word_address_0 & array_obj_ref_451_word_address_0 & array_obj_ref_445_word_address_0 & array_obj_ref_395_word_address_0 & array_obj_ref_479_word_address_0 & array_obj_ref_438_word_address_0 & array_obj_ref_388_word_address_0 & array_obj_ref_430_word_address_0 & array_obj_ref_376_word_address_0 & array_obj_ref_423_word_address_0 & array_obj_ref_473_word_address_0;
      data_in <= array_obj_ref_417_data_0 & array_obj_ref_466_data_0 & array_obj_ref_410_data_0 & array_obj_ref_458_data_0 & array_obj_ref_402_data_0 & array_obj_ref_451_data_0 & array_obj_ref_445_data_0 & array_obj_ref_395_data_0 & array_obj_ref_479_data_0 & array_obj_ref_438_data_0 & array_obj_ref_388_data_0 & array_obj_ref_430_data_0 & array_obj_ref_376_data_0 & array_obj_ref_423_data_0 & array_obj_ref_473_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 32,
        num_reqs => 15,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(4 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_bswap_i16 is -- 
  generic (tag_length : integer); 
  port ( -- 
    i : in  std_logic_vector(15 downto 0);
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_bswap_i16;
architecture Default of ahir_glue_bswap_i16 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_CP_969_start: Boolean;
  -- links between control-path and data-path
  signal binary_523_inst_ack_1 : boolean;
  signal binary_523_inst_ack_0 : boolean;
  signal binary_523_inst_req_1 : boolean;
  signal binary_528_inst_ack_1 : boolean;
  signal binary_528_inst_req_0 : boolean;
  signal binary_528_inst_ack_0 : boolean;
  signal binary_528_inst_req_1 : boolean;
  signal binary_523_inst_req_0 : boolean;
  signal binary_517_inst_req_1 : boolean;
  signal binary_517_inst_ack_1 : boolean;
  signal binary_517_inst_ack_0 : boolean;
  signal binary_517_inst_req_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  ret_val_x_x <= ret_val_x_x_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 3, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_bswap_i16_CP_969: Block -- control-path 
    signal cp_elements: BooleanArray(15 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(15);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(15), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    cpelement_group_2 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(4));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => binary_517_inst_req_0); -- 
    cp_elements(3) <= cp_elements(1);
    cp_elements(4) <= cp_elements(1);
    ra_993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_517_inst_ack_0, ack => cp_elements(5)); -- 
    cr_994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => binary_517_inst_req_1); -- 
    ca_995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_517_inst_ack_1, ack => cp_elements(6)); -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(8) & cp_elements(9));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => binary_523_inst_req_0); -- 
    cp_elements(8) <= cp_elements(1);
    cp_elements(9) <= cp_elements(1);
    ra_1005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_523_inst_ack_0, ack => cp_elements(10)); -- 
    cr_1006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => binary_523_inst_req_1); -- 
    ca_1007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_523_inst_ack_1, ack => cp_elements(11)); -- 
    cpelement_group_12 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(13) & cp_elements(6));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(12),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => binary_528_inst_req_0); -- 
    cp_elements(13) <= cp_elements(1);
    ra_1018_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_528_inst_ack_0, ack => cp_elements(14)); -- 
    cr_1019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => binary_528_inst_req_1); -- 
    ca_1020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_528_inst_ack_1, ack => cp_elements(15)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal tmp1_524 : std_logic_vector(15 downto 0);
    signal tmp_518 : std_logic_vector(15 downto 0);
    signal type_cast_516_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_522_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    type_cast_516_wire_constant <= "0000000000001000";
    type_cast_522_wire_constant <= "0000000000001000";
    -- shared split operator group (0) : binary_517_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i;
      tmp_518 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_517_inst_req_0,
          ackL => binary_517_inst_ack_0,
          reqR => binary_517_inst_req_1,
          ackR => binary_517_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_523_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i;
      tmp1_524 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_523_inst_req_0,
          ackL => binary_523_inst_ack_0,
          reqR => binary_523_inst_req_1,
          ackR => binary_523_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_528_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_524 & tmp_518;
      ret_val_x_x_buffer <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_528_inst_req_0,
          ackL => binary_528_inst_ack_0,
          reqR => binary_528_inst_req_1,
          ackR => binary_528_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_chk is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    chk_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    chk_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    chk_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    rtt_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    rtt_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    rtt_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    ahir_packet_free_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_free_call_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_free_call_data : out  std_logic_vector(31 downto 0);
    ahir_packet_free_call_tag  :  out  std_logic_vector(2 downto 0);
    ahir_packet_free_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_free_return_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_free_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_chk;
architecture Default of ahir_glue_chk is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_chk_CP_1053_start: Boolean;
  -- links between control-path and data-path
  signal binary_588_inst_ack_0 : boolean;
  signal binary_597_inst_req_1 : boolean;
  signal binary_588_inst_req_1 : boolean;
  signal ptr_deref_1060_addr_1_req_0 : boolean;
  signal binary_588_inst_ack_1 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal ptr_deref_616_addr_2_ack_0 : boolean;
  signal ptr_deref_616_load_3_req_1 : boolean;
  signal ptr_deref_616_load_1_req_1 : boolean;
  signal ptr_deref_960_addr_2_ack_1 : boolean;
  signal ptr_deref_616_load_2_ack_1 : boolean;
  signal if_stmt_968_branch_req_0 : boolean;
  signal ptr_deref_960_addr_1_ack_1 : boolean;
  signal ptr_deref_960_store_1_req_0 : boolean;
  signal ptr_deref_960_store_1_ack_0 : boolean;
  signal ptr_deref_960_addr_3_req_0 : boolean;
  signal ptr_deref_1060_addr_3_req_0 : boolean;
  signal binary_983_inst_ack_1 : boolean;
  signal ptr_deref_616_load_1_req_0 : boolean;
  signal ptr_deref_616_load_2_req_1 : boolean;
  signal binary_597_inst_ack_0 : boolean;
  signal ptr_deref_1060_addr_0_ack_1 : boolean;
  signal ptr_deref_616_load_1_ack_1 : boolean;
  signal ptr_deref_960_store_0_req_0 : boolean;
  signal ptr_deref_960_store_0_ack_0 : boolean;
  signal if_stmt_968_branch_ack_1 : boolean;
  signal ptr_deref_569_load_0_req_0 : boolean;
  signal ptr_deref_1060_addr_1_ack_0 : boolean;
  signal ptr_deref_569_load_0_ack_0 : boolean;
  signal ptr_deref_616_root_address_inst_req_0 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal ptr_deref_569_load_2_req_0 : boolean;
  signal ptr_deref_616_root_address_inst_ack_0 : boolean;
  signal call_stmt_607_call_req_0 : boolean;
  signal binary_1067_inst_ack_0 : boolean;
  signal ptr_deref_569_load_3_req_0 : boolean;
  signal type_cast_845_inst_req_0 : boolean;
  signal type_cast_612_inst_req_0 : boolean;
  signal ptr_deref_569_load_3_ack_0 : boolean;
  signal type_cast_612_inst_ack_0 : boolean;
  signal binary_1067_inst_req_1 : boolean;
  signal ptr_deref_569_load_1_req_0 : boolean;
  signal ptr_deref_616_load_2_ack_0 : boolean;
  signal ptr_deref_616_addr_3_ack_1 : boolean;
  signal phi_stmt_840_ack_0 : boolean;
  signal binary_1067_inst_ack_1 : boolean;
  signal binary_966_inst_ack_1 : boolean;
  signal call_stmt_607_call_ack_0 : boolean;
  signal ptr_deref_569_load_1_ack_0 : boolean;
  signal call_stmt_648_call_req_0 : boolean;
  signal call_stmt_648_call_ack_0 : boolean;
  signal ptr_deref_616_addr_0_req_0 : boolean;
  signal ptr_deref_1060_addr_2_req_1 : boolean;
  signal if_stmt_599_branch_ack_0 : boolean;
  signal ptr_deref_616_addr_0_ack_0 : boolean;
  signal ptr_deref_1060_store_3_req_1 : boolean;
  signal ptr_deref_616_addr_2_req_1 : boolean;
  signal ptr_deref_1060_addr_2_ack_0 : boolean;
  signal ptr_deref_616_addr_0_req_1 : boolean;
  signal call_stmt_648_call_req_1 : boolean;
  signal ptr_deref_616_addr_0_ack_1 : boolean;
  signal if_stmt_640_branch_req_0 : boolean;
  signal call_stmt_648_call_ack_1 : boolean;
  signal ptr_deref_569_load_0_req_1 : boolean;
  signal ptr_deref_569_load_0_ack_1 : boolean;
  signal ptr_deref_616_addr_1_req_0 : boolean;
  signal ptr_deref_616_addr_1_ack_0 : boolean;
  signal ptr_deref_1060_addr_0_req_0 : boolean;
  signal ptr_deref_1060_addr_1_req_1 : boolean;
  signal if_stmt_1069_branch_req_0 : boolean;
  signal if_stmt_640_branch_ack_1 : boolean;
  signal ptr_deref_616_addr_1_req_1 : boolean;
  signal ptr_deref_1060_addr_2_ack_1 : boolean;
  signal ptr_deref_569_load_1_req_1 : boolean;
  signal ptr_deref_616_addr_2_ack_1 : boolean;
  signal ptr_deref_616_load_0_ack_0 : boolean;
  signal type_cast_845_inst_ack_0 : boolean;
  signal ptr_deref_569_load_2_ack_1 : boolean;
  signal binary_655_inst_req_0 : boolean;
  signal ptr_deref_616_gather_scatter_ack_0 : boolean;
  signal ptr_deref_569_load_3_req_1 : boolean;
  signal binary_634_inst_req_0 : boolean;
  signal binary_634_inst_req_1 : boolean;
  signal binary_667_inst_ack_0 : boolean;
  signal ptr_deref_616_addr_2_req_0 : boolean;
  signal ptr_deref_616_load_0_req_1 : boolean;
  signal ptr_deref_616_load_0_ack_1 : boolean;
  signal binary_667_inst_ack_1 : boolean;
  signal type_cast_573_inst_req_0 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal binary_966_inst_req_0 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal call_stmt_677_call_req_0 : boolean;
  signal type_cast_573_inst_ack_0 : boolean;
  signal binary_966_inst_req_1 : boolean;
  signal ptr_deref_616_load_3_req_0 : boolean;
  signal if_stmt_669_branch_ack_0 : boolean;
  signal ptr_deref_960_addr_1_req_1 : boolean;
  signal type_cast_740_inst_ack_0 : boolean;
  signal phi_stmt_840_req_1 : boolean;
  signal binary_661_inst_req_1 : boolean;
  signal ptr_deref_1060_addr_1_ack_1 : boolean;
  signal binary_597_inst_req_0 : boolean;
  signal ptr_deref_569_load_2_ack_0 : boolean;
  signal binary_628_inst_req_0 : boolean;
  signal ptr_deref_616_load_3_ack_0 : boolean;
  signal ptr_deref_616_load_2_req_0 : boolean;
  signal if_stmt_1069_branch_ack_1 : boolean;
  signal ptr_deref_1060_addr_2_req_0 : boolean;
  signal binary_588_inst_req_0 : boolean;
  signal ptr_deref_960_addr_2_req_1 : boolean;
  signal binary_628_inst_ack_0 : boolean;
  signal ptr_deref_1060_addr_0_ack_0 : boolean;
  signal ptr_deref_616_addr_3_req_1 : boolean;
  signal ptr_deref_960_gather_scatter_ack_0 : boolean;
  signal ptr_deref_616_load_1_ack_0 : boolean;
  signal binary_628_inst_req_1 : boolean;
  signal ptr_deref_960_addr_2_ack_0 : boolean;
  signal ptr_deref_616_addr_3_ack_0 : boolean;
  signal phi_stmt_834_ack_0 : boolean;
  signal ptr_deref_1060_addr_0_req_1 : boolean;
  signal binary_628_inst_ack_1 : boolean;
  signal binary_1067_inst_req_0 : boolean;
  signal if_stmt_669_branch_ack_1 : boolean;
  signal binary_661_inst_ack_1 : boolean;
  signal ptr_deref_569_load_1_ack_1 : boolean;
  signal ptr_deref_1060_addr_3_ack_0 : boolean;
  signal binary_622_inst_req_0 : boolean;
  signal phi_stmt_734_req_1 : boolean;
  signal if_stmt_669_branch_req_0 : boolean;
  signal ptr_deref_616_base_resize_req_0 : boolean;
  signal binary_622_inst_ack_0 : boolean;
  signal binary_634_inst_ack_0 : boolean;
  signal binary_582_inst_ack_0 : boolean;
  signal ptr_deref_616_addr_1_ack_1 : boolean;
  signal call_stmt_677_call_ack_1 : boolean;
  signal if_stmt_1069_branch_ack_0 : boolean;
  signal binary_667_inst_req_0 : boolean;
  signal binary_597_inst_ack_1 : boolean;
  signal ptr_deref_616_load_3_ack_1 : boolean;
  signal binary_582_inst_req_0 : boolean;
  signal call_stmt_677_call_ack_0 : boolean;
  signal if_stmt_640_branch_ack_0 : boolean;
  signal call_stmt_682_call_req_1 : boolean;
  signal call_stmt_682_call_ack_1 : boolean;
  signal call_stmt_682_call_ack_0 : boolean;
  signal ptr_deref_1060_addr_3_req_1 : boolean;
  signal if_stmt_599_branch_req_0 : boolean;
  signal binary_966_inst_ack_0 : boolean;
  signal binary_622_inst_req_1 : boolean;
  signal binary_655_inst_req_1 : boolean;
  signal binary_582_inst_req_1 : boolean;
  signal ptr_deref_960_addr_1_ack_0 : boolean;
  signal ptr_deref_616_gather_scatter_req_0 : boolean;
  signal type_cast_740_inst_req_0 : boolean;
  signal type_cast_638_inst_req_0 : boolean;
  signal binary_582_inst_ack_1 : boolean;
  signal ptr_deref_616_load_0_req_0 : boolean;
  signal binary_622_inst_ack_1 : boolean;
  signal binary_661_inst_ack_0 : boolean;
  signal binary_655_inst_ack_1 : boolean;
  signal ptr_deref_616_base_resize_ack_0 : boolean;
  signal type_cast_638_inst_ack_0 : boolean;
  signal ptr_deref_569_load_2_req_1 : boolean;
  signal binary_661_inst_req_0 : boolean;
  signal ptr_deref_616_addr_3_req_0 : boolean;
  signal ptr_deref_1060_addr_3_ack_1 : boolean;
  signal call_stmt_607_call_req_1 : boolean;
  signal ptr_deref_569_load_3_ack_1 : boolean;
  signal ptr_deref_569_gather_scatter_req_0 : boolean;
  signal binary_634_inst_ack_1 : boolean;
  signal ptr_deref_569_gather_scatter_ack_0 : boolean;
  signal if_stmt_599_branch_ack_1 : boolean;
  signal call_stmt_682_call_req_0 : boolean;
  signal binary_655_inst_ack_0 : boolean;
  signal call_stmt_607_call_ack_1 : boolean;
  signal binary_690_inst_req_1 : boolean;
  signal binary_690_inst_ack_1 : boolean;
  signal binary_690_inst_req_0 : boolean;
  signal binary_690_inst_ack_0 : boolean;
  signal type_cast_685_inst_req_0 : boolean;
  signal type_cast_843_inst_ack_0 : boolean;
  signal binary_667_inst_req_1 : boolean;
  signal type_cast_685_inst_ack_0 : boolean;
  signal type_cast_843_inst_req_0 : boolean;
  signal ptr_deref_1060_gather_scatter_req_0 : boolean;
  signal call_stmt_677_call_req_1 : boolean;
  signal type_cast_747_inst_req_0 : boolean;
  signal type_cast_747_inst_ack_0 : boolean;
  signal ternary_989_inst_ack_0 : boolean;
  signal if_stmt_968_branch_ack_0 : boolean;
  signal ptr_deref_960_addr_3_ack_0 : boolean;
  signal ptr_deref_960_store_2_req_0 : boolean;
  signal ptr_deref_960_store_2_ack_0 : boolean;
  signal ptr_deref_960_store_3_req_0 : boolean;
  signal binary_995_inst_req_1 : boolean;
  signal ptr_deref_960_store_3_ack_0 : boolean;
  signal ptr_deref_960_addr_3_req_1 : boolean;
  signal ptr_deref_960_base_resize_req_0 : boolean;
  signal binary_983_inst_req_0 : boolean;
  signal ptr_deref_960_addr_3_ack_1 : boolean;
  signal binary_995_inst_ack_1 : boolean;
  signal ptr_deref_960_base_resize_ack_0 : boolean;
  signal ternary_989_inst_req_0 : boolean;
  signal binary_995_inst_ack_0 : boolean;
  signal ptr_deref_960_root_address_inst_req_0 : boolean;
  signal ptr_deref_960_root_address_inst_ack_0 : boolean;
  signal ptr_deref_960_store_0_req_1 : boolean;
  signal ptr_deref_960_store_0_ack_1 : boolean;
  signal ptr_deref_960_store_1_req_1 : boolean;
  signal ptr_deref_960_store_1_ack_1 : boolean;
  signal ptr_deref_960_store_2_req_1 : boolean;
  signal ptr_deref_960_store_2_ack_1 : boolean;
  signal ptr_deref_960_store_3_req_1 : boolean;
  signal ptr_deref_960_store_3_ack_1 : boolean;
  signal ptr_deref_960_addr_0_req_0 : boolean;
  signal binary_978_inst_req_0 : boolean;
  signal ptr_deref_960_addr_0_ack_0 : boolean;
  signal binary_995_inst_req_0 : boolean;
  signal binary_978_inst_ack_0 : boolean;
  signal binary_978_inst_req_1 : boolean;
  signal ptr_deref_960_addr_0_req_1 : boolean;
  signal simple_obj_ref_537_inst_req_0 : boolean;
  signal binary_978_inst_ack_1 : boolean;
  signal simple_obj_ref_537_inst_ack_0 : boolean;
  signal ptr_deref_960_addr_0_ack_1 : boolean;
  signal binary_983_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal binary_983_inst_req_1 : boolean;
  signal ptr_deref_960_addr_2_req_0 : boolean;
  signal ptr_deref_960_gather_scatter_req_0 : boolean;
  signal ptr_deref_960_addr_1_req_0 : boolean;
  signal type_cast_542_inst_req_0 : boolean;
  signal type_cast_542_inst_ack_0 : boolean;
  signal array_obj_ref_549_base_resize_req_0 : boolean;
  signal array_obj_ref_549_base_resize_ack_0 : boolean;
  signal array_obj_ref_549_root_address_inst_req_0 : boolean;
  signal array_obj_ref_549_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_549_root_address_inst_req_1 : boolean;
  signal array_obj_ref_549_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_549_final_reg_req_0 : boolean;
  signal array_obj_ref_549_final_reg_ack_0 : boolean;
  signal ptr_deref_553_base_resize_req_0 : boolean;
  signal ptr_deref_553_base_resize_ack_0 : boolean;
  signal ptr_deref_553_root_address_inst_req_0 : boolean;
  signal ptr_deref_553_root_address_inst_ack_0 : boolean;
  signal ptr_deref_553_addr_0_req_0 : boolean;
  signal ptr_deref_553_addr_0_ack_0 : boolean;
  signal ptr_deref_553_addr_0_req_1 : boolean;
  signal ptr_deref_553_addr_0_ack_1 : boolean;
  signal ptr_deref_553_addr_1_req_0 : boolean;
  signal ptr_deref_553_addr_1_ack_0 : boolean;
  signal ptr_deref_553_addr_1_req_1 : boolean;
  signal ptr_deref_553_addr_1_ack_1 : boolean;
  signal ptr_deref_553_addr_2_req_0 : boolean;
  signal ptr_deref_553_addr_2_ack_0 : boolean;
  signal ptr_deref_553_addr_2_req_1 : boolean;
  signal ptr_deref_553_addr_2_ack_1 : boolean;
  signal ptr_deref_553_addr_3_req_0 : boolean;
  signal ptr_deref_553_addr_3_ack_0 : boolean;
  signal ptr_deref_553_addr_3_req_1 : boolean;
  signal ptr_deref_553_addr_3_ack_1 : boolean;
  signal ptr_deref_553_load_0_req_0 : boolean;
  signal ptr_deref_553_load_0_ack_0 : boolean;
  signal ptr_deref_553_load_1_req_0 : boolean;
  signal ptr_deref_553_load_1_ack_0 : boolean;
  signal ptr_deref_553_load_2_req_0 : boolean;
  signal ptr_deref_553_load_2_ack_0 : boolean;
  signal ptr_deref_553_load_3_req_0 : boolean;
  signal ptr_deref_553_load_3_ack_0 : boolean;
  signal ptr_deref_553_load_0_req_1 : boolean;
  signal ptr_deref_553_load_0_ack_1 : boolean;
  signal ptr_deref_553_load_1_req_1 : boolean;
  signal ptr_deref_553_load_1_ack_1 : boolean;
  signal ptr_deref_553_load_2_req_1 : boolean;
  signal ptr_deref_553_load_2_ack_1 : boolean;
  signal ptr_deref_553_load_3_req_1 : boolean;
  signal ptr_deref_553_load_3_ack_1 : boolean;
  signal ptr_deref_553_gather_scatter_req_0 : boolean;
  signal ptr_deref_553_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_558_base_resize_req_0 : boolean;
  signal array_obj_ref_558_base_resize_ack_0 : boolean;
  signal array_obj_ref_558_root_address_inst_req_0 : boolean;
  signal array_obj_ref_558_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_558_root_address_inst_req_1 : boolean;
  signal array_obj_ref_558_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_558_final_reg_req_0 : boolean;
  signal array_obj_ref_558_final_reg_ack_0 : boolean;
  signal array_obj_ref_565_base_resize_req_0 : boolean;
  signal array_obj_ref_565_base_resize_ack_0 : boolean;
  signal array_obj_ref_565_root_address_inst_req_0 : boolean;
  signal array_obj_ref_565_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_565_root_address_inst_req_1 : boolean;
  signal array_obj_ref_565_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_565_final_reg_req_0 : boolean;
  signal array_obj_ref_565_final_reg_ack_0 : boolean;
  signal ptr_deref_569_base_resize_req_0 : boolean;
  signal ptr_deref_569_base_resize_ack_0 : boolean;
  signal ptr_deref_569_root_address_inst_req_0 : boolean;
  signal ptr_deref_569_root_address_inst_ack_0 : boolean;
  signal ptr_deref_569_addr_0_req_0 : boolean;
  signal ptr_deref_569_addr_0_ack_0 : boolean;
  signal ptr_deref_569_addr_0_req_1 : boolean;
  signal ptr_deref_569_addr_0_ack_1 : boolean;
  signal ptr_deref_569_addr_1_req_0 : boolean;
  signal ptr_deref_569_addr_1_ack_0 : boolean;
  signal ptr_deref_569_addr_1_req_1 : boolean;
  signal ptr_deref_569_addr_1_ack_1 : boolean;
  signal ptr_deref_569_addr_2_req_0 : boolean;
  signal ptr_deref_569_addr_2_ack_0 : boolean;
  signal ptr_deref_569_addr_2_req_1 : boolean;
  signal ptr_deref_569_addr_2_ack_1 : boolean;
  signal ptr_deref_569_addr_3_req_0 : boolean;
  signal ptr_deref_569_addr_3_ack_0 : boolean;
  signal ptr_deref_569_addr_3_req_1 : boolean;
  signal ptr_deref_569_addr_3_ack_1 : boolean;
  signal phi_stmt_741_req_1 : boolean;
  signal binary_695_inst_req_0 : boolean;
  signal binary_695_inst_ack_0 : boolean;
  signal ptr_deref_1060_gather_scatter_ack_0 : boolean;
  signal binary_695_inst_req_1 : boolean;
  signal binary_695_inst_ack_1 : boolean;
  signal binary_700_inst_req_0 : boolean;
  signal binary_700_inst_ack_0 : boolean;
  signal ptr_deref_1060_store_0_req_0 : boolean;
  signal binary_700_inst_req_1 : boolean;
  signal binary_700_inst_ack_1 : boolean;
  signal ptr_deref_1060_store_3_ack_1 : boolean;
  signal phi_stmt_875_ack_0 : boolean;
  signal if_stmt_702_branch_req_0 : boolean;
  signal if_stmt_702_branch_ack_1 : boolean;
  signal if_stmt_702_branch_ack_0 : boolean;
  signal phi_stmt_734_req_0 : boolean;
  signal ptr_deref_1060_store_0_ack_0 : boolean;
  signal call_stmt_710_call_req_0 : boolean;
  signal call_stmt_710_call_ack_0 : boolean;
  signal call_stmt_710_call_req_1 : boolean;
  signal call_stmt_710_call_ack_1 : boolean;
  signal binary_717_inst_req_0 : boolean;
  signal binary_717_inst_ack_0 : boolean;
  signal binary_717_inst_req_1 : boolean;
  signal ptr_deref_1060_store_1_req_0 : boolean;
  signal binary_717_inst_ack_1 : boolean;
  signal if_stmt_719_branch_req_0 : boolean;
  signal type_cast_1078_inst_req_0 : boolean;
  signal if_stmt_719_branch_ack_1 : boolean;
  signal if_stmt_719_branch_ack_0 : boolean;
  signal ptr_deref_1060_store_1_ack_0 : boolean;
  signal phi_stmt_741_req_0 : boolean;
  signal ptr_deref_1060_store_2_req_0 : boolean;
  signal binary_730_inst_req_0 : boolean;
  signal binary_730_inst_ack_0 : boolean;
  signal binary_730_inst_req_1 : boolean;
  signal ptr_deref_1060_store_2_ack_0 : boolean;
  signal binary_730_inst_ack_1 : boolean;
  signal phi_stmt_734_ack_0 : boolean;
  signal phi_stmt_741_ack_0 : boolean;
  signal type_cast_1078_inst_ack_0 : boolean;
  signal binary_753_inst_req_0 : boolean;
  signal binary_753_inst_ack_0 : boolean;
  signal binary_753_inst_req_1 : boolean;
  signal type_cast_830_inst_req_0 : boolean;
  signal binary_753_inst_ack_1 : boolean;
  signal ptr_deref_1060_store_3_req_0 : boolean;
  signal type_cast_830_inst_ack_0 : boolean;
  signal ptr_deref_1060_store_3_ack_0 : boolean;
  signal type_cast_878_inst_req_0 : boolean;
  signal binary_758_inst_req_0 : boolean;
  signal binary_758_inst_ack_0 : boolean;
  signal binary_758_inst_req_1 : boolean;
  signal binary_758_inst_ack_1 : boolean;
  signal type_cast_1082_inst_req_0 : boolean;
  signal phi_stmt_827_req_0 : boolean;
  signal type_cast_1082_inst_ack_0 : boolean;
  signal binary_764_inst_req_0 : boolean;
  signal binary_764_inst_ack_0 : boolean;
  signal binary_764_inst_req_1 : boolean;
  signal binary_764_inst_ack_1 : boolean;
  signal type_cast_880_inst_req_0 : boolean;
  signal phi_stmt_840_req_0 : boolean;
  signal binary_770_inst_req_0 : boolean;
  signal binary_770_inst_ack_0 : boolean;
  signal binary_770_inst_req_1 : boolean;
  signal binary_770_inst_ack_1 : boolean;
  signal array_obj_ref_774_index_0_resize_req_0 : boolean;
  signal array_obj_ref_774_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_774_index_0_rename_req_0 : boolean;
  signal phi_stmt_827_req_1 : boolean;
  signal array_obj_ref_774_index_0_rename_ack_0 : boolean;
  signal type_cast_880_inst_ack_0 : boolean;
  signal ptr_deref_1060_store_0_req_1 : boolean;
  signal array_obj_ref_774_offset_inst_req_0 : boolean;
  signal array_obj_ref_774_offset_inst_ack_0 : boolean;
  signal simple_obj_ref_1080_inst_req_0 : boolean;
  signal array_obj_ref_774_base_resize_req_0 : boolean;
  signal array_obj_ref_774_base_resize_ack_0 : boolean;
  signal ptr_deref_1060_store_0_ack_1 : boolean;
  signal simple_obj_ref_1080_inst_ack_0 : boolean;
  signal array_obj_ref_774_root_address_inst_req_0 : boolean;
  signal array_obj_ref_774_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_774_root_address_inst_req_1 : boolean;
  signal array_obj_ref_774_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_774_final_reg_req_0 : boolean;
  signal array_obj_ref_774_final_reg_ack_0 : boolean;
  signal type_cast_878_inst_ack_0 : boolean;
  signal type_cast_779_inst_req_0 : boolean;
  signal type_cast_779_inst_ack_0 : boolean;
  signal type_cast_837_inst_req_0 : boolean;
  signal ptr_deref_783_base_resize_req_0 : boolean;
  signal ptr_deref_783_base_resize_ack_0 : boolean;
  signal type_cast_837_inst_ack_0 : boolean;
  signal ptr_deref_783_root_address_inst_req_0 : boolean;
  signal ptr_deref_783_root_address_inst_ack_0 : boolean;
  signal ptr_deref_783_addr_0_req_0 : boolean;
  signal ptr_deref_783_addr_0_ack_0 : boolean;
  signal type_cast_839_inst_req_0 : boolean;
  signal ptr_deref_783_addr_0_req_1 : boolean;
  signal ptr_deref_783_addr_0_ack_1 : boolean;
  signal ptr_deref_783_addr_1_req_0 : boolean;
  signal ptr_deref_783_addr_1_ack_0 : boolean;
  signal type_cast_839_inst_ack_0 : boolean;
  signal ptr_deref_783_addr_1_req_1 : boolean;
  signal ptr_deref_1060_store_1_req_1 : boolean;
  signal ptr_deref_783_addr_1_ack_1 : boolean;
  signal ptr_deref_1060_store_1_ack_1 : boolean;
  signal ptr_deref_783_load_0_req_0 : boolean;
  signal ptr_deref_783_load_0_ack_0 : boolean;
  signal ptr_deref_783_load_1_req_0 : boolean;
  signal phi_stmt_834_req_1 : boolean;
  signal ptr_deref_783_load_1_ack_0 : boolean;
  signal ptr_deref_783_load_0_req_1 : boolean;
  signal ptr_deref_783_load_0_ack_1 : boolean;
  signal ptr_deref_783_load_1_req_1 : boolean;
  signal ptr_deref_783_load_1_ack_1 : boolean;
  signal ptr_deref_783_gather_scatter_req_0 : boolean;
  signal ptr_deref_783_gather_scatter_ack_0 : boolean;
  signal phi_stmt_827_ack_0 : boolean;
  signal type_cast_787_inst_req_0 : boolean;
  signal type_cast_787_inst_ack_0 : boolean;
  signal phi_stmt_834_req_0 : boolean;
  signal phi_stmt_875_req_0 : boolean;
  signal ptr_deref_1060_store_2_req_1 : boolean;
  signal phi_stmt_875_req_1 : boolean;
  signal binary_792_inst_req_0 : boolean;
  signal binary_792_inst_ack_0 : boolean;
  signal ptr_deref_1060_store_2_ack_1 : boolean;
  signal binary_792_inst_req_1 : boolean;
  signal binary_792_inst_ack_1 : boolean;
  signal type_cast_796_inst_req_0 : boolean;
  signal type_cast_796_inst_ack_0 : boolean;
  signal binary_800_inst_req_0 : boolean;
  signal binary_800_inst_ack_0 : boolean;
  signal binary_800_inst_req_1 : boolean;
  signal binary_800_inst_ack_1 : boolean;
  signal binary_806_inst_req_0 : boolean;
  signal binary_806_inst_ack_0 : boolean;
  signal binary_806_inst_req_1 : boolean;
  signal binary_806_inst_ack_1 : boolean;
  signal if_stmt_808_branch_req_0 : boolean;
  signal if_stmt_808_branch_ack_1 : boolean;
  signal if_stmt_808_branch_ack_0 : boolean;
  signal binary_819_inst_req_0 : boolean;
  signal binary_819_inst_ack_0 : boolean;
  signal binary_819_inst_req_1 : boolean;
  signal binary_819_inst_ack_1 : boolean;
  signal array_obj_ref_823_index_0_resize_req_0 : boolean;
  signal array_obj_ref_823_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_823_index_0_rename_req_0 : boolean;
  signal array_obj_ref_823_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_823_offset_inst_req_0 : boolean;
  signal array_obj_ref_823_offset_inst_ack_0 : boolean;
  signal array_obj_ref_823_base_resize_req_0 : boolean;
  signal array_obj_ref_823_base_resize_ack_0 : boolean;
  signal array_obj_ref_823_root_address_inst_req_0 : boolean;
  signal array_obj_ref_823_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_823_root_address_inst_req_1 : boolean;
  signal array_obj_ref_823_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_823_final_reg_req_0 : boolean;
  signal array_obj_ref_823_final_reg_ack_0 : boolean;
  signal binary_851_inst_req_0 : boolean;
  signal binary_851_inst_ack_0 : boolean;
  signal binary_851_inst_req_1 : boolean;
  signal binary_851_inst_ack_1 : boolean;
  signal if_stmt_853_branch_req_0 : boolean;
  signal if_stmt_853_branch_ack_1 : boolean;
  signal if_stmt_853_branch_ack_0 : boolean;
  signal ptr_deref_862_base_resize_req_0 : boolean;
  signal ptr_deref_862_base_resize_ack_0 : boolean;
  signal ptr_deref_862_root_address_inst_req_0 : boolean;
  signal ptr_deref_862_root_address_inst_ack_0 : boolean;
  signal ptr_deref_862_addr_0_req_0 : boolean;
  signal ptr_deref_862_addr_0_ack_0 : boolean;
  signal ptr_deref_862_load_0_req_0 : boolean;
  signal ptr_deref_862_load_0_ack_0 : boolean;
  signal ptr_deref_862_load_0_req_1 : boolean;
  signal ptr_deref_862_load_0_ack_1 : boolean;
  signal ptr_deref_862_gather_scatter_req_0 : boolean;
  signal ptr_deref_862_gather_scatter_ack_0 : boolean;
  signal type_cast_866_inst_req_0 : boolean;
  signal type_cast_866_inst_ack_0 : boolean;
  signal binary_871_inst_req_0 : boolean;
  signal binary_871_inst_ack_0 : boolean;
  signal binary_871_inst_req_1 : boolean;
  signal binary_871_inst_ack_1 : boolean;
  signal binary_886_inst_req_0 : boolean;
  signal binary_886_inst_ack_0 : boolean;
  signal binary_886_inst_req_1 : boolean;
  signal binary_886_inst_ack_1 : boolean;
  signal binary_892_inst_req_0 : boolean;
  signal binary_892_inst_ack_0 : boolean;
  signal binary_892_inst_req_1 : boolean;
  signal binary_892_inst_ack_1 : boolean;
  signal binary_897_inst_req_0 : boolean;
  signal binary_897_inst_ack_0 : boolean;
  signal binary_897_inst_req_1 : boolean;
  signal binary_897_inst_ack_1 : boolean;
  signal binary_903_inst_req_0 : boolean;
  signal binary_903_inst_ack_0 : boolean;
  signal binary_903_inst_req_1 : boolean;
  signal binary_903_inst_ack_1 : boolean;
  signal binary_908_inst_req_0 : boolean;
  signal binary_908_inst_ack_0 : boolean;
  signal binary_908_inst_req_1 : boolean;
  signal binary_908_inst_ack_1 : boolean;
  signal type_cast_912_inst_req_0 : boolean;
  signal type_cast_912_inst_ack_0 : boolean;
  signal binary_918_inst_req_0 : boolean;
  signal binary_918_inst_ack_0 : boolean;
  signal binary_918_inst_req_1 : boolean;
  signal binary_918_inst_ack_1 : boolean;
  signal if_stmt_920_branch_req_0 : boolean;
  signal if_stmt_920_branch_ack_1 : boolean;
  signal if_stmt_920_branch_ack_0 : boolean;
  signal call_stmt_928_call_req_0 : boolean;
  signal call_stmt_928_call_ack_0 : boolean;
  signal call_stmt_928_call_req_1 : boolean;
  signal call_stmt_928_call_ack_1 : boolean;
  signal array_obj_ref_936_base_resize_req_0 : boolean;
  signal array_obj_ref_936_base_resize_ack_0 : boolean;
  signal array_obj_ref_936_root_address_inst_req_0 : boolean;
  signal array_obj_ref_936_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_936_root_address_inst_req_1 : boolean;
  signal array_obj_ref_936_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_936_final_reg_req_0 : boolean;
  signal array_obj_ref_936_final_reg_ack_0 : boolean;
  signal ptr_deref_939_base_resize_req_0 : boolean;
  signal ptr_deref_939_base_resize_ack_0 : boolean;
  signal ptr_deref_939_root_address_inst_req_0 : boolean;
  signal ptr_deref_939_root_address_inst_ack_0 : boolean;
  signal ptr_deref_939_addr_0_req_0 : boolean;
  signal ptr_deref_939_addr_0_ack_0 : boolean;
  signal ptr_deref_939_addr_0_req_1 : boolean;
  signal ptr_deref_939_addr_0_ack_1 : boolean;
  signal ptr_deref_939_addr_1_req_0 : boolean;
  signal ptr_deref_939_addr_1_ack_0 : boolean;
  signal ptr_deref_939_addr_1_req_1 : boolean;
  signal ptr_deref_939_addr_1_ack_1 : boolean;
  signal ptr_deref_939_addr_2_req_0 : boolean;
  signal ptr_deref_939_addr_2_ack_0 : boolean;
  signal ptr_deref_939_addr_2_req_1 : boolean;
  signal ptr_deref_939_addr_2_ack_1 : boolean;
  signal ptr_deref_939_addr_3_req_0 : boolean;
  signal ptr_deref_939_addr_3_ack_0 : boolean;
  signal ptr_deref_939_addr_3_req_1 : boolean;
  signal ptr_deref_939_addr_3_ack_1 : boolean;
  signal ptr_deref_939_gather_scatter_req_0 : boolean;
  signal ptr_deref_939_gather_scatter_ack_0 : boolean;
  signal ptr_deref_939_store_0_req_0 : boolean;
  signal ptr_deref_939_store_0_ack_0 : boolean;
  signal ptr_deref_939_store_1_req_0 : boolean;
  signal ptr_deref_939_store_1_ack_0 : boolean;
  signal ptr_deref_939_store_2_req_0 : boolean;
  signal ptr_deref_939_store_2_ack_0 : boolean;
  signal ptr_deref_939_store_3_req_0 : boolean;
  signal ptr_deref_939_store_3_ack_0 : boolean;
  signal ptr_deref_939_store_0_req_1 : boolean;
  signal ptr_deref_939_store_0_ack_1 : boolean;
  signal ptr_deref_939_store_1_req_1 : boolean;
  signal ptr_deref_939_store_1_ack_1 : boolean;
  signal ptr_deref_939_store_2_req_1 : boolean;
  signal ptr_deref_939_store_2_ack_1 : boolean;
  signal ptr_deref_939_store_3_req_1 : boolean;
  signal ptr_deref_939_store_3_ack_1 : boolean;
  signal binary_946_inst_req_0 : boolean;
  signal binary_946_inst_ack_0 : boolean;
  signal binary_946_inst_req_1 : boolean;
  signal binary_946_inst_ack_1 : boolean;
  signal array_obj_ref_950_index_0_resize_req_0 : boolean;
  signal array_obj_ref_950_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_950_index_0_rename_req_0 : boolean;
  signal array_obj_ref_950_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_950_offset_inst_req_0 : boolean;
  signal array_obj_ref_950_offset_inst_ack_0 : boolean;
  signal array_obj_ref_950_base_resize_req_0 : boolean;
  signal array_obj_ref_950_base_resize_ack_0 : boolean;
  signal array_obj_ref_950_root_address_inst_req_0 : boolean;
  signal array_obj_ref_950_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_950_root_address_inst_req_1 : boolean;
  signal array_obj_ref_950_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_950_final_reg_req_0 : boolean;
  signal array_obj_ref_950_final_reg_ack_0 : boolean;
  signal array_obj_ref_957_base_resize_req_0 : boolean;
  signal array_obj_ref_957_base_resize_ack_0 : boolean;
  signal array_obj_ref_957_root_address_inst_req_0 : boolean;
  signal array_obj_ref_957_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_957_root_address_inst_req_1 : boolean;
  signal array_obj_ref_957_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_957_final_reg_req_0 : boolean;
  signal array_obj_ref_957_final_reg_ack_0 : boolean;
  signal array_obj_ref_999_index_0_resize_req_0 : boolean;
  signal array_obj_ref_999_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_999_index_0_rename_req_0 : boolean;
  signal array_obj_ref_999_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_999_offset_inst_req_0 : boolean;
  signal array_obj_ref_999_offset_inst_ack_0 : boolean;
  signal array_obj_ref_999_base_resize_req_0 : boolean;
  signal array_obj_ref_999_base_resize_ack_0 : boolean;
  signal array_obj_ref_999_root_address_inst_req_0 : boolean;
  signal array_obj_ref_999_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_999_root_address_inst_req_1 : boolean;
  signal array_obj_ref_999_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_999_final_reg_req_0 : boolean;
  signal array_obj_ref_999_final_reg_ack_0 : boolean;
  signal ptr_deref_1002_base_resize_req_0 : boolean;
  signal ptr_deref_1002_base_resize_ack_0 : boolean;
  signal ptr_deref_1002_root_address_inst_req_0 : boolean;
  signal ptr_deref_1002_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1002_addr_0_req_0 : boolean;
  signal ptr_deref_1002_addr_0_ack_0 : boolean;
  signal ptr_deref_1002_addr_0_req_1 : boolean;
  signal ptr_deref_1002_addr_0_ack_1 : boolean;
  signal ptr_deref_1002_addr_1_req_0 : boolean;
  signal ptr_deref_1002_addr_1_ack_0 : boolean;
  signal ptr_deref_1002_addr_1_req_1 : boolean;
  signal ptr_deref_1002_addr_1_ack_1 : boolean;
  signal ptr_deref_1002_addr_2_req_0 : boolean;
  signal ptr_deref_1002_addr_2_ack_0 : boolean;
  signal ptr_deref_1002_addr_2_req_1 : boolean;
  signal ptr_deref_1002_addr_2_ack_1 : boolean;
  signal ptr_deref_1002_addr_3_req_0 : boolean;
  signal ptr_deref_1002_addr_3_ack_0 : boolean;
  signal ptr_deref_1002_addr_3_req_1 : boolean;
  signal ptr_deref_1002_addr_3_ack_1 : boolean;
  signal ptr_deref_1002_gather_scatter_req_0 : boolean;
  signal ptr_deref_1002_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1002_store_0_req_0 : boolean;
  signal ptr_deref_1002_store_0_ack_0 : boolean;
  signal ptr_deref_1002_store_1_req_0 : boolean;
  signal ptr_deref_1002_store_1_ack_0 : boolean;
  signal ptr_deref_1002_store_2_req_0 : boolean;
  signal ptr_deref_1002_store_2_ack_0 : boolean;
  signal ptr_deref_1002_store_3_req_0 : boolean;
  signal ptr_deref_1002_store_3_ack_0 : boolean;
  signal ptr_deref_1002_store_0_req_1 : boolean;
  signal ptr_deref_1002_store_0_ack_1 : boolean;
  signal ptr_deref_1002_store_1_req_1 : boolean;
  signal ptr_deref_1002_store_1_ack_1 : boolean;
  signal ptr_deref_1002_store_2_req_1 : boolean;
  signal ptr_deref_1002_store_2_ack_1 : boolean;
  signal ptr_deref_1002_store_3_req_1 : boolean;
  signal ptr_deref_1002_store_3_ack_1 : boolean;
  signal array_obj_ref_1008_base_resize_req_0 : boolean;
  signal array_obj_ref_1008_base_resize_ack_0 : boolean;
  signal array_obj_ref_1008_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1008_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1008_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1008_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1008_final_reg_req_0 : boolean;
  signal array_obj_ref_1008_final_reg_ack_0 : boolean;
  signal type_cast_1012_inst_req_0 : boolean;
  signal type_cast_1012_inst_ack_0 : boolean;
  signal ptr_deref_1016_base_resize_req_0 : boolean;
  signal ptr_deref_1016_base_resize_ack_0 : boolean;
  signal ptr_deref_1016_root_address_inst_req_0 : boolean;
  signal ptr_deref_1016_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1016_addr_0_req_0 : boolean;
  signal ptr_deref_1016_addr_0_ack_0 : boolean;
  signal ptr_deref_1016_addr_0_req_1 : boolean;
  signal ptr_deref_1016_addr_0_ack_1 : boolean;
  signal ptr_deref_1016_addr_1_req_0 : boolean;
  signal ptr_deref_1016_addr_1_ack_0 : boolean;
  signal ptr_deref_1016_addr_1_req_1 : boolean;
  signal ptr_deref_1016_addr_1_ack_1 : boolean;
  signal ptr_deref_1016_addr_2_req_0 : boolean;
  signal ptr_deref_1016_addr_2_ack_0 : boolean;
  signal ptr_deref_1016_addr_2_req_1 : boolean;
  signal ptr_deref_1016_addr_2_ack_1 : boolean;
  signal ptr_deref_1016_addr_3_req_0 : boolean;
  signal ptr_deref_1016_addr_3_ack_0 : boolean;
  signal ptr_deref_1016_addr_3_req_1 : boolean;
  signal ptr_deref_1016_addr_3_ack_1 : boolean;
  signal ptr_deref_1016_load_0_req_0 : boolean;
  signal ptr_deref_1016_load_0_ack_0 : boolean;
  signal ptr_deref_1016_load_1_req_0 : boolean;
  signal ptr_deref_1016_load_1_ack_0 : boolean;
  signal ptr_deref_1016_load_2_req_0 : boolean;
  signal ptr_deref_1016_load_2_ack_0 : boolean;
  signal ptr_deref_1016_load_3_req_0 : boolean;
  signal ptr_deref_1016_load_3_ack_0 : boolean;
  signal ptr_deref_1016_load_0_req_1 : boolean;
  signal ptr_deref_1016_load_0_ack_1 : boolean;
  signal ptr_deref_1016_load_1_req_1 : boolean;
  signal ptr_deref_1016_load_1_ack_1 : boolean;
  signal ptr_deref_1016_load_2_req_1 : boolean;
  signal ptr_deref_1016_load_2_ack_1 : boolean;
  signal ptr_deref_1016_load_3_req_1 : boolean;
  signal ptr_deref_1016_load_3_ack_1 : boolean;
  signal ptr_deref_1016_gather_scatter_req_0 : boolean;
  signal ptr_deref_1016_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1023_base_resize_req_0 : boolean;
  signal array_obj_ref_1023_base_resize_ack_0 : boolean;
  signal array_obj_ref_1023_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1023_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1023_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1023_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1023_final_reg_req_0 : boolean;
  signal array_obj_ref_1023_final_reg_ack_0 : boolean;
  signal type_cast_1027_inst_req_0 : boolean;
  signal type_cast_1027_inst_ack_0 : boolean;
  signal ptr_deref_1030_base_resize_req_0 : boolean;
  signal ptr_deref_1030_base_resize_ack_0 : boolean;
  signal ptr_deref_1030_root_address_inst_req_0 : boolean;
  signal ptr_deref_1030_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1030_addr_0_req_0 : boolean;
  signal ptr_deref_1030_addr_0_ack_0 : boolean;
  signal ptr_deref_1030_addr_0_req_1 : boolean;
  signal ptr_deref_1030_addr_0_ack_1 : boolean;
  signal ptr_deref_1030_addr_1_req_0 : boolean;
  signal ptr_deref_1030_addr_1_ack_0 : boolean;
  signal ptr_deref_1030_addr_1_req_1 : boolean;
  signal ptr_deref_1030_addr_1_ack_1 : boolean;
  signal ptr_deref_1030_addr_2_req_0 : boolean;
  signal ptr_deref_1030_addr_2_ack_0 : boolean;
  signal ptr_deref_1030_addr_2_req_1 : boolean;
  signal ptr_deref_1030_addr_2_ack_1 : boolean;
  signal ptr_deref_1030_addr_3_req_0 : boolean;
  signal ptr_deref_1030_addr_3_ack_0 : boolean;
  signal ptr_deref_1030_addr_3_req_1 : boolean;
  signal ptr_deref_1030_addr_3_ack_1 : boolean;
  signal ptr_deref_1030_gather_scatter_req_0 : boolean;
  signal ptr_deref_1030_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1030_store_0_req_0 : boolean;
  signal ptr_deref_1030_store_0_ack_0 : boolean;
  signal ptr_deref_1030_store_1_req_0 : boolean;
  signal ptr_deref_1030_store_1_ack_0 : boolean;
  signal ptr_deref_1030_store_2_req_0 : boolean;
  signal ptr_deref_1030_store_2_ack_0 : boolean;
  signal ptr_deref_1030_store_3_req_0 : boolean;
  signal ptr_deref_1030_store_3_ack_0 : boolean;
  signal ptr_deref_1030_store_0_req_1 : boolean;
  signal ptr_deref_1030_store_0_ack_1 : boolean;
  signal ptr_deref_1030_store_1_req_1 : boolean;
  signal ptr_deref_1030_store_1_ack_1 : boolean;
  signal ptr_deref_1030_store_2_req_1 : boolean;
  signal ptr_deref_1030_store_2_ack_1 : boolean;
  signal ptr_deref_1030_store_3_req_1 : boolean;
  signal ptr_deref_1030_store_3_ack_1 : boolean;
  signal array_obj_ref_1038_base_resize_req_0 : boolean;
  signal array_obj_ref_1038_base_resize_ack_0 : boolean;
  signal array_obj_ref_1038_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1038_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1038_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1038_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1038_final_reg_req_0 : boolean;
  signal array_obj_ref_1038_final_reg_ack_0 : boolean;
  signal type_cast_1042_inst_req_0 : boolean;
  signal type_cast_1042_inst_ack_0 : boolean;
  signal ptr_deref_1046_base_resize_req_0 : boolean;
  signal ptr_deref_1046_base_resize_ack_0 : boolean;
  signal ptr_deref_1046_root_address_inst_req_0 : boolean;
  signal ptr_deref_1046_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1046_addr_0_req_0 : boolean;
  signal ptr_deref_1046_addr_0_ack_0 : boolean;
  signal ptr_deref_1046_addr_0_req_1 : boolean;
  signal ptr_deref_1046_addr_0_ack_1 : boolean;
  signal ptr_deref_1046_addr_1_req_0 : boolean;
  signal ptr_deref_1046_addr_1_ack_0 : boolean;
  signal ptr_deref_1046_addr_1_req_1 : boolean;
  signal ptr_deref_1046_addr_1_ack_1 : boolean;
  signal ptr_deref_1046_addr_2_req_0 : boolean;
  signal ptr_deref_1046_addr_2_ack_0 : boolean;
  signal ptr_deref_1046_addr_2_req_1 : boolean;
  signal ptr_deref_1046_addr_2_ack_1 : boolean;
  signal ptr_deref_1046_addr_3_req_0 : boolean;
  signal ptr_deref_1046_addr_3_ack_0 : boolean;
  signal ptr_deref_1046_addr_3_req_1 : boolean;
  signal ptr_deref_1046_addr_3_ack_1 : boolean;
  signal ptr_deref_1046_load_0_req_0 : boolean;
  signal ptr_deref_1046_load_0_ack_0 : boolean;
  signal ptr_deref_1046_load_1_req_0 : boolean;
  signal ptr_deref_1046_load_1_ack_0 : boolean;
  signal ptr_deref_1046_load_2_req_0 : boolean;
  signal ptr_deref_1046_load_2_ack_0 : boolean;
  signal ptr_deref_1046_load_3_req_0 : boolean;
  signal ptr_deref_1046_load_3_ack_0 : boolean;
  signal ptr_deref_1046_load_0_req_1 : boolean;
  signal ptr_deref_1046_load_0_ack_1 : boolean;
  signal ptr_deref_1046_load_1_req_1 : boolean;
  signal ptr_deref_1046_load_1_ack_1 : boolean;
  signal ptr_deref_1046_load_2_req_1 : boolean;
  signal ptr_deref_1046_load_2_ack_1 : boolean;
  signal ptr_deref_1046_load_3_req_1 : boolean;
  signal ptr_deref_1046_load_3_ack_1 : boolean;
  signal ptr_deref_1046_gather_scatter_req_0 : boolean;
  signal ptr_deref_1046_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1053_base_resize_req_0 : boolean;
  signal array_obj_ref_1053_base_resize_ack_0 : boolean;
  signal array_obj_ref_1053_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1053_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1053_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1053_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1053_final_reg_req_0 : boolean;
  signal array_obj_ref_1053_final_reg_ack_0 : boolean;
  signal type_cast_1057_inst_req_0 : boolean;
  signal type_cast_1057_inst_ack_0 : boolean;
  signal ptr_deref_1060_base_resize_req_0 : boolean;
  signal ptr_deref_1060_base_resize_ack_0 : boolean;
  signal ptr_deref_1060_root_address_inst_req_0 : boolean;
  signal ptr_deref_1060_root_address_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_chk_CP_1053: Block -- control-path 
    signal cp_elements: BooleanArray(974 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(974);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(974), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(145);
    cp_elements(2) <= OrReduce(cp_elements(152) & cp_elements(893));
    crr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_607_call_req_0); -- 
    cp_elements(3) <= cp_elements(215);
    cp_elements(4) <= OrReduce(cp_elements(224) & cp_elements(895));
    crr_1775_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => call_stmt_648_call_req_0); -- 
    cp_elements(5) <= OrReduce(cp_elements(247) & cp_elements(897));
    crr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => call_stmt_677_call_req_0); -- 
    cp_elements(6) <= OrReduce(cp_elements(281) & cp_elements(899));
    crr_1958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => call_stmt_710_call_req_0); -- 
    cp_elements(7) <= OrReduce(cp_elements(298) & cp_elements(901));
    cp_elements(8) <= cp_elements(916);
    cp_elements(9) <= cp_elements(383);
    cp_elements(10) <= OrReduce(cp_elements(392) & cp_elements(918));
    cp_elements(11) <= cp_elements(951);
    cp_elements(12) <= OrReduce(cp_elements(422) & cp_elements(953));
    cp_elements(13) <= OrReduce(cp_elements(483) & cp_elements(966));
    crr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => call_stmt_928_call_req_0); -- 
    cp_elements(14) <= cp_elements(597);
    cp_elements(15) <= OrReduce(cp_elements(604) & cp_elements(968));
    cp_elements(16) <= cp_elements(771);
    cp_elements(17) <= cp_elements(871);
    cp_elements(18) <= OrReduce(cp_elements(970) & cp_elements(972));
    cp_elements(19) <= cp_elements(0);
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(21) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_538_inst_req_0); -- 
    cp_elements(21) <= cp_elements(19);
    cp_elements(22) <= cp_elements(19);
    req_1180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => simple_obj_ref_537_inst_req_0); -- 
    ack_1181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_537_inst_ack_0, ack => cp_elements(23)); -- 
    ack_1186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => cp_elements(24)); -- 
    cp_elements(25) <= cp_elements(24);
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(28));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => type_cast_542_inst_req_0); -- 
    cp_elements(27) <= cp_elements(25);
    cp_elements(28) <= cp_elements(25);
    cp_elements(29) <= type_cast_542_inst_ack_0;
    cp_elements(30) <= cp_elements(25);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(35));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_549_final_reg_req_0); -- 
    cp_elements(32) <= cp_elements(29);
    base_resize_req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_549_base_resize_req_0); -- 
    base_resize_ack_1211_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_base_resize_ack_0, ack => cp_elements(33)); -- 
    plus_base_rr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_549_root_address_inst_req_0); -- 
    plus_base_ra_1217_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_root_address_inst_ack_0, ack => cp_elements(34)); -- 
    plus_base_cr_1218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_549_root_address_inst_req_1); -- 
    plus_base_ca_1219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_root_address_inst_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= array_obj_ref_549_final_reg_ack_0;
    cpelement_group_37 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(36) & cp_elements(53));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(37),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(38) <= cp_elements(36);
    base_resize_req_1237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => ptr_deref_553_base_resize_req_0); -- 
    base_resize_ack_1238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_base_resize_ack_0, ack => cp_elements(39)); -- 
    sum_rename_req_1242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => ptr_deref_553_root_address_inst_req_0); -- 
    cp_elements(40) <= ptr_deref_553_root_address_inst_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_553_addr_0_req_0); -- 
    ra_1251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_0_ack_0, ack => cp_elements(42)); -- 
    cr_1252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_553_addr_0_req_1); -- 
    ca_1253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_0_ack_1, ack => cp_elements(43)); -- 
    cp_elements(44) <= cp_elements(40);
    rr_1257_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_553_addr_1_req_0); -- 
    ra_1258_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_1_ack_0, ack => cp_elements(45)); -- 
    cr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_553_addr_1_req_1); -- 
    ca_1260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_1_ack_1, ack => cp_elements(46)); -- 
    cp_elements(47) <= cp_elements(40);
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_553_addr_2_req_0); -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_2_ack_0, ack => cp_elements(48)); -- 
    cr_1266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_553_addr_2_req_1); -- 
    ca_1267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_2_ack_1, ack => cp_elements(49)); -- 
    cp_elements(50) <= cp_elements(40);
    rr_1271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => ptr_deref_553_addr_3_req_0); -- 
    ra_1272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_3_ack_0, ack => cp_elements(51)); -- 
    cr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => ptr_deref_553_addr_3_req_1); -- 
    ca_1274_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_3_ack_1, ack => cp_elements(52)); -- 
    cpelement_group_53 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(43) & cp_elements(46) & cp_elements(49) & cp_elements(52));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(53),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(54) <= cp_elements(37);
    rr_1284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_553_load_0_req_0); -- 
    ra_1285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_0_ack_0, ack => cp_elements(55)); -- 
    cp_elements(56) <= cp_elements(37);
    rr_1289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => ptr_deref_553_load_1_req_0); -- 
    ra_1290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_1_ack_0, ack => cp_elements(57)); -- 
    cp_elements(58) <= cp_elements(37);
    rr_1294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_553_load_2_req_0); -- 
    ra_1295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_2_ack_0, ack => cp_elements(59)); -- 
    cp_elements(60) <= cp_elements(37);
    rr_1299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => ptr_deref_553_load_3_req_0); -- 
    ra_1300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_3_ack_0, ack => cp_elements(61)); -- 
    cpelement_group_62 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(55) & cp_elements(57) & cp_elements(59) & cp_elements(61));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(62),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(63) <= cp_elements(62);
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_553_load_0_req_1); -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_0_ack_1, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(62);
    cr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_553_load_1_req_1); -- 
    ca_1316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_1_ack_1, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(62);
    cr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => ptr_deref_553_load_2_req_1); -- 
    ca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_2_ack_1, ack => cp_elements(68)); -- 
    cp_elements(69) <= cp_elements(62);
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_553_load_3_req_1); -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_3_ack_1, ack => cp_elements(70)); -- 
    cpelement_group_71 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66) & cp_elements(68) & cp_elements(70));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(71),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_1327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => ptr_deref_553_gather_scatter_req_0); -- 
    cp_elements(72) <= ptr_deref_553_gather_scatter_ack_0;
    cp_elements(73) <= cp_elements(25);
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(73) & cp_elements(78));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_558_final_reg_req_0); -- 
    cp_elements(75) <= cp_elements(72);
    base_resize_req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_558_base_resize_req_0); -- 
    base_resize_ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_base_resize_ack_0, ack => cp_elements(76)); -- 
    plus_base_rr_1345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => array_obj_ref_558_root_address_inst_req_0); -- 
    plus_base_ra_1346_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_root_address_inst_ack_0, ack => cp_elements(77)); -- 
    plus_base_cr_1347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => array_obj_ref_558_root_address_inst_req_1); -- 
    plus_base_ca_1348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_root_address_inst_ack_1, ack => cp_elements(78)); -- 
    final_reg_ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_final_reg_ack_0, ack => cp_elements(79)); -- 
    cp_elements(80) <= cp_elements(25);
    cpelement_group_81 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(80) & cp_elements(85));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(81),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_565_final_reg_req_0); -- 
    cp_elements(82) <= cp_elements(29);
    base_resize_req_1364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_565_base_resize_req_0); -- 
    base_resize_ack_1365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_base_resize_ack_0, ack => cp_elements(83)); -- 
    plus_base_rr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => array_obj_ref_565_root_address_inst_req_0); -- 
    plus_base_ra_1371_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_root_address_inst_ack_0, ack => cp_elements(84)); -- 
    plus_base_cr_1372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => array_obj_ref_565_root_address_inst_req_1); -- 
    plus_base_ca_1373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_root_address_inst_ack_1, ack => cp_elements(85)); -- 
    cp_elements(86) <= array_obj_ref_565_final_reg_ack_0;
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(86) & cp_elements(103));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(88) <= cp_elements(86);
    base_resize_req_1391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_569_base_resize_req_0); -- 
    base_resize_ack_1392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_base_resize_ack_0, ack => cp_elements(89)); -- 
    sum_rename_req_1396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_569_root_address_inst_req_0); -- 
    cp_elements(90) <= ptr_deref_569_root_address_inst_ack_0;
    cp_elements(91) <= cp_elements(90);
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => ptr_deref_569_addr_0_req_0); -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_0_ack_0, ack => cp_elements(92)); -- 
    cr_1406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_569_addr_0_req_1); -- 
    ca_1407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_0_ack_1, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(90);
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_569_addr_1_req_0); -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_1_ack_0, ack => cp_elements(95)); -- 
    cr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => ptr_deref_569_addr_1_req_1); -- 
    ca_1414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_1_ack_1, ack => cp_elements(96)); -- 
    cp_elements(97) <= cp_elements(90);
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => ptr_deref_569_addr_2_req_0); -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_2_ack_0, ack => cp_elements(98)); -- 
    cr_1420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_569_addr_2_req_1); -- 
    ca_1421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_2_ack_1, ack => cp_elements(99)); -- 
    cp_elements(100) <= cp_elements(90);
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_569_addr_3_req_0); -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_3_ack_0, ack => cp_elements(101)); -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_569_addr_3_req_1); -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_3_ack_1, ack => cp_elements(102)); -- 
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(96) & cp_elements(99) & cp_elements(102));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(104) <= cp_elements(87);
    rr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_569_load_0_req_0); -- 
    ra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_0_ack_0, ack => cp_elements(105)); -- 
    cp_elements(106) <= cp_elements(87);
    rr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_569_load_1_req_0); -- 
    ra_1444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_1_ack_0, ack => cp_elements(107)); -- 
    cp_elements(108) <= cp_elements(87);
    rr_1448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => ptr_deref_569_load_2_req_0); -- 
    ra_1449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_2_ack_0, ack => cp_elements(109)); -- 
    cp_elements(110) <= cp_elements(87);
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ptr_deref_569_load_3_req_0); -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_3_ack_0, ack => cp_elements(111)); -- 
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(105) & cp_elements(107) & cp_elements(109) & cp_elements(111));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(113) <= cp_elements(112);
    cr_1464_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_569_load_0_req_1); -- 
    ca_1465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_0_ack_1, ack => cp_elements(114)); -- 
    cp_elements(115) <= cp_elements(112);
    cr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_569_load_1_req_1); -- 
    ca_1470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_1_ack_1, ack => cp_elements(116)); -- 
    cp_elements(117) <= cp_elements(112);
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_569_load_2_req_1); -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_2_ack_1, ack => cp_elements(118)); -- 
    cp_elements(119) <= cp_elements(112);
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_569_load_3_req_1); -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_3_ack_1, ack => cp_elements(120)); -- 
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(116) & cp_elements(118) & cp_elements(120));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_1481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => ptr_deref_569_gather_scatter_req_0); -- 
    merge_ack_1482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_gather_scatter_ack_0, ack => cp_elements(122)); -- 
    cpelement_group_123 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(122) & cp_elements(124));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(123),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1491_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => type_cast_573_inst_req_0); -- 
    cp_elements(124) <= cp_elements(25);
    ack_1492_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_0, ack => cp_elements(125)); -- 
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(128));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => type_cast_577_inst_req_0); -- 
    cp_elements(127) <= cp_elements(25);
    cp_elements(128) <= cp_elements(72);
    ack_1502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => cp_elements(129)); -- 
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(129) & cp_elements(131));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => binary_582_inst_req_0); -- 
    cp_elements(131) <= cp_elements(25);
    ra_1513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_582_inst_ack_0, ack => cp_elements(132)); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => binary_582_inst_req_1); -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_582_inst_ack_1, ack => cp_elements(133)); -- 
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(135));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => binary_588_inst_req_0); -- 
    cp_elements(135) <= cp_elements(25);
    ra_1525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_588_inst_ack_0, ack => cp_elements(136)); -- 
    cr_1526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => binary_588_inst_req_1); -- 
    ca_1527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_588_inst_ack_1, ack => cp_elements(137)); -- 
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(142));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => binary_597_inst_req_0); -- 
    cp_elements(139) <= cp_elements(25);
    cpelement_group_140 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(141));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(140),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => type_cast_593_inst_req_0); -- 
    cp_elements(141) <= cp_elements(25);
    ack_1539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => cp_elements(142)); -- 
    ra_1544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_597_inst_ack_0, ack => cp_elements(143)); -- 
    cr_1545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => binary_597_inst_req_1); -- 
    ca_1546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_597_inst_ack_1, ack => cp_elements(144)); -- 
    cpelement_group_145 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(79) & cp_elements(144));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(145),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(146) <= cp_elements(1);
    cp_elements(147) <= false;
    cp_elements(148) <= cp_elements(147);
    cp_elements(149) <= cp_elements(1);
    branch_req_1554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => if_stmt_599_branch_req_0); -- 
    cp_elements(150) <= cp_elements(149);
    cp_elements(151) <= cp_elements(150);
    if_choice_transition_1559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_599_branch_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(150);
    else_choice_transition_1563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_599_branch_ack_0, ack => cp_elements(154)); -- 
    cra_1576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_607_call_ack_0, ack => cp_elements(155)); -- 
    ccr_1580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => call_stmt_607_call_req_1); -- 
    cca_1581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_607_call_ack_1, ack => cp_elements(156)); -- 
    cp_elements(157) <= cp_elements(154);
    cpelement_group_158 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(159) & cp_elements(160));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => type_cast_612_inst_req_0); -- 
    cp_elements(159) <= cp_elements(157);
    cp_elements(160) <= cp_elements(157);
    cp_elements(161) <= type_cast_612_inst_ack_0;
    cpelement_group_162 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(161) & cp_elements(178));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(162),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(163) <= cp_elements(161);
    base_resize_req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => ptr_deref_616_base_resize_req_0); -- 
    base_resize_ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_base_resize_ack_0, ack => cp_elements(164)); -- 
    sum_rename_req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => ptr_deref_616_root_address_inst_req_0); -- 
    cp_elements(165) <= ptr_deref_616_root_address_inst_ack_0;
    cp_elements(166) <= cp_elements(165);
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => ptr_deref_616_addr_0_req_0); -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_0_ack_0, ack => cp_elements(167)); -- 
    cr_1624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => ptr_deref_616_addr_0_req_1); -- 
    ca_1625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_0_ack_1, ack => cp_elements(168)); -- 
    cp_elements(169) <= cp_elements(165);
    rr_1629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => ptr_deref_616_addr_1_req_0); -- 
    ra_1630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_1_ack_0, ack => cp_elements(170)); -- 
    cr_1631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => ptr_deref_616_addr_1_req_1); -- 
    ca_1632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_1_ack_1, ack => cp_elements(171)); -- 
    cp_elements(172) <= cp_elements(165);
    rr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(172), ack => ptr_deref_616_addr_2_req_0); -- 
    ra_1637_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_2_ack_0, ack => cp_elements(173)); -- 
    cr_1638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => ptr_deref_616_addr_2_req_1); -- 
    ca_1639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_2_ack_1, ack => cp_elements(174)); -- 
    cp_elements(175) <= cp_elements(165);
    rr_1643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(175), ack => ptr_deref_616_addr_3_req_0); -- 
    ra_1644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_3_ack_0, ack => cp_elements(176)); -- 
    cr_1645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => ptr_deref_616_addr_3_req_1); -- 
    ca_1646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_addr_3_ack_1, ack => cp_elements(177)); -- 
    cpelement_group_178 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(168) & cp_elements(171) & cp_elements(174) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(178),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(179) <= cp_elements(162);
    rr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => ptr_deref_616_load_0_req_0); -- 
    ra_1657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_0_ack_0, ack => cp_elements(180)); -- 
    cp_elements(181) <= cp_elements(162);
    rr_1661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => ptr_deref_616_load_1_req_0); -- 
    ra_1662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_1_ack_0, ack => cp_elements(182)); -- 
    cp_elements(183) <= cp_elements(162);
    rr_1666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => ptr_deref_616_load_2_req_0); -- 
    ra_1667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_2_ack_0, ack => cp_elements(184)); -- 
    cp_elements(185) <= cp_elements(162);
    rr_1671_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => ptr_deref_616_load_3_req_0); -- 
    ra_1672_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_3_ack_0, ack => cp_elements(186)); -- 
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(180) & cp_elements(182) & cp_elements(184) & cp_elements(186));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(188) <= cp_elements(187);
    cr_1682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => ptr_deref_616_load_0_req_1); -- 
    ca_1683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_0_ack_1, ack => cp_elements(189)); -- 
    cp_elements(190) <= cp_elements(187);
    cr_1687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_616_load_1_req_1); -- 
    ca_1688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_1_ack_1, ack => cp_elements(191)); -- 
    cp_elements(192) <= cp_elements(187);
    cr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => ptr_deref_616_load_2_req_1); -- 
    ca_1693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_2_ack_1, ack => cp_elements(193)); -- 
    cp_elements(194) <= cp_elements(187);
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => ptr_deref_616_load_3_req_1); -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_616_load_3_ack_1, ack => cp_elements(195)); -- 
    cpelement_group_196 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(189) & cp_elements(191) & cp_elements(193) & cp_elements(195));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(196),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_1699_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => ptr_deref_616_gather_scatter_req_0); -- 
    cp_elements(197) <= ptr_deref_616_gather_scatter_ack_0;
    cpelement_group_198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(199) & cp_elements(200));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1709_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => binary_622_inst_req_0); -- 
    cp_elements(199) <= cp_elements(157);
    cp_elements(200) <= cp_elements(197);
    ra_1710_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_622_inst_ack_0, ack => cp_elements(201)); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => binary_622_inst_req_1); -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_622_inst_ack_1, ack => cp_elements(202)); -- 
    cpelement_group_203 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(202) & cp_elements(204));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(203),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => binary_628_inst_req_0); -- 
    cp_elements(204) <= cp_elements(157);
    ra_1722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_628_inst_ack_0, ack => cp_elements(205)); -- 
    cr_1723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => binary_628_inst_req_1); -- 
    ca_1724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_628_inst_ack_1, ack => cp_elements(206)); -- 
    cpelement_group_207 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(208) & cp_elements(209));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(207),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => binary_634_inst_req_0); -- 
    cp_elements(208) <= cp_elements(157);
    cp_elements(209) <= cp_elements(197);
    ra_1734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_634_inst_ack_0, ack => cp_elements(210)); -- 
    cr_1735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => binary_634_inst_req_1); -- 
    ca_1736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_634_inst_ack_1, ack => cp_elements(211)); -- 
    cpelement_group_212 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(213));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => type_cast_638_inst_req_0); -- 
    cp_elements(213) <= cp_elements(157);
    ack_1746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_638_inst_ack_0, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(206) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= cp_elements(3);
    cp_elements(217) <= false;
    cp_elements(218) <= cp_elements(217);
    cp_elements(219) <= cp_elements(3);
    branch_req_1754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => if_stmt_640_branch_req_0); -- 
    cp_elements(220) <= cp_elements(219);
    cp_elements(221) <= cp_elements(220);
    if_choice_transition_1759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_640_branch_ack_1, ack => cp_elements(222)); -- 
    cp_elements(223) <= cp_elements(220);
    else_choice_transition_1763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_640_branch_ack_0, ack => cp_elements(224)); -- 
    cra_1776_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_648_call_ack_0, ack => cp_elements(225)); -- 
    ccr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => call_stmt_648_call_req_1); -- 
    cca_1781_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_648_call_ack_1, ack => cp_elements(226)); -- 
    cp_elements(227) <= cp_elements(222);
    cpelement_group_228 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(229) & cp_elements(230));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(228),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => binary_655_inst_req_0); -- 
    cp_elements(229) <= cp_elements(227);
    cp_elements(230) <= cp_elements(227);
    ra_1796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_655_inst_ack_0, ack => cp_elements(231)); -- 
    cr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => binary_655_inst_req_1); -- 
    ca_1798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_655_inst_ack_1, ack => cp_elements(232)); -- 
    cpelement_group_233 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(232) & cp_elements(234));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(233),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => binary_661_inst_req_0); -- 
    cp_elements(234) <= cp_elements(227);
    ra_1808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_661_inst_ack_0, ack => cp_elements(235)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => binary_661_inst_req_1); -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_661_inst_ack_1, ack => cp_elements(236)); -- 
    cpelement_group_237 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(236) & cp_elements(238));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(237),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => binary_667_inst_req_0); -- 
    cp_elements(238) <= cp_elements(227);
    ra_1820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_667_inst_ack_0, ack => cp_elements(239)); -- 
    cr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => binary_667_inst_req_1); -- 
    ca_1822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_667_inst_ack_1, ack => cp_elements(240)); -- 
    cp_elements(241) <= cp_elements(240);
    cp_elements(242) <= false;
    cp_elements(243) <= cp_elements(242);
    cp_elements(244) <= cp_elements(240);
    branch_req_1830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => if_stmt_669_branch_req_0); -- 
    cp_elements(245) <= cp_elements(244);
    cp_elements(246) <= cp_elements(245);
    if_choice_transition_1835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_669_branch_ack_1, ack => cp_elements(247)); -- 
    cp_elements(248) <= cp_elements(245);
    else_choice_transition_1839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_669_branch_ack_0, ack => cp_elements(249)); -- 
    crr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => call_stmt_682_call_req_0); -- 
    cra_1852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_677_call_ack_0, ack => cp_elements(250)); -- 
    ccr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => call_stmt_677_call_req_1); -- 
    cca_1857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_677_call_ack_1, ack => cp_elements(251)); -- 
    cra_1870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_682_call_ack_0, ack => cp_elements(252)); -- 
    ccr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => call_stmt_682_call_req_1); -- 
    cca_1875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_682_call_ack_1, ack => cp_elements(253)); -- 
    cp_elements(254) <= cp_elements(253);
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(256) & cp_elements(257));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => type_cast_685_inst_req_0); -- 
    cp_elements(256) <= cp_elements(254);
    cp_elements(257) <= cp_elements(254);
    cp_elements(258) <= type_cast_685_inst_ack_0;
    cpelement_group_259 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(260) & cp_elements(261) & cp_elements(262));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => binary_690_inst_req_0); -- 
    cp_elements(260) <= cp_elements(254);
    cp_elements(261) <= cp_elements(258);
    cp_elements(262) <= cp_elements(254);
    ra_1901_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_690_inst_ack_0, ack => cp_elements(263)); -- 
    cr_1902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => binary_690_inst_req_1); -- 
    ca_1903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_690_inst_ack_1, ack => cp_elements(264)); -- 
    cpelement_group_265 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(266) & cp_elements(267) & cp_elements(268));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(265),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => binary_695_inst_req_0); -- 
    cp_elements(266) <= cp_elements(254);
    cp_elements(267) <= cp_elements(258);
    cp_elements(268) <= cp_elements(254);
    ra_1914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_695_inst_ack_0, ack => cp_elements(269)); -- 
    cr_1915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => binary_695_inst_req_1); -- 
    ca_1916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_695_inst_ack_1, ack => cp_elements(270)); -- 
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(264) & cp_elements(270) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => binary_700_inst_req_0); -- 
    cp_elements(272) <= cp_elements(254);
    ra_1927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_700_inst_ack_0, ack => cp_elements(273)); -- 
    cr_1928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => binary_700_inst_req_1); -- 
    ca_1929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_700_inst_ack_1, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(274);
    cp_elements(276) <= false;
    cp_elements(277) <= cp_elements(276);
    cp_elements(278) <= cp_elements(274);
    branch_req_1937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(278), ack => if_stmt_702_branch_req_0); -- 
    cp_elements(279) <= cp_elements(278);
    cp_elements(280) <= cp_elements(279);
    if_choice_transition_1942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_702_branch_ack_1, ack => cp_elements(281)); -- 
    cp_elements(282) <= cp_elements(279);
    else_choice_transition_1946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_702_branch_ack_0, ack => cp_elements(283)); -- 
    cra_1959_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_0, ack => cp_elements(284)); -- 
    ccr_1963_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => call_stmt_710_call_req_1); -- 
    cca_1964_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(283);
    cpelement_group_287 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(288) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(287),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(287), ack => binary_717_inst_req_0); -- 
    cp_elements(288) <= cp_elements(286);
    cp_elements(289) <= cp_elements(286);
    ra_1979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_717_inst_ack_0, ack => cp_elements(290)); -- 
    cr_1980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => binary_717_inst_req_1); -- 
    ca_1981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_717_inst_ack_1, ack => cp_elements(291)); -- 
    cp_elements(292) <= cp_elements(291);
    cp_elements(293) <= false;
    cp_elements(294) <= cp_elements(293);
    cp_elements(295) <= cp_elements(291);
    branch_req_1989_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => if_stmt_719_branch_req_0); -- 
    cp_elements(296) <= cp_elements(295);
    cp_elements(297) <= cp_elements(296);
    if_choice_transition_1994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_719_branch_ack_1, ack => cp_elements(298)); -- 
    cp_elements(299) <= cp_elements(296);
    else_choice_transition_1998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_719_branch_ack_0, ack => cp_elements(300)); -- 
    cp_elements(301) <= cp_elements(7);
    cpelement_group_302 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(303) & cp_elements(304));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(302),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(302), ack => binary_730_inst_req_0); -- 
    cp_elements(303) <= cp_elements(301);
    cp_elements(304) <= cp_elements(301);
    ra_2013_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_730_inst_ack_0, ack => cp_elements(305)); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(305), ack => binary_730_inst_req_1); -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_730_inst_ack_1, ack => cp_elements(306)); -- 
    cp_elements(307) <= cp_elements(8);
    cpelement_group_308 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(309) & cp_elements(310));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => binary_753_inst_req_0); -- 
    cp_elements(309) <= cp_elements(307);
    cp_elements(310) <= cp_elements(307);
    ra_2028_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_753_inst_ack_0, ack => cp_elements(311)); -- 
    cr_2029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(311), ack => binary_753_inst_req_1); -- 
    ca_2030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_753_inst_ack_1, ack => cp_elements(312)); -- 
    cpelement_group_313 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(312) & cp_elements(314) & cp_elements(315));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(313),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(313), ack => binary_758_inst_req_0); -- 
    cp_elements(314) <= cp_elements(307);
    cp_elements(315) <= cp_elements(307);
    ra_2041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_758_inst_ack_0, ack => cp_elements(316)); -- 
    cr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => binary_758_inst_req_1); -- 
    ca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_758_inst_ack_1, ack => cp_elements(317)); -- 
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(319) & cp_elements(320));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => binary_764_inst_req_0); -- 
    cp_elements(319) <= cp_elements(307);
    cp_elements(320) <= cp_elements(307);
    ra_2053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_764_inst_ack_0, ack => cp_elements(321)); -- 
    cr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => binary_764_inst_req_1); -- 
    ca_2055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_764_inst_ack_1, ack => cp_elements(322)); -- 
    cpelement_group_323 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(322) & cp_elements(324));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(323),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(323), ack => binary_770_inst_req_0); -- 
    cp_elements(324) <= cp_elements(307);
    ra_2065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_770_inst_ack_0, ack => cp_elements(325)); -- 
    cr_2066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => binary_770_inst_req_1); -- 
    ca_2067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_770_inst_ack_1, ack => cp_elements(326)); -- 
    index_resize_req_2082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(326), ack => array_obj_ref_774_index_0_resize_req_0); -- 
    cp_elements(327) <= cp_elements(307);
    cpelement_group_328 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(327) & cp_elements(336));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => array_obj_ref_774_final_reg_req_0); -- 
    cp_elements(329) <= cp_elements(307);
    base_resize_req_2098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => array_obj_ref_774_base_resize_req_0); -- 
    index_resize_ack_2083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_index_0_resize_ack_0, ack => cp_elements(330)); -- 
    scale_rename_req_2087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => array_obj_ref_774_index_0_rename_req_0); -- 
    scale_rename_ack_2088_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_index_0_rename_ack_0, ack => cp_elements(331)); -- 
    final_index_req_2092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => array_obj_ref_774_offset_inst_req_0); -- 
    final_index_ack_2093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_offset_inst_ack_0, ack => cp_elements(332)); -- 
    base_resize_ack_2099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_base_resize_ack_0, ack => cp_elements(333)); -- 
    cpelement_group_334 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(332) & cp_elements(333));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(334),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(334), ack => array_obj_ref_774_root_address_inst_req_0); -- 
    plus_base_ra_2105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_root_address_inst_ack_0, ack => cp_elements(335)); -- 
    plus_base_cr_2106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => array_obj_ref_774_root_address_inst_req_1); -- 
    plus_base_ca_2107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_root_address_inst_ack_1, ack => cp_elements(336)); -- 
    final_reg_ack_2112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_774_final_reg_ack_0, ack => cp_elements(337)); -- 
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(337) & cp_elements(339));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => type_cast_779_inst_req_0); -- 
    cp_elements(339) <= cp_elements(307);
    cp_elements(340) <= type_cast_779_inst_ack_0;
    cpelement_group_341 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(340) & cp_elements(351));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(341),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(342) <= cp_elements(340);
    base_resize_req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(342), ack => ptr_deref_783_base_resize_req_0); -- 
    base_resize_ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_base_resize_ack_0, ack => cp_elements(343)); -- 
    sum_rename_req_2140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(343), ack => ptr_deref_783_root_address_inst_req_0); -- 
    cp_elements(344) <= ptr_deref_783_root_address_inst_ack_0;
    cp_elements(345) <= cp_elements(344);
    rr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => ptr_deref_783_addr_0_req_0); -- 
    ra_2149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_addr_0_ack_0, ack => cp_elements(346)); -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(346), ack => ptr_deref_783_addr_0_req_1); -- 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_addr_0_ack_1, ack => cp_elements(347)); -- 
    cp_elements(348) <= cp_elements(344);
    rr_2155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => ptr_deref_783_addr_1_req_0); -- 
    ra_2156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_addr_1_ack_0, ack => cp_elements(349)); -- 
    cr_2157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(349), ack => ptr_deref_783_addr_1_req_1); -- 
    ca_2158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_addr_1_ack_1, ack => cp_elements(350)); -- 
    cpelement_group_351 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(350));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(351),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(352) <= cp_elements(341);
    rr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(352), ack => ptr_deref_783_load_0_req_0); -- 
    ra_2169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_load_0_ack_0, ack => cp_elements(353)); -- 
    cp_elements(354) <= cp_elements(341);
    rr_2173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(354), ack => ptr_deref_783_load_1_req_0); -- 
    ra_2174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_load_1_ack_0, ack => cp_elements(355)); -- 
    cpelement_group_356 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(353) & cp_elements(355));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(356),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(357) <= cp_elements(356);
    cr_2184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => ptr_deref_783_load_0_req_1); -- 
    ca_2185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_load_0_ack_1, ack => cp_elements(358)); -- 
    cp_elements(359) <= cp_elements(356);
    cr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(359), ack => ptr_deref_783_load_1_req_1); -- 
    ca_2190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_load_1_ack_1, ack => cp_elements(360)); -- 
    cpelement_group_361 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(358) & cp_elements(360));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(361),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(361), ack => ptr_deref_783_gather_scatter_req_0); -- 
    merge_ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_783_gather_scatter_ack_0, ack => cp_elements(362)); -- 
    cpelement_group_363 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(362) & cp_elements(364));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(363),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(363), ack => type_cast_787_inst_req_0); -- 
    cp_elements(364) <= cp_elements(307);
    ack_2202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_0, ack => cp_elements(365)); -- 
    cpelement_group_366 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(365) & cp_elements(367) & cp_elements(368));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(366),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(366), ack => binary_792_inst_req_0); -- 
    cp_elements(367) <= cp_elements(307);
    cp_elements(368) <= cp_elements(307);
    ra_2213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_792_inst_ack_0, ack => cp_elements(369)); -- 
    cr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(369), ack => binary_792_inst_req_1); -- 
    ca_2215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_792_inst_ack_1, ack => cp_elements(370)); -- 
    cpelement_group_371 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(372) & cp_elements(375));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => binary_800_inst_req_0); -- 
    cp_elements(372) <= cp_elements(307);
    cpelement_group_373 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(317) & cp_elements(374));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(373),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(373), ack => type_cast_796_inst_req_0); -- 
    cp_elements(374) <= cp_elements(307);
    ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_0, ack => cp_elements(375)); -- 
    ra_2232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_800_inst_ack_0, ack => cp_elements(376)); -- 
    cr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(376), ack => binary_800_inst_req_1); -- 
    ca_2234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_800_inst_ack_1, ack => cp_elements(377)); -- 
    cpelement_group_378 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(379) & cp_elements(380));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(378),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(378), ack => binary_806_inst_req_0); -- 
    cp_elements(379) <= cp_elements(307);
    cp_elements(380) <= cp_elements(307);
    ra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_806_inst_ack_0, ack => cp_elements(381)); -- 
    cr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => binary_806_inst_req_1); -- 
    ca_2246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_806_inst_ack_1, ack => cp_elements(382)); -- 
    cpelement_group_383 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(370) & cp_elements(377) & cp_elements(382));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(383),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(384) <= cp_elements(9);
    cp_elements(385) <= false;
    cp_elements(386) <= cp_elements(385);
    cp_elements(387) <= cp_elements(9);
    branch_req_2254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(387), ack => if_stmt_808_branch_req_0); -- 
    cp_elements(388) <= cp_elements(387);
    cp_elements(389) <= cp_elements(388);
    if_choice_transition_2259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_808_branch_ack_1, ack => cp_elements(390)); -- 
    cp_elements(391) <= cp_elements(388);
    else_choice_transition_2263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_808_branch_ack_0, ack => cp_elements(392)); -- 
    cp_elements(393) <= cp_elements(10);
    cpelement_group_394 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(395) & cp_elements(396));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(394),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(394), ack => binary_819_inst_req_0); -- 
    cp_elements(395) <= cp_elements(393);
    cp_elements(396) <= cp_elements(393);
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_819_inst_ack_0, ack => cp_elements(397)); -- 
    cr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(397), ack => binary_819_inst_req_1); -- 
    ca_2280_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_819_inst_ack_1, ack => cp_elements(398)); -- 
    index_resize_req_2295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(398), ack => array_obj_ref_823_index_0_resize_req_0); -- 
    cp_elements(399) <= cp_elements(393);
    cpelement_group_400 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(399) & cp_elements(408));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(400),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(400), ack => array_obj_ref_823_final_reg_req_0); -- 
    cp_elements(401) <= cp_elements(393);
    base_resize_req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(401), ack => array_obj_ref_823_base_resize_req_0); -- 
    index_resize_ack_2296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_index_0_resize_ack_0, ack => cp_elements(402)); -- 
    scale_rename_req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => array_obj_ref_823_index_0_rename_req_0); -- 
    scale_rename_ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_index_0_rename_ack_0, ack => cp_elements(403)); -- 
    final_index_req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(403), ack => array_obj_ref_823_offset_inst_req_0); -- 
    final_index_ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_offset_inst_ack_0, ack => cp_elements(404)); -- 
    base_resize_ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_base_resize_ack_0, ack => cp_elements(405)); -- 
    cpelement_group_406 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(404) & cp_elements(405));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(406),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => array_obj_ref_823_root_address_inst_req_0); -- 
    plus_base_ra_2318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_root_address_inst_ack_0, ack => cp_elements(407)); -- 
    plus_base_cr_2319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(407), ack => array_obj_ref_823_root_address_inst_req_1); -- 
    plus_base_ca_2320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_root_address_inst_ack_1, ack => cp_elements(408)); -- 
    final_reg_ack_2325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_823_final_reg_ack_0, ack => cp_elements(409)); -- 
    cp_elements(410) <= cp_elements(11);
    cpelement_group_411 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(412) & cp_elements(413));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(411),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => binary_851_inst_req_0); -- 
    cp_elements(412) <= cp_elements(410);
    cp_elements(413) <= cp_elements(410);
    ra_2338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_851_inst_ack_0, ack => cp_elements(414)); -- 
    cr_2339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(414), ack => binary_851_inst_req_1); -- 
    ca_2340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_851_inst_ack_1, ack => cp_elements(415)); -- 
    cp_elements(416) <= cp_elements(415);
    cp_elements(417) <= false;
    cp_elements(418) <= cp_elements(417);
    cp_elements(419) <= cp_elements(415);
    branch_req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(419), ack => if_stmt_853_branch_req_0); -- 
    cp_elements(420) <= cp_elements(419);
    cp_elements(421) <= cp_elements(420);
    if_choice_transition_2353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_853_branch_ack_1, ack => cp_elements(422)); -- 
    cp_elements(423) <= cp_elements(420);
    cp_elements(424) <= if_stmt_853_branch_ack_0;
    cp_elements(425) <= cp_elements(12);
    cpelement_group_426 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(427) & cp_elements(431));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(426),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(426), ack => ptr_deref_862_load_0_req_0); -- 
    cp_elements(427) <= cp_elements(425);
    cp_elements(428) <= cp_elements(427);
    base_resize_req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(428), ack => ptr_deref_862_base_resize_req_0); -- 
    base_resize_ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_862_base_resize_ack_0, ack => cp_elements(429)); -- 
    sum_rename_req_2380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(429), ack => ptr_deref_862_root_address_inst_req_0); -- 
    sum_rename_ack_2381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_862_root_address_inst_ack_0, ack => cp_elements(430)); -- 
    root_rename_req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(430), ack => ptr_deref_862_addr_0_req_0); -- 
    root_rename_ack_2386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_862_addr_0_ack_0, ack => cp_elements(431)); -- 
    ra_2397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_862_load_0_ack_0, ack => cp_elements(432)); -- 
    cr_2407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(432), ack => ptr_deref_862_load_0_req_1); -- 
    ca_2408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_862_load_0_ack_1, ack => cp_elements(433)); -- 
    merge_req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(433), ack => ptr_deref_862_gather_scatter_req_0); -- 
    merge_ack_2410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_862_gather_scatter_ack_0, ack => cp_elements(434)); -- 
    cpelement_group_435 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(434) & cp_elements(436));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(435),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => type_cast_866_inst_req_0); -- 
    cp_elements(436) <= cp_elements(425);
    ack_2420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_866_inst_ack_0, ack => cp_elements(437)); -- 
    cpelement_group_438 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(437) & cp_elements(439) & cp_elements(440));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(438),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => binary_871_inst_req_0); -- 
    cp_elements(439) <= cp_elements(425);
    cp_elements(440) <= cp_elements(425);
    ra_2431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_871_inst_ack_0, ack => cp_elements(441)); -- 
    cr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(441), ack => binary_871_inst_req_1); -- 
    cp_elements(442) <= binary_871_inst_ack_1;
    cp_elements(443) <= cp_elements(964);
    cpelement_group_444 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(445) & cp_elements(446));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(444),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => binary_886_inst_req_0); -- 
    cp_elements(445) <= cp_elements(443);
    cp_elements(446) <= cp_elements(443);
    ra_2446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_886_inst_ack_0, ack => cp_elements(447)); -- 
    cr_2447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(447), ack => binary_886_inst_req_1); -- 
    ca_2448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_886_inst_ack_1, ack => cp_elements(448)); -- 
    cpelement_group_449 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(450) & cp_elements(451));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(449),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => binary_892_inst_req_0); -- 
    cp_elements(450) <= cp_elements(443);
    cp_elements(451) <= cp_elements(443);
    ra_2458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_892_inst_ack_0, ack => cp_elements(452)); -- 
    cr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(452), ack => binary_892_inst_req_1); -- 
    ca_2460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_892_inst_ack_1, ack => cp_elements(453)); -- 
    cpelement_group_454 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(448) & cp_elements(453) & cp_elements(455));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(454),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(454), ack => binary_897_inst_req_0); -- 
    cp_elements(455) <= cp_elements(443);
    ra_2471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_897_inst_ack_0, ack => cp_elements(456)); -- 
    cr_2472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(456), ack => binary_897_inst_req_1); -- 
    cp_elements(457) <= binary_897_inst_ack_1;
    cpelement_group_458 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(459) & cp_elements(460));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(458),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => binary_903_inst_req_0); -- 
    cp_elements(459) <= cp_elements(443);
    cp_elements(460) <= cp_elements(457);
    ra_2483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_903_inst_ack_0, ack => cp_elements(461)); -- 
    cr_2484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => binary_903_inst_req_1); -- 
    ca_2485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_903_inst_ack_1, ack => cp_elements(462)); -- 
    cpelement_group_463 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(462) & cp_elements(464) & cp_elements(465));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(463),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(463), ack => binary_908_inst_req_0); -- 
    cp_elements(464) <= cp_elements(443);
    cp_elements(465) <= cp_elements(457);
    ra_2496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_908_inst_ack_0, ack => cp_elements(466)); -- 
    cr_2497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(466), ack => binary_908_inst_req_1); -- 
    ca_2498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_908_inst_ack_1, ack => cp_elements(467)); -- 
    cpelement_group_468 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(467) & cp_elements(469));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(468),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2507_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(468), ack => type_cast_912_inst_req_0); -- 
    cp_elements(469) <= cp_elements(443);
    ack_2508_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_912_inst_ack_0, ack => cp_elements(470)); -- 
    cpelement_group_471 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(470) & cp_elements(472));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(471),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(471), ack => binary_918_inst_req_0); -- 
    cp_elements(472) <= cp_elements(443);
    ra_2518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_918_inst_ack_0, ack => cp_elements(473)); -- 
    cr_2519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(473), ack => binary_918_inst_req_1); -- 
    ca_2520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_918_inst_ack_1, ack => cp_elements(474)); -- 
    cp_elements(475) <= cp_elements(474);
    cp_elements(476) <= false;
    cp_elements(477) <= cp_elements(476);
    cp_elements(478) <= cp_elements(474);
    branch_req_2528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(478), ack => if_stmt_920_branch_req_0); -- 
    cp_elements(479) <= cp_elements(478);
    cp_elements(480) <= cp_elements(479);
    if_choice_transition_2533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_920_branch_ack_1, ack => cp_elements(481)); -- 
    cp_elements(482) <= cp_elements(479);
    else_choice_transition_2537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_920_branch_ack_0, ack => cp_elements(483)); -- 
    cra_2550_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_928_call_ack_0, ack => cp_elements(484)); -- 
    ccr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(484), ack => call_stmt_928_call_req_1); -- 
    cca_2555_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_928_call_ack_1, ack => cp_elements(485)); -- 
    cp_elements(486) <= cp_elements(481);
    cp_elements(487) <= cp_elements(486);
    cpelement_group_488 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(487) & cp_elements(492));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(488),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2584_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(488), ack => array_obj_ref_936_final_reg_req_0); -- 
    cp_elements(489) <= cp_elements(486);
    base_resize_req_2571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(489), ack => array_obj_ref_936_base_resize_req_0); -- 
    base_resize_ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_936_base_resize_ack_0, ack => cp_elements(490)); -- 
    plus_base_rr_2577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => array_obj_ref_936_root_address_inst_req_0); -- 
    plus_base_ra_2578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_936_root_address_inst_ack_0, ack => cp_elements(491)); -- 
    plus_base_cr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(491), ack => array_obj_ref_936_root_address_inst_req_1); -- 
    plus_base_ca_2580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_936_root_address_inst_ack_1, ack => cp_elements(492)); -- 
    cp_elements(493) <= array_obj_ref_936_final_reg_ack_0;
    cp_elements(494) <= cp_elements(486);
    cpelement_group_495 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(493) & cp_elements(494) & cp_elements(511));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(495),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(495), ack => ptr_deref_939_gather_scatter_req_0); -- 
    cp_elements(496) <= cp_elements(493);
    base_resize_req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => ptr_deref_939_base_resize_req_0); -- 
    base_resize_ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_base_resize_ack_0, ack => cp_elements(497)); -- 
    sum_rename_req_2604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(497), ack => ptr_deref_939_root_address_inst_req_0); -- 
    cp_elements(498) <= ptr_deref_939_root_address_inst_ack_0;
    cp_elements(499) <= cp_elements(498);
    rr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => ptr_deref_939_addr_0_req_0); -- 
    ra_2613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_0_ack_0, ack => cp_elements(500)); -- 
    cr_2614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => ptr_deref_939_addr_0_req_1); -- 
    ca_2615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_0_ack_1, ack => cp_elements(501)); -- 
    cp_elements(502) <= cp_elements(498);
    rr_2619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(502), ack => ptr_deref_939_addr_1_req_0); -- 
    ra_2620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_1_ack_0, ack => cp_elements(503)); -- 
    cr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => ptr_deref_939_addr_1_req_1); -- 
    ca_2622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_1_ack_1, ack => cp_elements(504)); -- 
    cp_elements(505) <= cp_elements(498);
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(505), ack => ptr_deref_939_addr_2_req_0); -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_2_ack_0, ack => cp_elements(506)); -- 
    cr_2628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => ptr_deref_939_addr_2_req_1); -- 
    ca_2629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_2_ack_1, ack => cp_elements(507)); -- 
    cp_elements(508) <= cp_elements(498);
    rr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(508), ack => ptr_deref_939_addr_3_req_0); -- 
    ra_2634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_3_ack_0, ack => cp_elements(509)); -- 
    cr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => ptr_deref_939_addr_3_req_1); -- 
    ca_2636_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_addr_3_ack_1, ack => cp_elements(510)); -- 
    cpelement_group_511 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(501) & cp_elements(504) & cp_elements(507) & cp_elements(510));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(511),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(512) <= ptr_deref_939_gather_scatter_ack_0;
    cp_elements(513) <= cp_elements(512);
    rr_2648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(513), ack => ptr_deref_939_store_0_req_0); -- 
    ra_2649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_0_ack_0, ack => cp_elements(514)); -- 
    cp_elements(515) <= cp_elements(512);
    rr_2653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => ptr_deref_939_store_1_req_0); -- 
    ra_2654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_1_ack_0, ack => cp_elements(516)); -- 
    cp_elements(517) <= cp_elements(512);
    rr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => ptr_deref_939_store_2_req_0); -- 
    ra_2659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_2_ack_0, ack => cp_elements(518)); -- 
    cp_elements(519) <= cp_elements(512);
    rr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => ptr_deref_939_store_3_req_0); -- 
    ra_2664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_3_ack_0, ack => cp_elements(520)); -- 
    cpelement_group_521 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(514) & cp_elements(516) & cp_elements(518) & cp_elements(520));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(521),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(522) <= cp_elements(521);
    cp_elements(523) <= cp_elements(522);
    cr_2674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(523), ack => ptr_deref_939_store_0_req_1); -- 
    ca_2675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_0_ack_1, ack => cp_elements(524)); -- 
    cp_elements(525) <= cp_elements(522);
    cr_2679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(525), ack => ptr_deref_939_store_1_req_1); -- 
    ca_2680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_1_ack_1, ack => cp_elements(526)); -- 
    cp_elements(527) <= cp_elements(522);
    cr_2684_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(527), ack => ptr_deref_939_store_2_req_1); -- 
    ca_2685_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_2_ack_1, ack => cp_elements(528)); -- 
    cp_elements(529) <= cp_elements(522);
    cr_2689_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(529), ack => ptr_deref_939_store_3_req_1); -- 
    ca_2690_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_939_store_3_ack_1, ack => cp_elements(530)); -- 
    cpelement_group_531 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(524) & cp_elements(526) & cp_elements(528) & cp_elements(530));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(531),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_532 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(533) & cp_elements(534));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(532),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2699_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(532), ack => binary_946_inst_req_0); -- 
    cp_elements(533) <= cp_elements(486);
    cp_elements(534) <= cp_elements(486);
    ra_2700_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_946_inst_ack_0, ack => cp_elements(535)); -- 
    cr_2701_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(535), ack => binary_946_inst_req_1); -- 
    ca_2702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_946_inst_ack_1, ack => cp_elements(536)); -- 
    index_resize_req_2717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(536), ack => array_obj_ref_950_index_0_resize_req_0); -- 
    cp_elements(537) <= cp_elements(486);
    cpelement_group_538 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(537) & cp_elements(546));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(538),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => array_obj_ref_950_final_reg_req_0); -- 
    cp_elements(539) <= cp_elements(486);
    base_resize_req_2733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(539), ack => array_obj_ref_950_base_resize_req_0); -- 
    index_resize_ack_2718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_0_resize_ack_0, ack => cp_elements(540)); -- 
    scale_rename_req_2722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(540), ack => array_obj_ref_950_index_0_rename_req_0); -- 
    scale_rename_ack_2723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_0_rename_ack_0, ack => cp_elements(541)); -- 
    final_index_req_2727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => array_obj_ref_950_offset_inst_req_0); -- 
    final_index_ack_2728_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_offset_inst_ack_0, ack => cp_elements(542)); -- 
    base_resize_ack_2734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_base_resize_ack_0, ack => cp_elements(543)); -- 
    cpelement_group_544 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(542) & cp_elements(543));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(544),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(544), ack => array_obj_ref_950_root_address_inst_req_0); -- 
    plus_base_ra_2740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_root_address_inst_ack_0, ack => cp_elements(545)); -- 
    plus_base_cr_2741_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => array_obj_ref_950_root_address_inst_req_1); -- 
    plus_base_ca_2742_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_root_address_inst_ack_1, ack => cp_elements(546)); -- 
    final_reg_ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_final_reg_ack_0, ack => cp_elements(547)); -- 
    cp_elements(548) <= cp_elements(486);
    cpelement_group_549 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(548) & cp_elements(553));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(549),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(549), ack => array_obj_ref_957_final_reg_req_0); -- 
    cp_elements(550) <= cp_elements(486);
    base_resize_req_2758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => array_obj_ref_957_base_resize_req_0); -- 
    base_resize_ack_2759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_957_base_resize_ack_0, ack => cp_elements(551)); -- 
    plus_base_rr_2764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(551), ack => array_obj_ref_957_root_address_inst_req_0); -- 
    plus_base_ra_2765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_957_root_address_inst_ack_0, ack => cp_elements(552)); -- 
    plus_base_cr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => array_obj_ref_957_root_address_inst_req_1); -- 
    plus_base_ca_2767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_957_root_address_inst_ack_1, ack => cp_elements(553)); -- 
    cp_elements(554) <= array_obj_ref_957_final_reg_ack_0;
    cpelement_group_555 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(521) & cp_elements(547) & cp_elements(554) & cp_elements(571));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(555),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(555), ack => ptr_deref_960_gather_scatter_req_0); -- 
    cp_elements(556) <= cp_elements(554);
    base_resize_req_2786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(556), ack => ptr_deref_960_base_resize_req_0); -- 
    base_resize_ack_2787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_base_resize_ack_0, ack => cp_elements(557)); -- 
    sum_rename_req_2791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(557), ack => ptr_deref_960_root_address_inst_req_0); -- 
    cp_elements(558) <= ptr_deref_960_root_address_inst_ack_0;
    cp_elements(559) <= cp_elements(558);
    rr_2799_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(559), ack => ptr_deref_960_addr_0_req_0); -- 
    ra_2800_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_0_ack_0, ack => cp_elements(560)); -- 
    cr_2801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(560), ack => ptr_deref_960_addr_0_req_1); -- 
    ca_2802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_0_ack_1, ack => cp_elements(561)); -- 
    cp_elements(562) <= cp_elements(558);
    rr_2806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(562), ack => ptr_deref_960_addr_1_req_0); -- 
    ra_2807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_1_ack_0, ack => cp_elements(563)); -- 
    cr_2808_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(563), ack => ptr_deref_960_addr_1_req_1); -- 
    ca_2809_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_1_ack_1, ack => cp_elements(564)); -- 
    cp_elements(565) <= cp_elements(558);
    rr_2813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(565), ack => ptr_deref_960_addr_2_req_0); -- 
    ra_2814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_2_ack_0, ack => cp_elements(566)); -- 
    cr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => ptr_deref_960_addr_2_req_1); -- 
    ca_2816_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_2_ack_1, ack => cp_elements(567)); -- 
    cp_elements(568) <= cp_elements(558);
    rr_2820_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(568), ack => ptr_deref_960_addr_3_req_0); -- 
    ra_2821_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_3_ack_0, ack => cp_elements(569)); -- 
    cr_2822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(569), ack => ptr_deref_960_addr_3_req_1); -- 
    ca_2823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_addr_3_ack_1, ack => cp_elements(570)); -- 
    cpelement_group_571 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(561) & cp_elements(564) & cp_elements(567) & cp_elements(570));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(571),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(572) <= ptr_deref_960_gather_scatter_ack_0;
    cp_elements(573) <= cp_elements(572);
    rr_2835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(573), ack => ptr_deref_960_store_0_req_0); -- 
    ra_2836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_0_ack_0, ack => cp_elements(574)); -- 
    cp_elements(575) <= cp_elements(572);
    rr_2840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => ptr_deref_960_store_1_req_0); -- 
    ra_2841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_1_ack_0, ack => cp_elements(576)); -- 
    cp_elements(577) <= cp_elements(572);
    rr_2845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(577), ack => ptr_deref_960_store_2_req_0); -- 
    ra_2846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_2_ack_0, ack => cp_elements(578)); -- 
    cp_elements(579) <= cp_elements(572);
    rr_2850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(579), ack => ptr_deref_960_store_3_req_0); -- 
    ra_2851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_3_ack_0, ack => cp_elements(580)); -- 
    cpelement_group_581 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(574) & cp_elements(576) & cp_elements(578) & cp_elements(580));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(581),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(582) <= cp_elements(581);
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(582), ack => ptr_deref_960_store_0_req_1); -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_0_ack_1, ack => cp_elements(583)); -- 
    cp_elements(584) <= cp_elements(581);
    cr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(584), ack => ptr_deref_960_store_1_req_1); -- 
    ca_2867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_1_ack_1, ack => cp_elements(585)); -- 
    cp_elements(586) <= cp_elements(581);
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => ptr_deref_960_store_2_req_1); -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_2_ack_1, ack => cp_elements(587)); -- 
    cp_elements(588) <= cp_elements(581);
    cr_2876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(588), ack => ptr_deref_960_store_3_req_1); -- 
    ca_2877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_3_ack_1, ack => cp_elements(589)); -- 
    cpelement_group_590 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(583) & cp_elements(585) & cp_elements(587) & cp_elements(589));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(590),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_591 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(592) & cp_elements(593) & cp_elements(594));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(591),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2887_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => binary_966_inst_req_0); -- 
    cp_elements(592) <= cp_elements(486);
    cp_elements(593) <= cp_elements(486);
    cp_elements(594) <= cp_elements(486);
    ra_2888_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_966_inst_ack_0, ack => cp_elements(595)); -- 
    cr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => binary_966_inst_req_1); -- 
    ca_2890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_966_inst_ack_1, ack => cp_elements(596)); -- 
    cpelement_group_597 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(531) & cp_elements(590) & cp_elements(596));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(597),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(598) <= cp_elements(14);
    cp_elements(599) <= false;
    cp_elements(600) <= cp_elements(599);
    cp_elements(601) <= cp_elements(14);
    branch_req_2898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(601), ack => if_stmt_968_branch_req_0); -- 
    cp_elements(602) <= cp_elements(601);
    cp_elements(603) <= cp_elements(602);
    if_choice_transition_2903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_968_branch_ack_1, ack => cp_elements(604)); -- 
    cp_elements(605) <= cp_elements(602);
    else_choice_transition_2907_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_968_branch_ack_0, ack => cp_elements(606)); -- 
    cp_elements(607) <= cp_elements(15);
    cpelement_group_608 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(609) & cp_elements(610) & cp_elements(611));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(608),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(608), ack => binary_978_inst_req_0); -- 
    cp_elements(609) <= cp_elements(607);
    cp_elements(610) <= cp_elements(607);
    cp_elements(611) <= cp_elements(607);
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_978_inst_ack_0, ack => cp_elements(612)); -- 
    cr_2924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(612), ack => binary_978_inst_req_1); -- 
    cp_elements(613) <= binary_978_inst_ack_1;
    cpelement_group_614 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(615) & cp_elements(616) & cp_elements(617));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(614),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(614), ack => binary_983_inst_req_0); -- 
    cp_elements(615) <= cp_elements(607);
    cp_elements(616) <= cp_elements(607);
    cp_elements(617) <= cp_elements(613);
    ra_2936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_983_inst_ack_0, ack => cp_elements(618)); -- 
    cr_2937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(618), ack => binary_983_inst_req_1); -- 
    ca_2938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_983_inst_ack_1, ack => cp_elements(619)); -- 
    cp_elements(620) <= cp_elements(607);
    cpelement_group_621 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(619) & cp_elements(620) & cp_elements(622) & cp_elements(623));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(621), ack => ternary_989_inst_req_0); -- 
    cp_elements(622) <= cp_elements(607);
    cp_elements(623) <= cp_elements(613);
    ack_2950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ternary_989_inst_ack_0, ack => cp_elements(624)); -- 
    cpelement_group_625 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(624) & cp_elements(626));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(625),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(625), ack => binary_995_inst_req_0); -- 
    cp_elements(626) <= cp_elements(607);
    ra_2960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_995_inst_ack_0, ack => cp_elements(627)); -- 
    cr_2961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(627), ack => binary_995_inst_req_1); -- 
    ca_2962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_995_inst_ack_1, ack => cp_elements(628)); -- 
    index_resize_req_2977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(628), ack => array_obj_ref_999_index_0_resize_req_0); -- 
    cp_elements(629) <= cp_elements(607);
    cpelement_group_630 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(629) & cp_elements(638));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(630),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => array_obj_ref_999_final_reg_req_0); -- 
    cp_elements(631) <= cp_elements(607);
    base_resize_req_2993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(631), ack => array_obj_ref_999_base_resize_req_0); -- 
    index_resize_ack_2978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_index_0_resize_ack_0, ack => cp_elements(632)); -- 
    scale_rename_req_2982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(632), ack => array_obj_ref_999_index_0_rename_req_0); -- 
    scale_rename_ack_2983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_index_0_rename_ack_0, ack => cp_elements(633)); -- 
    final_index_req_2987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(633), ack => array_obj_ref_999_offset_inst_req_0); -- 
    final_index_ack_2988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_offset_inst_ack_0, ack => cp_elements(634)); -- 
    base_resize_ack_2994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_base_resize_ack_0, ack => cp_elements(635)); -- 
    cpelement_group_636 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(634) & cp_elements(635));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(636),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => array_obj_ref_999_root_address_inst_req_0); -- 
    plus_base_ra_3000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_root_address_inst_ack_0, ack => cp_elements(637)); -- 
    plus_base_cr_3001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(637), ack => array_obj_ref_999_root_address_inst_req_1); -- 
    plus_base_ca_3002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_root_address_inst_ack_1, ack => cp_elements(638)); -- 
    final_reg_ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_999_final_reg_ack_0, ack => cp_elements(639)); -- 
    cpelement_group_640 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(639) & cp_elements(641) & cp_elements(657));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(640),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => ptr_deref_1002_gather_scatter_req_0); -- 
    cp_elements(641) <= cp_elements(607);
    cp_elements(642) <= cp_elements(641);
    base_resize_req_3021_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(642), ack => ptr_deref_1002_base_resize_req_0); -- 
    base_resize_ack_3022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_base_resize_ack_0, ack => cp_elements(643)); -- 
    sum_rename_req_3026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => ptr_deref_1002_root_address_inst_req_0); -- 
    cp_elements(644) <= ptr_deref_1002_root_address_inst_ack_0;
    cp_elements(645) <= cp_elements(644);
    rr_3034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(645), ack => ptr_deref_1002_addr_0_req_0); -- 
    ra_3035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_0_ack_0, ack => cp_elements(646)); -- 
    cr_3036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(646), ack => ptr_deref_1002_addr_0_req_1); -- 
    ca_3037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_0_ack_1, ack => cp_elements(647)); -- 
    cp_elements(648) <= cp_elements(644);
    rr_3041_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(648), ack => ptr_deref_1002_addr_1_req_0); -- 
    ra_3042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_1_ack_0, ack => cp_elements(649)); -- 
    cr_3043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(649), ack => ptr_deref_1002_addr_1_req_1); -- 
    ca_3044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_1_ack_1, ack => cp_elements(650)); -- 
    cp_elements(651) <= cp_elements(644);
    rr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(651), ack => ptr_deref_1002_addr_2_req_0); -- 
    ra_3049_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_2_ack_0, ack => cp_elements(652)); -- 
    cr_3050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => ptr_deref_1002_addr_2_req_1); -- 
    ca_3051_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_2_ack_1, ack => cp_elements(653)); -- 
    cp_elements(654) <= cp_elements(644);
    rr_3055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ptr_deref_1002_addr_3_req_0); -- 
    ra_3056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_3_ack_0, ack => cp_elements(655)); -- 
    cr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => ptr_deref_1002_addr_3_req_1); -- 
    ca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_addr_3_ack_1, ack => cp_elements(656)); -- 
    cpelement_group_657 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(647) & cp_elements(650) & cp_elements(653) & cp_elements(656));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(657),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(658) <= ptr_deref_1002_gather_scatter_ack_0;
    cp_elements(659) <= cp_elements(658);
    rr_3070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(659), ack => ptr_deref_1002_store_0_req_0); -- 
    ra_3071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_0_ack_0, ack => cp_elements(660)); -- 
    cp_elements(661) <= cp_elements(658);
    rr_3075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(661), ack => ptr_deref_1002_store_1_req_0); -- 
    ra_3076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_1_ack_0, ack => cp_elements(662)); -- 
    cp_elements(663) <= cp_elements(658);
    rr_3080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => ptr_deref_1002_store_2_req_0); -- 
    ra_3081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_2_ack_0, ack => cp_elements(664)); -- 
    cp_elements(665) <= cp_elements(658);
    rr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(665), ack => ptr_deref_1002_store_3_req_0); -- 
    ra_3086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_3_ack_0, ack => cp_elements(666)); -- 
    cpelement_group_667 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(660) & cp_elements(662) & cp_elements(664) & cp_elements(666));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(667),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(668) <= cp_elements(667);
    cp_elements(669) <= cp_elements(668);
    cr_3096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(669), ack => ptr_deref_1002_store_0_req_1); -- 
    ca_3097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_0_ack_1, ack => cp_elements(670)); -- 
    cp_elements(671) <= cp_elements(668);
    cr_3101_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(671), ack => ptr_deref_1002_store_1_req_1); -- 
    ca_3102_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_1_ack_1, ack => cp_elements(672)); -- 
    cp_elements(673) <= cp_elements(668);
    cr_3106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(673), ack => ptr_deref_1002_store_2_req_1); -- 
    ca_3107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_2_ack_1, ack => cp_elements(674)); -- 
    cp_elements(675) <= cp_elements(668);
    cr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(675), ack => ptr_deref_1002_store_3_req_1); -- 
    ca_3112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_3_ack_1, ack => cp_elements(676)); -- 
    cpelement_group_677 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(670) & cp_elements(672) & cp_elements(674) & cp_elements(676));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(677),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(678) <= cp_elements(607);
    cpelement_group_679 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(678) & cp_elements(683));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(679),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(679), ack => array_obj_ref_1008_final_reg_req_0); -- 
    cp_elements(680) <= cp_elements(607);
    base_resize_req_3123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(680), ack => array_obj_ref_1008_base_resize_req_0); -- 
    base_resize_ack_3124_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_base_resize_ack_0, ack => cp_elements(681)); -- 
    plus_base_rr_3129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(681), ack => array_obj_ref_1008_root_address_inst_req_0); -- 
    plus_base_ra_3130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_root_address_inst_ack_0, ack => cp_elements(682)); -- 
    plus_base_cr_3131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => array_obj_ref_1008_root_address_inst_req_1); -- 
    plus_base_ca_3132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_root_address_inst_ack_1, ack => cp_elements(683)); -- 
    final_reg_ack_3137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_final_reg_ack_0, ack => cp_elements(684)); -- 
    cpelement_group_685 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(684) & cp_elements(686));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(685),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(685), ack => type_cast_1012_inst_req_0); -- 
    cp_elements(686) <= cp_elements(607);
    cp_elements(687) <= type_cast_1012_inst_ack_0;
    cpelement_group_688 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(667) & cp_elements(687) & cp_elements(704));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(688),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(689) <= cp_elements(687);
    base_resize_req_3160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(689), ack => ptr_deref_1016_base_resize_req_0); -- 
    base_resize_ack_3161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_base_resize_ack_0, ack => cp_elements(690)); -- 
    sum_rename_req_3165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => ptr_deref_1016_root_address_inst_req_0); -- 
    cp_elements(691) <= ptr_deref_1016_root_address_inst_ack_0;
    cp_elements(692) <= cp_elements(691);
    rr_3173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(692), ack => ptr_deref_1016_addr_0_req_0); -- 
    ra_3174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_0_ack_0, ack => cp_elements(693)); -- 
    cr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(693), ack => ptr_deref_1016_addr_0_req_1); -- 
    ca_3176_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_0_ack_1, ack => cp_elements(694)); -- 
    cp_elements(695) <= cp_elements(691);
    rr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(695), ack => ptr_deref_1016_addr_1_req_0); -- 
    ra_3181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_1_ack_0, ack => cp_elements(696)); -- 
    cr_3182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(696), ack => ptr_deref_1016_addr_1_req_1); -- 
    ca_3183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_1_ack_1, ack => cp_elements(697)); -- 
    cp_elements(698) <= cp_elements(691);
    rr_3187_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(698), ack => ptr_deref_1016_addr_2_req_0); -- 
    ra_3188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_2_ack_0, ack => cp_elements(699)); -- 
    cr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => ptr_deref_1016_addr_2_req_1); -- 
    ca_3190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_2_ack_1, ack => cp_elements(700)); -- 
    cp_elements(701) <= cp_elements(691);
    rr_3194_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => ptr_deref_1016_addr_3_req_0); -- 
    ra_3195_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_3_ack_0, ack => cp_elements(702)); -- 
    cr_3196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => ptr_deref_1016_addr_3_req_1); -- 
    ca_3197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_addr_3_ack_1, ack => cp_elements(703)); -- 
    cpelement_group_704 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(694) & cp_elements(697) & cp_elements(700) & cp_elements(703));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(704),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(705) <= cp_elements(688);
    rr_3207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => ptr_deref_1016_load_0_req_0); -- 
    ra_3208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_0_ack_0, ack => cp_elements(706)); -- 
    cp_elements(707) <= cp_elements(688);
    rr_3212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(707), ack => ptr_deref_1016_load_1_req_0); -- 
    ra_3213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_1_ack_0, ack => cp_elements(708)); -- 
    cp_elements(709) <= cp_elements(688);
    rr_3217_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(709), ack => ptr_deref_1016_load_2_req_0); -- 
    ra_3218_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_2_ack_0, ack => cp_elements(710)); -- 
    cp_elements(711) <= cp_elements(688);
    rr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => ptr_deref_1016_load_3_req_0); -- 
    ra_3223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_3_ack_0, ack => cp_elements(712)); -- 
    cpelement_group_713 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(706) & cp_elements(708) & cp_elements(710) & cp_elements(712));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(713),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(714) <= cp_elements(713);
    cp_elements(715) <= cp_elements(714);
    cr_3233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(715), ack => ptr_deref_1016_load_0_req_1); -- 
    ca_3234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_0_ack_1, ack => cp_elements(716)); -- 
    cp_elements(717) <= cp_elements(714);
    cr_3238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(717), ack => ptr_deref_1016_load_1_req_1); -- 
    ca_3239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_1_ack_1, ack => cp_elements(718)); -- 
    cp_elements(719) <= cp_elements(714);
    cr_3243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(719), ack => ptr_deref_1016_load_2_req_1); -- 
    ca_3244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_2_ack_1, ack => cp_elements(720)); -- 
    cp_elements(721) <= cp_elements(714);
    cr_3248_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(721), ack => ptr_deref_1016_load_3_req_1); -- 
    ca_3249_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_3_ack_1, ack => cp_elements(722)); -- 
    cpelement_group_723 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(716) & cp_elements(718) & cp_elements(720) & cp_elements(722));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(723),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_3250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(723), ack => ptr_deref_1016_gather_scatter_req_0); -- 
    merge_ack_3251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_gather_scatter_ack_0, ack => cp_elements(724)); -- 
    cp_elements(725) <= cp_elements(607);
    cpelement_group_726 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(725) & cp_elements(730));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(726),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(726), ack => array_obj_ref_1023_final_reg_req_0); -- 
    cp_elements(727) <= cp_elements(607);
    base_resize_req_3262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => array_obj_ref_1023_base_resize_req_0); -- 
    base_resize_ack_3263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1023_base_resize_ack_0, ack => cp_elements(728)); -- 
    plus_base_rr_3268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => array_obj_ref_1023_root_address_inst_req_0); -- 
    plus_base_ra_3269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1023_root_address_inst_ack_0, ack => cp_elements(729)); -- 
    plus_base_cr_3270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => array_obj_ref_1023_root_address_inst_req_1); -- 
    plus_base_ca_3271_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1023_root_address_inst_ack_1, ack => cp_elements(730)); -- 
    final_reg_ack_3276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1023_final_reg_ack_0, ack => cp_elements(731)); -- 
    cpelement_group_732 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(731) & cp_elements(733));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(732),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(732), ack => type_cast_1027_inst_req_0); -- 
    cp_elements(733) <= cp_elements(607);
    cp_elements(734) <= type_cast_1027_inst_ack_0;
    cpelement_group_735 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(713) & cp_elements(724) & cp_elements(734) & cp_elements(751));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(735),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => ptr_deref_1030_gather_scatter_req_0); -- 
    cp_elements(736) <= cp_elements(734);
    base_resize_req_3300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => ptr_deref_1030_base_resize_req_0); -- 
    base_resize_ack_3301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_base_resize_ack_0, ack => cp_elements(737)); -- 
    sum_rename_req_3305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(737), ack => ptr_deref_1030_root_address_inst_req_0); -- 
    cp_elements(738) <= ptr_deref_1030_root_address_inst_ack_0;
    cp_elements(739) <= cp_elements(738);
    rr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(739), ack => ptr_deref_1030_addr_0_req_0); -- 
    ra_3314_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_0_ack_0, ack => cp_elements(740)); -- 
    cr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => ptr_deref_1030_addr_0_req_1); -- 
    ca_3316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_0_ack_1, ack => cp_elements(741)); -- 
    cp_elements(742) <= cp_elements(738);
    rr_3320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(742), ack => ptr_deref_1030_addr_1_req_0); -- 
    ra_3321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_1_ack_0, ack => cp_elements(743)); -- 
    cr_3322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => ptr_deref_1030_addr_1_req_1); -- 
    ca_3323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_1_ack_1, ack => cp_elements(744)); -- 
    cp_elements(745) <= cp_elements(738);
    rr_3327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => ptr_deref_1030_addr_2_req_0); -- 
    ra_3328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_2_ack_0, ack => cp_elements(746)); -- 
    cr_3329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(746), ack => ptr_deref_1030_addr_2_req_1); -- 
    ca_3330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_2_ack_1, ack => cp_elements(747)); -- 
    cp_elements(748) <= cp_elements(738);
    rr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(748), ack => ptr_deref_1030_addr_3_req_0); -- 
    ra_3335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_3_ack_0, ack => cp_elements(749)); -- 
    cr_3336_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => ptr_deref_1030_addr_3_req_1); -- 
    ca_3337_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_3_ack_1, ack => cp_elements(750)); -- 
    cpelement_group_751 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(741) & cp_elements(744) & cp_elements(747) & cp_elements(750));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(751),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(752) <= ptr_deref_1030_gather_scatter_ack_0;
    cp_elements(753) <= cp_elements(752);
    rr_3349_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => ptr_deref_1030_store_0_req_0); -- 
    ra_3350_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_0_ack_0, ack => cp_elements(754)); -- 
    cp_elements(755) <= cp_elements(752);
    rr_3354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(755), ack => ptr_deref_1030_store_1_req_0); -- 
    ra_3355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_1_ack_0, ack => cp_elements(756)); -- 
    cp_elements(757) <= cp_elements(752);
    rr_3359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(757), ack => ptr_deref_1030_store_2_req_0); -- 
    ra_3360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_2_ack_0, ack => cp_elements(758)); -- 
    cp_elements(759) <= cp_elements(752);
    rr_3364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(759), ack => ptr_deref_1030_store_3_req_0); -- 
    ra_3365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_3_ack_0, ack => cp_elements(760)); -- 
    cpelement_group_761 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(754) & cp_elements(756) & cp_elements(758) & cp_elements(760));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(761),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(762) <= cp_elements(761);
    cr_3375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(762), ack => ptr_deref_1030_store_0_req_1); -- 
    ca_3376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_0_ack_1, ack => cp_elements(763)); -- 
    cp_elements(764) <= cp_elements(761);
    cr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(764), ack => ptr_deref_1030_store_1_req_1); -- 
    ca_3381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_1_ack_1, ack => cp_elements(765)); -- 
    cp_elements(766) <= cp_elements(761);
    cr_3385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(766), ack => ptr_deref_1030_store_2_req_1); -- 
    ca_3386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_2_ack_1, ack => cp_elements(767)); -- 
    cp_elements(768) <= cp_elements(761);
    cr_3390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(768), ack => ptr_deref_1030_store_3_req_1); -- 
    ca_3391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_store_3_ack_1, ack => cp_elements(769)); -- 
    cpelement_group_770 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(763) & cp_elements(765) & cp_elements(767) & cp_elements(769));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(770),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_771 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(677) & cp_elements(770));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(771),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(772) <= cp_elements(606);
    cp_elements(773) <= cp_elements(772);
    cpelement_group_774 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(773) & cp_elements(778));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(774),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => array_obj_ref_1038_final_reg_req_0); -- 
    cp_elements(775) <= cp_elements(772);
    base_resize_req_3405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(775), ack => array_obj_ref_1038_base_resize_req_0); -- 
    base_resize_ack_3406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_base_resize_ack_0, ack => cp_elements(776)); -- 
    plus_base_rr_3411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => array_obj_ref_1038_root_address_inst_req_0); -- 
    plus_base_ra_3412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_root_address_inst_ack_0, ack => cp_elements(777)); -- 
    plus_base_cr_3413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(777), ack => array_obj_ref_1038_root_address_inst_req_1); -- 
    plus_base_ca_3414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_root_address_inst_ack_1, ack => cp_elements(778)); -- 
    final_reg_ack_3419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_final_reg_ack_0, ack => cp_elements(779)); -- 
    cpelement_group_780 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(779) & cp_elements(781));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(780),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(780), ack => type_cast_1042_inst_req_0); -- 
    cp_elements(781) <= cp_elements(772);
    cp_elements(782) <= type_cast_1042_inst_ack_0;
    cpelement_group_783 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(782) & cp_elements(799));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(783),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(784) <= cp_elements(782);
    base_resize_req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => ptr_deref_1046_base_resize_req_0); -- 
    base_resize_ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_base_resize_ack_0, ack => cp_elements(785)); -- 
    sum_rename_req_3447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => ptr_deref_1046_root_address_inst_req_0); -- 
    cp_elements(786) <= ptr_deref_1046_root_address_inst_ack_0;
    cp_elements(787) <= cp_elements(786);
    rr_3455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(787), ack => ptr_deref_1046_addr_0_req_0); -- 
    ra_3456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_0_ack_0, ack => cp_elements(788)); -- 
    cr_3457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(788), ack => ptr_deref_1046_addr_0_req_1); -- 
    ca_3458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_0_ack_1, ack => cp_elements(789)); -- 
    cp_elements(790) <= cp_elements(786);
    rr_3462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => ptr_deref_1046_addr_1_req_0); -- 
    ra_3463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_1_ack_0, ack => cp_elements(791)); -- 
    cr_3464_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => ptr_deref_1046_addr_1_req_1); -- 
    ca_3465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_1_ack_1, ack => cp_elements(792)); -- 
    cp_elements(793) <= cp_elements(786);
    rr_3469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(793), ack => ptr_deref_1046_addr_2_req_0); -- 
    ra_3470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_2_ack_0, ack => cp_elements(794)); -- 
    cr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => ptr_deref_1046_addr_2_req_1); -- 
    ca_3472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_2_ack_1, ack => cp_elements(795)); -- 
    cp_elements(796) <= cp_elements(786);
    rr_3476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => ptr_deref_1046_addr_3_req_0); -- 
    ra_3477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_3_ack_0, ack => cp_elements(797)); -- 
    cr_3478_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => ptr_deref_1046_addr_3_req_1); -- 
    ca_3479_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_3_ack_1, ack => cp_elements(798)); -- 
    cpelement_group_799 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(789) & cp_elements(792) & cp_elements(795) & cp_elements(798));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(799),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(800) <= cp_elements(783);
    rr_3489_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(800), ack => ptr_deref_1046_load_0_req_0); -- 
    ra_3490_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_0_ack_0, ack => cp_elements(801)); -- 
    cp_elements(802) <= cp_elements(783);
    rr_3494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(802), ack => ptr_deref_1046_load_1_req_0); -- 
    ra_3495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_1_ack_0, ack => cp_elements(803)); -- 
    cp_elements(804) <= cp_elements(783);
    rr_3499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(804), ack => ptr_deref_1046_load_2_req_0); -- 
    ra_3500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_2_ack_0, ack => cp_elements(805)); -- 
    cp_elements(806) <= cp_elements(783);
    rr_3504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => ptr_deref_1046_load_3_req_0); -- 
    ra_3505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_3_ack_0, ack => cp_elements(807)); -- 
    cpelement_group_808 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(801) & cp_elements(803) & cp_elements(805) & cp_elements(807));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(808),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(809) <= cp_elements(808);
    cp_elements(810) <= cp_elements(809);
    cr_3515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => ptr_deref_1046_load_0_req_1); -- 
    ca_3516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_0_ack_1, ack => cp_elements(811)); -- 
    cp_elements(812) <= cp_elements(809);
    cr_3520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(812), ack => ptr_deref_1046_load_1_req_1); -- 
    ca_3521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_1_ack_1, ack => cp_elements(813)); -- 
    cp_elements(814) <= cp_elements(809);
    cr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(814), ack => ptr_deref_1046_load_2_req_1); -- 
    ca_3526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_2_ack_1, ack => cp_elements(815)); -- 
    cp_elements(816) <= cp_elements(809);
    cr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(816), ack => ptr_deref_1046_load_3_req_1); -- 
    ca_3531_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_load_3_ack_1, ack => cp_elements(817)); -- 
    cpelement_group_818 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(811) & cp_elements(813) & cp_elements(815) & cp_elements(817));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(818),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(818), ack => ptr_deref_1046_gather_scatter_req_0); -- 
    merge_ack_3533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_gather_scatter_ack_0, ack => cp_elements(819)); -- 
    cp_elements(820) <= cp_elements(772);
    cpelement_group_821 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(820) & cp_elements(825));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(821),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(821), ack => array_obj_ref_1053_final_reg_req_0); -- 
    cp_elements(822) <= cp_elements(772);
    base_resize_req_3544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(822), ack => array_obj_ref_1053_base_resize_req_0); -- 
    base_resize_ack_3545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1053_base_resize_ack_0, ack => cp_elements(823)); -- 
    plus_base_rr_3550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(823), ack => array_obj_ref_1053_root_address_inst_req_0); -- 
    plus_base_ra_3551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1053_root_address_inst_ack_0, ack => cp_elements(824)); -- 
    plus_base_cr_3552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(824), ack => array_obj_ref_1053_root_address_inst_req_1); -- 
    plus_base_ca_3553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1053_root_address_inst_ack_1, ack => cp_elements(825)); -- 
    final_reg_ack_3558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1053_final_reg_ack_0, ack => cp_elements(826)); -- 
    cpelement_group_827 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(826) & cp_elements(828));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(827),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(827), ack => type_cast_1057_inst_req_0); -- 
    cp_elements(828) <= cp_elements(772);
    cp_elements(829) <= type_cast_1057_inst_ack_0;
    cpelement_group_830 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(808) & cp_elements(819) & cp_elements(829) & cp_elements(846));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(830),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(830), ack => ptr_deref_1060_gather_scatter_req_0); -- 
    cp_elements(831) <= cp_elements(829);
    base_resize_req_3582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(831), ack => ptr_deref_1060_base_resize_req_0); -- 
    base_resize_ack_3583_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_base_resize_ack_0, ack => cp_elements(832)); -- 
    sum_rename_req_3587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(832), ack => ptr_deref_1060_root_address_inst_req_0); -- 
    cp_elements(833) <= ptr_deref_1060_root_address_inst_ack_0;
    cp_elements(834) <= cp_elements(833);
    rr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(834), ack => ptr_deref_1060_addr_0_req_0); -- 
    ra_3596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_0_ack_0, ack => cp_elements(835)); -- 
    cr_3597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => ptr_deref_1060_addr_0_req_1); -- 
    ca_3598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_0_ack_1, ack => cp_elements(836)); -- 
    cp_elements(837) <= cp_elements(833);
    rr_3602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(837), ack => ptr_deref_1060_addr_1_req_0); -- 
    ra_3603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_1_ack_0, ack => cp_elements(838)); -- 
    cr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(838), ack => ptr_deref_1060_addr_1_req_1); -- 
    ca_3605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_1_ack_1, ack => cp_elements(839)); -- 
    cp_elements(840) <= cp_elements(833);
    rr_3609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => ptr_deref_1060_addr_2_req_0); -- 
    ra_3610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_2_ack_0, ack => cp_elements(841)); -- 
    cr_3611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(841), ack => ptr_deref_1060_addr_2_req_1); -- 
    ca_3612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_2_ack_1, ack => cp_elements(842)); -- 
    cp_elements(843) <= cp_elements(833);
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(843), ack => ptr_deref_1060_addr_3_req_0); -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_3_ack_0, ack => cp_elements(844)); -- 
    cr_3618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(844), ack => ptr_deref_1060_addr_3_req_1); -- 
    ca_3619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_addr_3_ack_1, ack => cp_elements(845)); -- 
    cpelement_group_846 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(836) & cp_elements(839) & cp_elements(842) & cp_elements(845));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(846),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(847) <= ptr_deref_1060_gather_scatter_ack_0;
    cp_elements(848) <= cp_elements(847);
    rr_3631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(848), ack => ptr_deref_1060_store_0_req_0); -- 
    ra_3632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_0_ack_0, ack => cp_elements(849)); -- 
    cp_elements(850) <= cp_elements(847);
    rr_3636_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(850), ack => ptr_deref_1060_store_1_req_0); -- 
    ra_3637_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_1_ack_0, ack => cp_elements(851)); -- 
    cp_elements(852) <= cp_elements(847);
    rr_3641_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(852), ack => ptr_deref_1060_store_2_req_0); -- 
    ra_3642_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_2_ack_0, ack => cp_elements(853)); -- 
    cp_elements(854) <= cp_elements(847);
    rr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(854), ack => ptr_deref_1060_store_3_req_0); -- 
    ra_3647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_3_ack_0, ack => cp_elements(855)); -- 
    cpelement_group_856 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(849) & cp_elements(851) & cp_elements(853) & cp_elements(855));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(856),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(857) <= cp_elements(856);
    cr_3657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(857), ack => ptr_deref_1060_store_0_req_1); -- 
    ca_3658_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_0_ack_1, ack => cp_elements(858)); -- 
    cp_elements(859) <= cp_elements(856);
    cr_3662_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(859), ack => ptr_deref_1060_store_1_req_1); -- 
    ca_3663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_1_ack_1, ack => cp_elements(860)); -- 
    cp_elements(861) <= cp_elements(856);
    cr_3667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(861), ack => ptr_deref_1060_store_2_req_1); -- 
    ca_3668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_2_ack_1, ack => cp_elements(862)); -- 
    cp_elements(863) <= cp_elements(856);
    cr_3672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(863), ack => ptr_deref_1060_store_3_req_1); -- 
    ca_3673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1060_store_3_ack_1, ack => cp_elements(864)); -- 
    cpelement_group_865 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(858) & cp_elements(860) & cp_elements(862) & cp_elements(864));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(865),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_866 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(867) & cp_elements(868));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(866),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_3682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(866), ack => binary_1067_inst_req_0); -- 
    cp_elements(867) <= cp_elements(772);
    cp_elements(868) <= cp_elements(772);
    ra_3683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1067_inst_ack_0, ack => cp_elements(869)); -- 
    cr_3684_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(869), ack => binary_1067_inst_req_1); -- 
    ca_3685_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1067_inst_ack_1, ack => cp_elements(870)); -- 
    cpelement_group_871 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(865) & cp_elements(870));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(871),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(872) <= cp_elements(17);
    cp_elements(873) <= false;
    cp_elements(874) <= cp_elements(873);
    cp_elements(875) <= cp_elements(17);
    branch_req_3693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(875), ack => if_stmt_1069_branch_req_0); -- 
    cp_elements(876) <= cp_elements(875);
    cp_elements(877) <= cp_elements(876);
    if_choice_transition_3698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1069_branch_ack_1, ack => cp_elements(878)); -- 
    cp_elements(879) <= cp_elements(876);
    else_choice_transition_3702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1069_branch_ack_0, ack => cp_elements(880)); -- 
    cp_elements(881) <= cp_elements(18);
    cpelement_group_882 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(883) & cp_elements(884));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(882),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(882), ack => type_cast_1078_inst_req_0); -- 
    cp_elements(883) <= cp_elements(881);
    cp_elements(884) <= cp_elements(881);
    ack_3717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1078_inst_ack_0, ack => cp_elements(885)); -- 
    cp_elements(886) <= cp_elements(885);
    cpelement_group_887 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(888) & cp_elements(889));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(887),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(887), ack => type_cast_1082_inst_req_0); -- 
    cp_elements(888) <= cp_elements(886);
    cp_elements(889) <= cp_elements(886);
    ack_3730_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1082_inst_ack_0, ack => cp_elements(890)); -- 
    pipe_wreq_3735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(890), ack => simple_obj_ref_1080_inst_req_0); -- 
    pipe_wack_3736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1080_inst_ack_0, ack => cp_elements(891)); -- 
    cp_elements(892) <= false;
    cp_elements(893) <= cp_elements(892);
    cp_elements(894) <= false;
    cp_elements(895) <= cp_elements(894);
    cp_elements(896) <= false;
    cp_elements(897) <= cp_elements(896);
    cp_elements(898) <= false;
    cp_elements(899) <= cp_elements(898);
    cp_elements(900) <= false;
    cp_elements(901) <= cp_elements(900);
    cp_elements(902) <= cp_elements(390);
    cp_elements(903) <= cp_elements(902);
    req_3841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(903), ack => type_cast_740_inst_req_0); -- 
    ack_3842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_0, ack => cp_elements(904)); -- 
    phi_stmt_734_req_3843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(904), ack => phi_stmt_734_req_1); -- 
    cp_elements(905) <= cp_elements(902);
    req_3853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(905), ack => type_cast_747_inst_req_0); -- 
    ack_3854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_0, ack => cp_elements(906)); -- 
    phi_stmt_741_req_3855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(906), ack => phi_stmt_741_req_1); -- 
    cpelement_group_907 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(904) & cp_elements(906));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(907),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(908) <= cp_elements(306);
    cp_elements(909) <= cp_elements(908);
    phi_stmt_734_req_3870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(909), ack => phi_stmt_734_req_0); -- 
    cp_elements(910) <= cp_elements(908);
    phi_stmt_741_req_3882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(910), ack => phi_stmt_741_req_0); -- 
    cpelement_group_911 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(909) & cp_elements(910));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(911),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(912) <= OrReduce(cp_elements(907) & cp_elements(911));
    cp_elements(913) <= cp_elements(912);
    phi_stmt_734_ack_3887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_734_ack_0, ack => cp_elements(914)); -- 
    phi_stmt_741_ack_3888_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_741_ack_0, ack => cp_elements(915)); -- 
    cpelement_group_916 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(914) & cp_elements(915));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(916),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(917) <= false;
    cp_elements(918) <= cp_elements(917);
    cp_elements(919) <= cp_elements(300);
    cp_elements(920) <= cp_elements(919);
    phi_stmt_827_req_3915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(920), ack => phi_stmt_827_req_1); -- 
    cp_elements(921) <= cp_elements(919);
    cp_elements(922) <= cp_elements(921);
    cp_elements(923) <= cp_elements(921);
    req_3930_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(923), ack => type_cast_839_inst_req_0); -- 
    ack_3931_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_0, ack => cp_elements(924)); -- 
    cpelement_group_925 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(922) & cp_elements(924));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(925),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_834_req_3932_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(925), ack => phi_stmt_834_req_1); -- 
    cp_elements(926) <= cp_elements(919);
    cp_elements(927) <= cp_elements(926);
    cp_elements(928) <= cp_elements(926);
    req_3947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(928), ack => type_cast_845_inst_req_0); -- 
    ack_3948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_845_inst_ack_0, ack => cp_elements(929)); -- 
    cpelement_group_930 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(927) & cp_elements(929));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(930),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_840_req_3949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(930), ack => phi_stmt_840_req_1); -- 
    cpelement_group_931 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(920) & cp_elements(925) & cp_elements(930));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(931),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(932) <= cp_elements(409);
    cp_elements(933) <= cp_elements(932);
    req_3962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(933), ack => type_cast_830_inst_req_0); -- 
    ack_3963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_830_inst_ack_0, ack => cp_elements(934)); -- 
    phi_stmt_827_req_3964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(934), ack => phi_stmt_827_req_0); -- 
    cp_elements(935) <= cp_elements(932);
    cp_elements(936) <= cp_elements(935);
    req_3974_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(936), ack => type_cast_837_inst_req_0); -- 
    ack_3975_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_0, ack => cp_elements(937)); -- 
    cp_elements(938) <= cp_elements(935);
    cpelement_group_939 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(937) & cp_elements(938));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(939),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_834_req_3981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => phi_stmt_834_req_0); -- 
    cp_elements(940) <= cp_elements(932);
    cp_elements(941) <= cp_elements(940);
    req_3991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(941), ack => type_cast_843_inst_req_0); -- 
    ack_3992_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_0, ack => cp_elements(942)); -- 
    cp_elements(943) <= cp_elements(940);
    cpelement_group_944 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(942) & cp_elements(943));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(944),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_840_req_3998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => phi_stmt_840_req_0); -- 
    cpelement_group_945 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(934) & cp_elements(939) & cp_elements(944));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(945),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(946) <= OrReduce(cp_elements(931) & cp_elements(945));
    cp_elements(947) <= cp_elements(946);
    phi_stmt_827_ack_4003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_827_ack_0, ack => cp_elements(948)); -- 
    phi_stmt_834_ack_4004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_834_ack_0, ack => cp_elements(949)); -- 
    phi_stmt_840_ack_4005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_840_ack_0, ack => cp_elements(950)); -- 
    cpelement_group_951 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(948) & cp_elements(949) & cp_elements(950));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(951),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(952) <= false;
    cp_elements(953) <= cp_elements(952);
    cp_elements(954) <= cp_elements(424);
    cp_elements(955) <= cp_elements(424);
    req_4035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(955), ack => type_cast_880_inst_req_0); -- 
    ack_4036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_0, ack => cp_elements(956)); -- 
    cpelement_group_957 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(954) & cp_elements(956));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(957),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_875_req_4037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(957), ack => phi_stmt_875_req_1); -- 
    cp_elements(958) <= cp_elements(442);
    req_4050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(958), ack => type_cast_878_inst_req_0); -- 
    ack_4051_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_0, ack => cp_elements(959)); -- 
    cp_elements(960) <= cp_elements(442);
    cpelement_group_961 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(959) & cp_elements(960));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(961),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_875_req_4057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(961), ack => phi_stmt_875_req_0); -- 
    cp_elements(962) <= OrReduce(cp_elements(957) & cp_elements(961));
    cp_elements(963) <= cp_elements(962);
    phi_stmt_875_ack_4062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_875_ack_0, ack => cp_elements(964)); -- 
    cp_elements(965) <= false;
    cp_elements(966) <= cp_elements(965);
    cp_elements(967) <= false;
    cp_elements(968) <= cp_elements(967);
    cp_elements(969) <= false;
    cp_elements(970) <= cp_elements(969);
    cp_elements(971) <= OrReduce(cp_elements(16) & cp_elements(880));
    cp_elements(972) <= cp_elements(971);
    cp_elements(973) <= OrReduce(cp_elements(156) & cp_elements(226) & cp_elements(251) & cp_elements(285) & cp_elements(485) & cp_elements(878) & cp_elements(891));
    cp_elements(974) <= cp_elements(973);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1008_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1008_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1008_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1023_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1023_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1023_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1038_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1038_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1038_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1053_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1053_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1053_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_549_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_549_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_549_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_558_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_558_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_558_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_565_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_565_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_565_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_774_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_774_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_774_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_774_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_823_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_823_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_823_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_823_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_936_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_936_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_936_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_950_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_950_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_950_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_950_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_957_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_957_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_957_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_999_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_999_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_999_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_999_root_address : std_logic_vector(15 downto 0);
    signal elt5x_xi11_1013 : std_logic_vector(31 downto 0);
    signal elt5x_xi_1043 : std_logic_vector(31 downto 0);
    signal indvarx_xi12x_xi_734 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xi14x_xi_807 : std_logic_vector(31 downto 0);
    signal orx_xcondx_xi_701 : std_logic_vector(0 downto 0);
    signal ptr_deref_1002_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1002_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1002_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1002_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1002_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1002_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1002_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1016_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1016_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1016_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1016_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1030_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1030_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1030_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1030_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1030_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1030_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1046_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1046_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1046_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1046_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1046_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1060_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1060_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1060_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1060_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1060_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1060_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_553_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_569_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_616_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_616_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_616_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_616_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_616_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_616_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_783_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_783_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_783_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_783_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_783_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_783_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_783_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_783_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_862_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_862_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_862_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_862_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_862_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_939_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_939_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_939_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_939_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_939_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_939_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_939_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_939_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_960_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_960_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_960_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_960_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_960_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_960_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_960_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_960_word_offset_3 : std_logic_vector(15 downto 0);
    signal scevgep12x_xix_xi_780 : std_logic_vector(31 downto 0);
    signal scevgep14x_xix_xi_824 : std_logic_vector(31 downto 0);
    signal scevgep_775 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_537_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_773_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_773_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_822_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_822_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_949_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_949_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_998_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_998_scaled : std_logic_vector(15 downto 0);
    signal tmp13_539 : std_logic_vector(31 downto 0);
    signal tmp14_543 : std_logic_vector(31 downto 0);
    signal tmp15_550 : std_logic_vector(31 downto 0);
    signal tmp16_554 : std_logic_vector(31 downto 0);
    signal tmp17_559 : std_logic_vector(31 downto 0);
    signal tmp17x_xix_xi_759 : std_logic_vector(31 downto 0);
    signal tmp18_566 : std_logic_vector(31 downto 0);
    signal tmp19_570 : std_logic_vector(31 downto 0);
    signal tmp20_574 : std_logic_vector(31 downto 0);
    signal tmp21_578 : std_logic_vector(31 downto 0);
    signal tmp22_583 : std_logic_vector(31 downto 0);
    signal tmp23_589 : std_logic_vector(31 downto 0);
    signal tmp24_598 : std_logic_vector(0 downto 0);
    signal tmp25_613 : std_logic_vector(31 downto 0);
    signal tmp26_617 : std_logic_vector(31 downto 0);
    signal tmp27_623 : std_logic_vector(31 downto 0);
    signal tmp28_629 : std_logic_vector(0 downto 0);
    signal tmp29_656 : std_logic_vector(31 downto 0);
    signal tmp30_662 : std_logic_vector(31 downto 0);
    signal tmp31_668 : std_logic_vector(0 downto 0);
    signal tmp32_682 : std_logic_vector(15 downto 0);
    signal tmp33_686 : std_logic_vector(31 downto 0);
    signal tmp34_691 : std_logic_vector(0 downto 0);
    signal tmp34x_xi_635 : std_logic_vector(31 downto 0);
    signal tmp35_696 : std_logic_vector(0 downto 0);
    signal tmp35x_xi_639 : std_logic_vector(15 downto 0);
    signal tmp36_718 : std_logic_vector(0 downto 0);
    signal tmp37_741 : std_logic_vector(31 downto 0);
    signal tmp38_784 : std_logic_vector(15 downto 0);
    signal tmp39_788 : std_logic_vector(31 downto 0);
    signal tmp40_793 : std_logic_vector(31 downto 0);
    signal tmp41_801 : std_logic_vector(0 downto 0);
    signal tmp42_852 : std_logic_vector(0 downto 0);
    signal tmp43_863 : std_logic_vector(7 downto 0);
    signal tmp44_867 : std_logic_vector(31 downto 0);
    signal tmp45_872 : std_logic_vector(31 downto 0);
    signal tmp46_875 : std_logic_vector(31 downto 0);
    signal tmp47_887 : std_logic_vector(31 downto 0);
    signal tmp48_893 : std_logic_vector(31 downto 0);
    signal tmp49_898 : std_logic_vector(31 downto 0);
    signal tmp50_904 : std_logic_vector(31 downto 0);
    signal tmp51_909 : std_logic_vector(31 downto 0);
    signal tmp52_913 : std_logic_vector(15 downto 0);
    signal tmp53_919 : std_logic_vector(0 downto 0);
    signal tmp54_937 : std_logic_vector(31 downto 0);
    signal tmp55_951 : std_logic_vector(31 downto 0);
    signal tmp56_958 : std_logic_vector(31 downto 0);
    signal tmp57_967 : std_logic_vector(0 downto 0);
    signal tmp58_979 : std_logic_vector(31 downto 0);
    signal tmp59_984 : std_logic_vector(0 downto 0);
    signal tmp5_731 : std_logic_vector(31 downto 0);
    signal tmp60_990 : std_logic_vector(31 downto 0);
    signal tmp61_996 : std_logic_vector(31 downto 0);
    signal tmp62_1000 : std_logic_vector(31 downto 0);
    signal tmp63_1009 : std_logic_vector(31 downto 0);
    signal tmp64_1024 : std_logic_vector(31 downto 0);
    signal tmp65_1028 : std_logic_vector(31 downto 0);
    signal tmp66_1039 : std_logic_vector(31 downto 0);
    signal tmp67_1054 : std_logic_vector(31 downto 0);
    signal tmp68_1058 : std_logic_vector(31 downto 0);
    signal tmp69_1068 : std_logic_vector(0 downto 0);
    signal tmp70_1079 : std_logic_vector(31 downto 0);
    signal tmp8_771 : std_logic_vector(31 downto 0);
    signal tmp_754 : std_logic_vector(31 downto 0);
    signal tmpx_xix_xi_765 : std_logic_vector(31 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1082_wire : std_logic_vector(31 downto 0);
    signal type_cast_587_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_593_wire : std_logic_vector(31 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_621_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_627_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_633_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_666_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_729_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_740_wire : std_logic_vector(31 downto 0);
    signal type_cast_745_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_747_wire : std_logic_vector(31 downto 0);
    signal type_cast_752_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_763_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_769_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_796_wire : std_logic_vector(31 downto 0);
    signal type_cast_799_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_805_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_818_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_830_wire : std_logic_vector(31 downto 0);
    signal type_cast_833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_837_wire : std_logic_vector(31 downto 0);
    signal type_cast_839_wire : std_logic_vector(31 downto 0);
    signal type_cast_843_wire : std_logic_vector(31 downto 0);
    signal type_cast_845_wire : std_logic_vector(31 downto 0);
    signal type_cast_850_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_878_wire : std_logic_vector(31 downto 0);
    signal type_cast_880_wire : std_logic_vector(31 downto 0);
    signal type_cast_885_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_902_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_917_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_945_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_993_wire_constant : std_logic_vector(31 downto 0);
    signal val6x_xi12_1017 : std_logic_vector(31 downto 0);
    signal val6x_xi_1047 : std_logic_vector(31 downto 0);
    signal xx_xinx_xlcssax_xix_xi_834 : std_logic_vector(31 downto 0);
    signal xx_xlcssa5x_xix_xi_827 : std_logic_vector(31 downto 0);
    signal xx_xlcssax_xix_xi_840 : std_logic_vector(31 downto 0);
    signal xx_xsum20x_xi_820 : std_logic_vector(31 downto 0);
    signal xx_xsumx_xi_947 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1008_final_offset <= "0000000000011110";
    array_obj_ref_1023_final_offset <= "0000000000011100";
    array_obj_ref_1038_final_offset <= "0000000000011110";
    array_obj_ref_1053_final_offset <= "0000000000011100";
    array_obj_ref_549_final_offset <= "0000000000001100";
    array_obj_ref_558_final_offset <= "0000000000001110";
    array_obj_ref_565_final_offset <= "0000000000010000";
    array_obj_ref_774_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_823_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_936_final_offset <= "0000000001010000";
    array_obj_ref_950_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_957_final_offset <= "0000000001010100";
    array_obj_ref_999_offset_scale_factor_0 <= "0000000000000001";
    ptr_deref_1002_word_offset_0 <= "0000000000000000";
    ptr_deref_1002_word_offset_1 <= "0000000000000001";
    ptr_deref_1002_word_offset_2 <= "0000000000000010";
    ptr_deref_1002_word_offset_3 <= "0000000000000011";
    ptr_deref_1016_word_offset_0 <= "0000000000000000";
    ptr_deref_1016_word_offset_1 <= "0000000000000001";
    ptr_deref_1016_word_offset_2 <= "0000000000000010";
    ptr_deref_1016_word_offset_3 <= "0000000000000011";
    ptr_deref_1030_word_offset_0 <= "0000000000000000";
    ptr_deref_1030_word_offset_1 <= "0000000000000001";
    ptr_deref_1030_word_offset_2 <= "0000000000000010";
    ptr_deref_1030_word_offset_3 <= "0000000000000011";
    ptr_deref_1046_word_offset_0 <= "0000000000000000";
    ptr_deref_1046_word_offset_1 <= "0000000000000001";
    ptr_deref_1046_word_offset_2 <= "0000000000000010";
    ptr_deref_1046_word_offset_3 <= "0000000000000011";
    ptr_deref_1060_word_offset_0 <= "0000000000000000";
    ptr_deref_1060_word_offset_1 <= "0000000000000001";
    ptr_deref_1060_word_offset_2 <= "0000000000000010";
    ptr_deref_1060_word_offset_3 <= "0000000000000011";
    ptr_deref_553_word_offset_0 <= "0000000000000000";
    ptr_deref_553_word_offset_1 <= "0000000000000001";
    ptr_deref_553_word_offset_2 <= "0000000000000010";
    ptr_deref_553_word_offset_3 <= "0000000000000011";
    ptr_deref_569_word_offset_0 <= "0000000000000000";
    ptr_deref_569_word_offset_1 <= "0000000000000001";
    ptr_deref_569_word_offset_2 <= "0000000000000010";
    ptr_deref_569_word_offset_3 <= "0000000000000011";
    ptr_deref_616_word_offset_0 <= "0000000000000000";
    ptr_deref_616_word_offset_1 <= "0000000000000001";
    ptr_deref_616_word_offset_2 <= "0000000000000010";
    ptr_deref_616_word_offset_3 <= "0000000000000011";
    ptr_deref_783_word_offset_0 <= "0000000000000000";
    ptr_deref_783_word_offset_1 <= "0000000000000001";
    ptr_deref_862_word_offset_0 <= "0000000000000000";
    ptr_deref_939_word_offset_0 <= "0000000000000000";
    ptr_deref_939_word_offset_1 <= "0000000000000001";
    ptr_deref_939_word_offset_2 <= "0000000000000010";
    ptr_deref_939_word_offset_3 <= "0000000000000011";
    ptr_deref_960_word_offset_0 <= "0000000000000000";
    ptr_deref_960_word_offset_1 <= "0000000000000001";
    ptr_deref_960_word_offset_2 <= "0000000000000010";
    ptr_deref_960_word_offset_3 <= "0000000000000011";
    type_cast_1066_wire_constant <= "11111111111111111111111111111111";
    type_cast_587_wire_constant <= "11111111111111111111111111110010";
    type_cast_596_wire_constant <= "00000000000000000000000000010100";
    type_cast_621_wire_constant <= "00000000000000000000000011110000";
    type_cast_627_wire_constant <= "00000000000000000000000001000000";
    type_cast_633_wire_constant <= "00000000000000000000000000010000";
    type_cast_654_wire_constant <= "00000000000000000000000000000010";
    type_cast_660_wire_constant <= "00000000000000000000000000111100";
    type_cast_666_wire_constant <= "00000000000000000000000000010100";
    type_cast_716_wire_constant <= "00000000000000000000000000000001";
    type_cast_729_wire_constant <= "11111111111111111111111111111110";
    type_cast_738_wire_constant <= "00000000000000000000000000000000";
    type_cast_745_wire_constant <= "00000000000000000000000000000000";
    type_cast_752_wire_constant <= "11111111111111111111111111111110";
    type_cast_763_wire_constant <= "00000000000000000000000000000001";
    type_cast_769_wire_constant <= "00000000000000000000000000001110";
    type_cast_799_wire_constant <= "00000000000000000000000000000001";
    type_cast_805_wire_constant <= "00000000000000000000000000000001";
    type_cast_818_wire_constant <= "00000000000000000000000000010000";
    type_cast_833_wire_constant <= "00000000000000000000000000000000";
    type_cast_850_wire_constant <= "00000000000000000000000000000001";
    type_cast_885_wire_constant <= "00000000000000001111111111111111";
    type_cast_891_wire_constant <= "00000000000000000000000000010000";
    type_cast_902_wire_constant <= "00000000000000000000000000010000";
    type_cast_917_wire_constant <= "1111111111111111";
    type_cast_945_wire_constant <= "00000000000000000000000000001110";
    type_cast_993_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_734: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_738_wire_constant & type_cast_740_wire;
      req <= phi_stmt_734_req_0 & phi_stmt_734_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_734_ack_0,
          idata => idata,
          odata => indvarx_xi12x_xi_734,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_734
    phi_stmt_741: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_745_wire_constant & type_cast_747_wire;
      req <= phi_stmt_741_req_0 & phi_stmt_741_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_741_ack_0,
          idata => idata,
          odata => tmp37_741,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_741
    phi_stmt_827: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_830_wire & type_cast_833_wire_constant;
      req <= phi_stmt_827_req_0 & phi_stmt_827_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_827_ack_0,
          idata => idata,
          odata => xx_xlcssa5x_xix_xi_827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_827
    phi_stmt_834: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_837_wire & type_cast_839_wire;
      req <= phi_stmt_834_req_0 & phi_stmt_834_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_834_ack_0,
          idata => idata,
          odata => xx_xinx_xlcssax_xix_xi_834,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_834
    phi_stmt_840: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_843_wire & type_cast_845_wire;
      req <= phi_stmt_840_req_0 & phi_stmt_840_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_840_ack_0,
          idata => idata,
          odata => xx_xlcssax_xix_xi_840,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_840
    phi_stmt_875: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_878_wire & type_cast_880_wire;
      req <= phi_stmt_875_req_0 & phi_stmt_875_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_875_ack_0,
          idata => idata,
          odata => tmp46_875,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_875
    ternary_989_inst: SelectBase generic map(data_width => 32) -- 
      port map( x => tmp22_583, y => tmp58_979, sel => tmp59_984, z => tmp60_990, req => ternary_989_inst_req_0, ack => ternary_989_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1008_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_1008_resized_base_address, req => array_obj_ref_1008_base_resize_req_0, ack => array_obj_ref_1008_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1008_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1008_root_address, dout => tmp63_1009, req => array_obj_ref_1008_final_reg_req_0, ack => array_obj_ref_1008_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1023_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_1023_resized_base_address, req => array_obj_ref_1023_base_resize_req_0, ack => array_obj_ref_1023_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1023_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1023_root_address, dout => tmp64_1024, req => array_obj_ref_1023_final_reg_req_0, ack => array_obj_ref_1023_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1038_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_1038_resized_base_address, req => array_obj_ref_1038_base_resize_req_0, ack => array_obj_ref_1038_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1038_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1038_root_address, dout => tmp66_1039, req => array_obj_ref_1038_final_reg_req_0, ack => array_obj_ref_1038_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1053_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_1053_resized_base_address, req => array_obj_ref_1053_base_resize_req_0, ack => array_obj_ref_1053_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1053_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1053_root_address, dout => tmp67_1054, req => array_obj_ref_1053_final_reg_req_0, ack => array_obj_ref_1053_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_549_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_549_resized_base_address, req => array_obj_ref_549_base_resize_req_0, ack => array_obj_ref_549_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_549_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_549_root_address, dout => tmp15_550, req => array_obj_ref_549_final_reg_req_0, ack => array_obj_ref_549_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_558_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_558_resized_base_address, req => array_obj_ref_558_base_resize_req_0, ack => array_obj_ref_558_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_558_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_558_root_address, dout => tmp17_559, req => array_obj_ref_558_final_reg_req_0, ack => array_obj_ref_558_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_565_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_565_resized_base_address, req => array_obj_ref_565_base_resize_req_0, ack => array_obj_ref_565_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_565_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_565_root_address, dout => tmp18_566, req => array_obj_ref_565_final_reg_req_0, ack => array_obj_ref_565_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_774_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_774_resized_base_address, req => array_obj_ref_774_base_resize_req_0, ack => array_obj_ref_774_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_774_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_774_root_address, dout => scevgep_775, req => array_obj_ref_774_final_reg_req_0, ack => array_obj_ref_774_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_774_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_771, dout => simple_obj_ref_773_resized, req => array_obj_ref_774_index_0_resize_req_0, ack => array_obj_ref_774_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_774_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_773_scaled, dout => array_obj_ref_774_final_offset, req => array_obj_ref_774_offset_inst_req_0, ack => array_obj_ref_774_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_823_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_823_resized_base_address, req => array_obj_ref_823_base_resize_req_0, ack => array_obj_ref_823_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_823_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_823_root_address, dout => scevgep14x_xix_xi_824, req => array_obj_ref_823_final_reg_req_0, ack => array_obj_ref_823_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_823_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xsum20x_xi_820, dout => simple_obj_ref_822_resized, req => array_obj_ref_823_index_0_resize_req_0, ack => array_obj_ref_823_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_823_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_822_scaled, dout => array_obj_ref_823_final_offset, req => array_obj_ref_823_offset_inst_req_0, ack => array_obj_ref_823_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_936_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_936_resized_base_address, req => array_obj_ref_936_base_resize_req_0, ack => array_obj_ref_936_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_936_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_936_root_address, dout => tmp54_937, req => array_obj_ref_936_final_reg_req_0, ack => array_obj_ref_936_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_950_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_950_resized_base_address, req => array_obj_ref_950_base_resize_req_0, ack => array_obj_ref_950_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_950_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_950_root_address, dout => tmp55_951, req => array_obj_ref_950_final_reg_req_0, ack => array_obj_ref_950_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_950_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xsumx_xi_947, dout => simple_obj_ref_949_resized, req => array_obj_ref_950_index_0_resize_req_0, ack => array_obj_ref_950_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_950_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_949_scaled, dout => array_obj_ref_950_final_offset, req => array_obj_ref_950_offset_inst_req_0, ack => array_obj_ref_950_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_957_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_957_resized_base_address, req => array_obj_ref_957_base_resize_req_0, ack => array_obj_ref_957_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_957_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_957_root_address, dout => tmp56_958, req => array_obj_ref_957_final_reg_req_0, ack => array_obj_ref_957_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_999_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp19_570, dout => array_obj_ref_999_resized_base_address, req => array_obj_ref_999_base_resize_req_0, ack => array_obj_ref_999_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_999_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_999_root_address, dout => tmp62_1000, req => array_obj_ref_999_final_reg_req_0, ack => array_obj_ref_999_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_999_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp61_996, dout => simple_obj_ref_998_resized, req => array_obj_ref_999_index_0_resize_req_0, ack => array_obj_ref_999_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_999_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_998_scaled, dout => array_obj_ref_999_final_offset, req => array_obj_ref_999_offset_inst_req_0, ack => array_obj_ref_999_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1002_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_566, dout => ptr_deref_1002_resized_base_address, req => ptr_deref_1002_base_resize_req_0, ack => ptr_deref_1002_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1016_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => elt5x_xi11_1013, dout => ptr_deref_1016_resized_base_address, req => ptr_deref_1016_base_resize_req_0, ack => ptr_deref_1016_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1030_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp65_1028, dout => ptr_deref_1030_resized_base_address, req => ptr_deref_1030_base_resize_req_0, ack => ptr_deref_1030_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1046_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => elt5x_xi_1043, dout => ptr_deref_1046_resized_base_address, req => ptr_deref_1046_base_resize_req_0, ack => ptr_deref_1046_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1060_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp68_1058, dout => ptr_deref_1060_resized_base_address, req => ptr_deref_1060_base_resize_req_0, ack => ptr_deref_1060_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_553_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp15_550, dout => ptr_deref_553_resized_base_address, req => ptr_deref_553_base_resize_req_0, ack => ptr_deref_553_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_569_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_566, dout => ptr_deref_569_resized_base_address, req => ptr_deref_569_base_resize_req_0, ack => ptr_deref_569_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_616_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp25_613, dout => ptr_deref_616_resized_base_address, req => ptr_deref_616_base_resize_req_0, ack => ptr_deref_616_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_783_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => scevgep12x_xix_xi_780, dout => ptr_deref_783_resized_base_address, req => ptr_deref_783_base_resize_req_0, ack => ptr_deref_783_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_862_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xinx_xlcssax_xix_xi_834, dout => ptr_deref_862_resized_base_address, req => ptr_deref_862_base_resize_req_0, ack => ptr_deref_862_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_939_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp54_937, dout => ptr_deref_939_resized_base_address, req => ptr_deref_939_base_resize_req_0, ack => ptr_deref_939_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_960_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp56_958, dout => ptr_deref_960_resized_base_address, req => ptr_deref_960_base_resize_req_0, ack => ptr_deref_960_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1012_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp63_1009, dout => elt5x_xi11_1013, req => type_cast_1012_inst_req_0, ack => type_cast_1012_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1027_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp64_1024, dout => tmp65_1028, req => type_cast_1027_inst_req_0, ack => type_cast_1027_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1042_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp66_1039, dout => elt5x_xi_1043, req => type_cast_1042_inst_req_0, ack => type_cast_1042_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1057_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp67_1054, dout => tmp68_1058, req => type_cast_1057_inst_req_0, ack => type_cast_1057_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1078_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp14_543, dout => tmp70_1079, req => type_cast_1078_inst_req_0, ack => type_cast_1078_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1082_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp70_1079, dout => type_cast_1082_wire, req => type_cast_1082_inst_req_0, ack => type_cast_1082_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_538_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_537_wire, dout => tmp13_539, req => type_cast_538_inst_req_0, ack => type_cast_538_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_542_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_539, dout => tmp14_543, req => type_cast_542_inst_req_0, ack => type_cast_542_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_573_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp19_570, dout => tmp20_574, req => type_cast_573_inst_req_0, ack => type_cast_573_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_577_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp16_554, dout => tmp21_578, req => type_cast_577_inst_req_0, ack => type_cast_577_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_593_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp23_589, dout => type_cast_593_wire, req => type_cast_593_inst_req_0, ack => type_cast_593_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_612_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_559, dout => tmp25_613, req => type_cast_612_inst_req_0, ack => type_cast_612_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_638_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp34x_xi_635, dout => tmp35x_xi_639, req => type_cast_638_inst_req_0, ack => type_cast_638_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_685_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp32_682, dout => tmp33_686, req => type_cast_685_inst_req_0, ack => type_cast_685_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_740_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnextx_xi14x_xi_807, dout => type_cast_740_wire, req => type_cast_740_inst_req_0, ack => type_cast_740_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_747_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_793, dout => type_cast_747_wire, req => type_cast_747_inst_req_0, ack => type_cast_747_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_779_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => scevgep_775, dout => scevgep12x_xix_xi_780, req => type_cast_779_inst_req_0, ack => type_cast_779_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_787_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp38_784, dout => tmp39_788, req => type_cast_787_inst_req_0, ack => type_cast_787_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_796_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17x_xix_xi_759, dout => type_cast_796_wire, req => type_cast_796_inst_req_0, ack => type_cast_796_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_830_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_793, dout => type_cast_830_wire, req => type_cast_830_inst_req_0, ack => type_cast_830_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_837_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => scevgep14x_xix_xi_824, dout => type_cast_837_wire, req => type_cast_837_inst_req_0, ack => type_cast_837_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_839_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17_559, dout => type_cast_839_wire, req => type_cast_839_inst_req_0, ack => type_cast_839_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_843_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17x_xix_xi_759, dout => type_cast_843_wire, req => type_cast_843_inst_req_0, ack => type_cast_843_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_845_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp30_662, dout => type_cast_845_wire, req => type_cast_845_inst_req_0, ack => type_cast_845_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_866_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 32, flow_through => false ) 
      port map( din => tmp43_863, dout => tmp44_867, req => type_cast_866_inst_req_0, ack => type_cast_866_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_878_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp45_872, dout => type_cast_878_wire, req => type_cast_878_inst_req_0, ack => type_cast_878_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_880_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => xx_xlcssa5x_xix_xi_827, dout => type_cast_880_wire, req => type_cast_880_inst_req_0, ack => type_cast_880_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_912_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp51_909, dout => tmp52_913, req => type_cast_912_inst_req_0, ack => type_cast_912_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_774_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_774_index_0_rename_ack_0 <= array_obj_ref_774_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_773_resized;
      simple_obj_ref_773_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_823_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_823_index_0_rename_ack_0 <= array_obj_ref_823_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_822_resized;
      simple_obj_ref_822_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_950_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_950_index_0_rename_ack_0 <= array_obj_ref_950_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_949_resized;
      simple_obj_ref_949_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_999_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_999_index_0_rename_ack_0 <= array_obj_ref_999_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_998_resized;
      simple_obj_ref_998_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1002_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1002_gather_scatter_ack_0 <= ptr_deref_1002_gather_scatter_req_0;
      aggregated_sig <= tmp62_1000;
      ptr_deref_1002_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1002_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1002_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1002_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1002_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1002_root_address_inst_ack_0 <= ptr_deref_1002_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1002_resized_base_address;
      ptr_deref_1002_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1016_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1016_gather_scatter_ack_0 <= ptr_deref_1016_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1016_data_3 & ptr_deref_1016_data_2 & ptr_deref_1016_data_1 & ptr_deref_1016_data_0;
      val6x_xi12_1017 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1016_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1016_root_address_inst_ack_0 <= ptr_deref_1016_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1016_resized_base_address;
      ptr_deref_1016_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1030_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1030_gather_scatter_ack_0 <= ptr_deref_1030_gather_scatter_req_0;
      aggregated_sig <= val6x_xi12_1017;
      ptr_deref_1030_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1030_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1030_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1030_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1030_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1030_root_address_inst_ack_0 <= ptr_deref_1030_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1030_resized_base_address;
      ptr_deref_1030_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1046_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1046_gather_scatter_ack_0 <= ptr_deref_1046_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1046_data_3 & ptr_deref_1046_data_2 & ptr_deref_1046_data_1 & ptr_deref_1046_data_0;
      val6x_xi_1047 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1046_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1046_root_address_inst_ack_0 <= ptr_deref_1046_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1046_resized_base_address;
      ptr_deref_1046_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1060_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1060_gather_scatter_ack_0 <= ptr_deref_1060_gather_scatter_req_0;
      aggregated_sig <= val6x_xi_1047;
      ptr_deref_1060_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1060_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1060_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1060_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1060_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1060_root_address_inst_ack_0 <= ptr_deref_1060_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1060_resized_base_address;
      ptr_deref_1060_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_553_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_553_gather_scatter_ack_0 <= ptr_deref_553_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_553_data_3 & ptr_deref_553_data_2 & ptr_deref_553_data_1 & ptr_deref_553_data_0;
      tmp16_554 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_553_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_553_root_address_inst_ack_0 <= ptr_deref_553_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_553_resized_base_address;
      ptr_deref_553_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_569_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_569_gather_scatter_ack_0 <= ptr_deref_569_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_569_data_3 & ptr_deref_569_data_2 & ptr_deref_569_data_1 & ptr_deref_569_data_0;
      tmp19_570 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_569_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_569_root_address_inst_ack_0 <= ptr_deref_569_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_569_resized_base_address;
      ptr_deref_569_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_616_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_616_gather_scatter_ack_0 <= ptr_deref_616_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_616_data_3 & ptr_deref_616_data_2 & ptr_deref_616_data_1 & ptr_deref_616_data_0;
      tmp26_617 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_616_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_616_root_address_inst_ack_0 <= ptr_deref_616_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_616_resized_base_address;
      ptr_deref_616_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_783_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_783_gather_scatter_ack_0 <= ptr_deref_783_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_783_data_1 & ptr_deref_783_data_0;
      tmp38_784 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_783_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_783_root_address_inst_ack_0 <= ptr_deref_783_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_783_resized_base_address;
      ptr_deref_783_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_862_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_862_addr_0_ack_0 <= ptr_deref_862_addr_0_req_0;
      aggregated_sig <= ptr_deref_862_root_address;
      ptr_deref_862_word_address_0 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_862_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_862_gather_scatter_ack_0 <= ptr_deref_862_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_862_data_0;
      tmp43_863 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_862_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_862_root_address_inst_ack_0 <= ptr_deref_862_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_862_resized_base_address;
      ptr_deref_862_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_939_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_939_gather_scatter_ack_0 <= ptr_deref_939_gather_scatter_req_0;
      aggregated_sig <= tmp17_559;
      ptr_deref_939_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_939_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_939_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_939_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_939_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_939_root_address_inst_ack_0 <= ptr_deref_939_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_939_resized_base_address;
      ptr_deref_939_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_960_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_960_gather_scatter_ack_0 <= ptr_deref_960_gather_scatter_req_0;
      aggregated_sig <= tmp55_951;
      ptr_deref_960_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_960_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_960_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_960_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_960_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_960_root_address_inst_ack_0 <= ptr_deref_960_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_960_resized_base_address;
      ptr_deref_960_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_1069_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp69_1068;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1069_branch_req_0,
          ack0 => if_stmt_1069_branch_ack_0,
          ack1 => if_stmt_1069_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_599_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp24_598;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_599_branch_req_0,
          ack0 => if_stmt_599_branch_ack_0,
          ack1 => if_stmt_599_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_640_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp28_629;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_640_branch_req_0,
          ack0 => if_stmt_640_branch_ack_0,
          ack1 => if_stmt_640_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_669_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp31_668;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_669_branch_req_0,
          ack0 => if_stmt_669_branch_ack_0,
          ack1 => if_stmt_669_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_702_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xi_701;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_702_branch_req_0,
          ack0 => if_stmt_702_branch_ack_0,
          ack1 => if_stmt_702_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_719_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp36_718;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_719_branch_req_0,
          ack0 => if_stmt_719_branch_ack_0,
          ack1 => if_stmt_719_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_808_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp41_801;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_808_branch_req_0,
          ack0 => if_stmt_808_branch_ack_0,
          ack1 => if_stmt_808_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_853_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp42_852;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_853_branch_req_0,
          ack0 => if_stmt_853_branch_ack_0,
          ack1 => if_stmt_853_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_920_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp53_919;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_920_branch_req_0,
          ack0 => if_stmt_920_branch_ack_0,
          ack1 => if_stmt_920_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_968_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp57_967;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_968_branch_req_0,
          ack0 => if_stmt_968_branch_ack_0,
          ack1 => if_stmt_968_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1008_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1008_resized_base_address;
      array_obj_ref_1008_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1008_root_address_inst_req_0,
          ackL => array_obj_ref_1008_root_address_inst_ack_0,
          reqR => array_obj_ref_1008_root_address_inst_req_1,
          ackR => array_obj_ref_1008_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1023_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1023_resized_base_address;
      array_obj_ref_1023_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1023_root_address_inst_req_0,
          ackL => array_obj_ref_1023_root_address_inst_ack_0,
          reqR => array_obj_ref_1023_root_address_inst_req_1,
          ackR => array_obj_ref_1023_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1038_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1038_resized_base_address;
      array_obj_ref_1038_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1038_root_address_inst_req_0,
          ackL => array_obj_ref_1038_root_address_inst_ack_0,
          reqR => array_obj_ref_1038_root_address_inst_req_1,
          ackR => array_obj_ref_1038_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1053_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1053_resized_base_address;
      array_obj_ref_1053_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1053_root_address_inst_req_0,
          ackL => array_obj_ref_1053_root_address_inst_ack_0,
          reqR => array_obj_ref_1053_root_address_inst_req_1,
          ackR => array_obj_ref_1053_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_549_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_549_resized_base_address;
      array_obj_ref_549_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_549_root_address_inst_req_0,
          ackL => array_obj_ref_549_root_address_inst_ack_0,
          reqR => array_obj_ref_549_root_address_inst_req_1,
          ackR => array_obj_ref_549_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_558_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_558_resized_base_address;
      array_obj_ref_558_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_558_root_address_inst_req_0,
          ackL => array_obj_ref_558_root_address_inst_ack_0,
          reqR => array_obj_ref_558_root_address_inst_req_1,
          ackR => array_obj_ref_558_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_565_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_565_resized_base_address;
      array_obj_ref_565_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_565_root_address_inst_req_0,
          ackL => array_obj_ref_565_root_address_inst_ack_0,
          reqR => array_obj_ref_565_root_address_inst_req_1,
          ackR => array_obj_ref_565_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_774_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_774_final_offset & array_obj_ref_774_resized_base_address;
      array_obj_ref_774_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_774_root_address_inst_req_0,
          ackL => array_obj_ref_774_root_address_inst_ack_0,
          reqR => array_obj_ref_774_root_address_inst_req_1,
          ackR => array_obj_ref_774_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_823_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_823_final_offset & array_obj_ref_823_resized_base_address;
      array_obj_ref_823_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_823_root_address_inst_req_0,
          ackL => array_obj_ref_823_root_address_inst_ack_0,
          reqR => array_obj_ref_823_root_address_inst_req_1,
          ackR => array_obj_ref_823_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_936_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_936_resized_base_address;
      array_obj_ref_936_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_936_root_address_inst_req_0,
          ackL => array_obj_ref_936_root_address_inst_ack_0,
          reqR => array_obj_ref_936_root_address_inst_req_1,
          ackR => array_obj_ref_936_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_950_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_950_final_offset & array_obj_ref_950_resized_base_address;
      array_obj_ref_950_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_950_root_address_inst_req_0,
          ackL => array_obj_ref_950_root_address_inst_ack_0,
          reqR => array_obj_ref_950_root_address_inst_req_1,
          ackR => array_obj_ref_950_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_957_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_957_resized_base_address;
      array_obj_ref_957_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001010100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_957_root_address_inst_req_0,
          ackL => array_obj_ref_957_root_address_inst_ack_0,
          reqR => array_obj_ref_957_root_address_inst_req_1,
          ackR => array_obj_ref_957_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_999_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_999_final_offset & array_obj_ref_999_resized_base_address;
      array_obj_ref_999_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_999_root_address_inst_req_0,
          ackL => array_obj_ref_999_root_address_inst_ack_0,
          reqR => array_obj_ref_999_root_address_inst_req_1,
          ackR => array_obj_ref_999_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_1067_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp14_543;
      tmp69_1068 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1067_inst_req_0,
          ackL => binary_1067_inst_ack_0,
          reqR => binary_1067_inst_req_1,
          ackR => binary_1067_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_582_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_574 & tmp21_578;
      tmp22_583 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_582_inst_req_0,
          ackL => binary_582_inst_ack_0,
          reqR => binary_582_inst_req_1,
          ackR => binary_582_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_588_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp22_583;
      tmp23_589 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111110010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_588_inst_req_0,
          ackL => binary_588_inst_ack_0,
          reqR => binary_588_inst_req_1,
          ackR => binary_588_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_597_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_593_wire;
      tmp24_598 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_597_inst_req_0,
          ackL => binary_597_inst_ack_0,
          reqR => binary_597_inst_req_1,
          ackR => binary_597_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_622_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_617;
      tmp27_623 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011110000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_622_inst_req_0,
          ackL => binary_622_inst_ack_0,
          reqR => binary_622_inst_req_1,
          ackR => binary_622_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_628_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp27_623;
      tmp28_629 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_628_inst_req_0,
          ackL => binary_628_inst_ack_0,
          reqR => binary_628_inst_req_1,
          ackR => binary_628_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_634_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_617;
      tmp34x_xi_635 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_634_inst_req_0,
          ackL => binary_634_inst_ack_0,
          reqR => binary_634_inst_req_1,
          ackR => binary_634_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_655_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_617;
      tmp29_656 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_655_inst_req_0,
          ackL => binary_655_inst_ack_0,
          reqR => binary_655_inst_req_1,
          ackR => binary_655_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_661_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp29_656;
      tmp30_662 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000111100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_661_inst_req_0,
          ackL => binary_661_inst_ack_0,
          reqR => binary_661_inst_req_1,
          ackR => binary_661_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_667_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_662;
      tmp31_668 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_667_inst_req_0,
          ackL => binary_667_inst_ack_0,
          reqR => binary_667_inst_req_1,
          ackR => binary_667_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_690_inst binary_966_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp33_686 & tmp23_589 & tmp23_589 & tmp33_686;
      tmp34_691 <= data_out(1 downto 1);
      tmp57_967 <= data_out(0 downto 0);
      reqL(1) <= binary_690_inst_req_0;
      reqL(0) <= binary_966_inst_req_0;
      binary_690_inst_ack_0 <= ackL(1);
      binary_966_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_690_inst_req_1;
      reqR(0) <= binary_966_inst_req_1;
      binary_690_inst_ack_1 <= ackR(1);
      binary_966_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_695_inst binary_983_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp33_686 & tmp30_662 & tmp22_583 & tmp58_979;
      tmp35_696 <= data_out(1 downto 1);
      tmp59_984 <= data_out(0 downto 0);
      reqL(1) <= binary_695_inst_req_0;
      reqL(0) <= binary_983_inst_req_0;
      binary_695_inst_ack_0 <= ackL(1);
      binary_983_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_695_inst_req_1;
      reqR(0) <= binary_983_inst_req_1;
      binary_695_inst_ack_1 <= ackR(1);
      binary_983_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_700_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp34_691 & tmp35_696;
      orx_xcondx_xi_701 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_700_inst_req_0,
          ackL => binary_700_inst_ack_0,
          reqR => binary_700_inst_req_1,
          ackR => binary_700_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_717_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_662;
      tmp36_718 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_717_inst_req_0,
          ackL => binary_717_inst_ack_0,
          reqR => binary_717_inst_req_1,
          ackR => binary_717_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_730_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_662;
      tmp5_731 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_730_inst_req_0,
          ackL => binary_730_inst_ack_0,
          reqR => binary_730_inst_req_1,
          ackR => binary_730_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_753_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_734;
      tmp_754 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_753_inst_req_0,
          ackL => binary_753_inst_ack_0,
          reqR => binary_753_inst_req_1,
          ackR => binary_753_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_758_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp5_731 & tmp_754;
      tmp17x_xix_xi_759 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_758_inst_req_0,
          ackL => binary_758_inst_ack_0,
          reqR => binary_758_inst_req_1,
          ackR => binary_758_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_764_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_734;
      tmpx_xix_xi_765 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_764_inst_req_0,
          ackL => binary_764_inst_ack_0,
          reqR => binary_764_inst_req_1,
          ackR => binary_764_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_770_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xix_xi_765;
      tmp8_771 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_770_inst_req_0,
          ackL => binary_770_inst_ack_0,
          reqR => binary_770_inst_req_1,
          ackR => binary_770_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_792_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp39_788 & tmp37_741;
      tmp40_793 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_792_inst_req_0,
          ackL => binary_792_inst_ack_0,
          reqR => binary_792_inst_req_1,
          ackR => binary_792_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_800_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_796_wire;
      tmp41_801 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_800_inst_req_0,
          ackL => binary_800_inst_ack_0,
          reqR => binary_800_inst_req_1,
          ackR => binary_800_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_806_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_734;
      indvarx_xnextx_xi14x_xi_807 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_806_inst_req_0,
          ackL => binary_806_inst_ack_0,
          reqR => binary_806_inst_req_1,
          ackR => binary_806_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_819_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xix_xi_765;
      xx_xsum20x_xi_820 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_819_inst_req_0,
          ackL => binary_819_inst_ack_0,
          reqR => binary_819_inst_req_1,
          ackR => binary_819_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_851_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xlcssax_xix_xi_840;
      tmp42_852 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_851_inst_req_0,
          ackL => binary_851_inst_ack_0,
          reqR => binary_851_inst_req_1,
          ackR => binary_851_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_871_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp44_867 & xx_xlcssa5x_xix_xi_827;
      tmp45_872 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_871_inst_req_0,
          ackL => binary_871_inst_ack_0,
          reqR => binary_871_inst_req_1,
          ackR => binary_871_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_886_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp46_875;
      tmp47_887 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_886_inst_req_0,
          ackL => binary_886_inst_ack_0,
          reqR => binary_886_inst_req_1,
          ackR => binary_886_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_892_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp46_875;
      tmp48_893 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_892_inst_req_0,
          ackL => binary_892_inst_ack_0,
          reqR => binary_892_inst_req_1,
          ackR => binary_892_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_897_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp47_887 & tmp48_893;
      tmp49_898 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_897_inst_req_0,
          ackL => binary_897_inst_ack_0,
          reqR => binary_897_inst_req_1,
          ackR => binary_897_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_903_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp49_898;
      tmp50_904 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_903_inst_req_0,
          ackL => binary_903_inst_ack_0,
          reqR => binary_903_inst_req_1,
          ackR => binary_903_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_908_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp50_904 & tmp49_898;
      tmp51_909 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_908_inst_req_0,
          ackL => binary_908_inst_ack_0,
          reqR => binary_908_inst_req_1,
          ackR => binary_908_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_918_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp52_913;
      tmp53_919 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1111111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_918_inst_req_0,
          ackL => binary_918_inst_ack_0,
          reqR => binary_918_inst_req_1,
          ackR => binary_918_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_946_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_662;
      xx_xsumx_xi_947 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_946_inst_req_0,
          ackL => binary_946_inst_ack_0,
          reqR => binary_946_inst_req_1,
          ackR => binary_946_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_978_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp23_589 & tmp33_686;
      tmp58_979 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_978_inst_req_0,
          ackL => binary_978_inst_ack_0,
          reqR => binary_978_inst_req_1,
          ackR => binary_978_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_995_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_993_wire_constant & tmp60_990;
      tmp61_996 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_995_inst_req_0,
          ackL => binary_995_inst_ack_0,
          reqR => binary_995_inst_req_1,
          ackR => binary_995_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : ptr_deref_1002_addr_0 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1002_root_address;
      ptr_deref_1002_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1002_addr_0_req_0,
          ackL => ptr_deref_1002_addr_0_ack_0,
          reqR => ptr_deref_1002_addr_0_req_1,
          ackR => ptr_deref_1002_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : ptr_deref_1002_addr_1 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1002_root_address;
      ptr_deref_1002_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1002_addr_1_req_0,
          ackL => ptr_deref_1002_addr_1_ack_0,
          reqR => ptr_deref_1002_addr_1_req_1,
          ackR => ptr_deref_1002_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : ptr_deref_1002_addr_2 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1002_root_address;
      ptr_deref_1002_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1002_addr_2_req_0,
          ackL => ptr_deref_1002_addr_2_ack_0,
          reqR => ptr_deref_1002_addr_2_req_1,
          ackR => ptr_deref_1002_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : ptr_deref_1002_addr_3 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1002_root_address;
      ptr_deref_1002_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1002_addr_3_req_0,
          ackL => ptr_deref_1002_addr_3_ack_0,
          reqR => ptr_deref_1002_addr_3_req_1,
          ackR => ptr_deref_1002_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : ptr_deref_1016_addr_0 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1016_root_address;
      ptr_deref_1016_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1016_addr_0_req_0,
          ackL => ptr_deref_1016_addr_0_ack_0,
          reqR => ptr_deref_1016_addr_0_req_1,
          ackR => ptr_deref_1016_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_1016_addr_1 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1016_root_address;
      ptr_deref_1016_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1016_addr_1_req_0,
          ackL => ptr_deref_1016_addr_1_ack_0,
          reqR => ptr_deref_1016_addr_1_req_1,
          ackR => ptr_deref_1016_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_1016_addr_2 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1016_root_address;
      ptr_deref_1016_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1016_addr_2_req_0,
          ackL => ptr_deref_1016_addr_2_ack_0,
          reqR => ptr_deref_1016_addr_2_req_1,
          ackR => ptr_deref_1016_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_1016_addr_3 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1016_root_address;
      ptr_deref_1016_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1016_addr_3_req_0,
          ackL => ptr_deref_1016_addr_3_ack_0,
          reqR => ptr_deref_1016_addr_3_req_1,
          ackR => ptr_deref_1016_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_1030_addr_0 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1030_root_address;
      ptr_deref_1030_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1030_addr_0_req_0,
          ackL => ptr_deref_1030_addr_0_ack_0,
          reqR => ptr_deref_1030_addr_0_req_1,
          ackR => ptr_deref_1030_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_1030_addr_1 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1030_root_address;
      ptr_deref_1030_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1030_addr_1_req_0,
          ackL => ptr_deref_1030_addr_1_ack_0,
          reqR => ptr_deref_1030_addr_1_req_1,
          ackR => ptr_deref_1030_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_1030_addr_2 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1030_root_address;
      ptr_deref_1030_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1030_addr_2_req_0,
          ackL => ptr_deref_1030_addr_2_ack_0,
          reqR => ptr_deref_1030_addr_2_req_1,
          ackR => ptr_deref_1030_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_1030_addr_3 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1030_root_address;
      ptr_deref_1030_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1030_addr_3_req_0,
          ackL => ptr_deref_1030_addr_3_ack_0,
          reqR => ptr_deref_1030_addr_3_req_1,
          ackR => ptr_deref_1030_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : ptr_deref_1046_addr_0 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1046_root_address;
      ptr_deref_1046_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1046_addr_0_req_0,
          ackL => ptr_deref_1046_addr_0_ack_0,
          reqR => ptr_deref_1046_addr_0_req_1,
          ackR => ptr_deref_1046_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : ptr_deref_1046_addr_1 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1046_root_address;
      ptr_deref_1046_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1046_addr_1_req_0,
          ackL => ptr_deref_1046_addr_1_ack_0,
          reqR => ptr_deref_1046_addr_1_req_1,
          ackR => ptr_deref_1046_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : ptr_deref_1046_addr_2 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1046_root_address;
      ptr_deref_1046_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1046_addr_2_req_0,
          ackL => ptr_deref_1046_addr_2_ack_0,
          reqR => ptr_deref_1046_addr_2_req_1,
          ackR => ptr_deref_1046_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : ptr_deref_1046_addr_3 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1046_root_address;
      ptr_deref_1046_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1046_addr_3_req_0,
          ackL => ptr_deref_1046_addr_3_ack_0,
          reqR => ptr_deref_1046_addr_3_req_1,
          ackR => ptr_deref_1046_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : ptr_deref_1060_addr_0 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1060_root_address;
      ptr_deref_1060_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1060_addr_0_req_0,
          ackL => ptr_deref_1060_addr_0_ack_0,
          reqR => ptr_deref_1060_addr_0_req_1,
          ackR => ptr_deref_1060_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : ptr_deref_1060_addr_1 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1060_root_address;
      ptr_deref_1060_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1060_addr_1_req_0,
          ackL => ptr_deref_1060_addr_1_ack_0,
          reqR => ptr_deref_1060_addr_1_req_1,
          ackR => ptr_deref_1060_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : ptr_deref_1060_addr_2 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1060_root_address;
      ptr_deref_1060_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1060_addr_2_req_0,
          ackL => ptr_deref_1060_addr_2_ack_0,
          reqR => ptr_deref_1060_addr_2_req_1,
          ackR => ptr_deref_1060_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : ptr_deref_1060_addr_3 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1060_root_address;
      ptr_deref_1060_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1060_addr_3_req_0,
          ackL => ptr_deref_1060_addr_3_ack_0,
          reqR => ptr_deref_1060_addr_3_req_1,
          ackR => ptr_deref_1060_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : ptr_deref_553_addr_0 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_0_req_0,
          ackL => ptr_deref_553_addr_0_ack_0,
          reqR => ptr_deref_553_addr_0_req_1,
          ackR => ptr_deref_553_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : ptr_deref_553_addr_1 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_1_req_0,
          ackL => ptr_deref_553_addr_1_ack_0,
          reqR => ptr_deref_553_addr_1_req_1,
          ackR => ptr_deref_553_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : ptr_deref_553_addr_2 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_2_req_0,
          ackL => ptr_deref_553_addr_2_ack_0,
          reqR => ptr_deref_553_addr_2_req_1,
          ackR => ptr_deref_553_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : ptr_deref_553_addr_3 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_3_req_0,
          ackL => ptr_deref_553_addr_3_ack_0,
          reqR => ptr_deref_553_addr_3_req_1,
          ackR => ptr_deref_553_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : ptr_deref_569_addr_0 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_0_req_0,
          ackL => ptr_deref_569_addr_0_ack_0,
          reqR => ptr_deref_569_addr_0_req_1,
          ackR => ptr_deref_569_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : ptr_deref_569_addr_1 
    SplitOperatorGroup72: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_1_req_0,
          ackL => ptr_deref_569_addr_1_ack_0,
          reqR => ptr_deref_569_addr_1_req_1,
          ackR => ptr_deref_569_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : ptr_deref_569_addr_2 
    SplitOperatorGroup73: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_2_req_0,
          ackL => ptr_deref_569_addr_2_ack_0,
          reqR => ptr_deref_569_addr_2_req_1,
          ackR => ptr_deref_569_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : ptr_deref_569_addr_3 
    SplitOperatorGroup74: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_3_req_0,
          ackL => ptr_deref_569_addr_3_ack_0,
          reqR => ptr_deref_569_addr_3_req_1,
          ackR => ptr_deref_569_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : ptr_deref_616_addr_0 
    SplitOperatorGroup75: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_616_root_address;
      ptr_deref_616_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_616_addr_0_req_0,
          ackL => ptr_deref_616_addr_0_ack_0,
          reqR => ptr_deref_616_addr_0_req_1,
          ackR => ptr_deref_616_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : ptr_deref_616_addr_1 
    SplitOperatorGroup76: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_616_root_address;
      ptr_deref_616_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_616_addr_1_req_0,
          ackL => ptr_deref_616_addr_1_ack_0,
          reqR => ptr_deref_616_addr_1_req_1,
          ackR => ptr_deref_616_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : ptr_deref_616_addr_2 
    SplitOperatorGroup77: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_616_root_address;
      ptr_deref_616_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_616_addr_2_req_0,
          ackL => ptr_deref_616_addr_2_ack_0,
          reqR => ptr_deref_616_addr_2_req_1,
          ackR => ptr_deref_616_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared split operator group (78) : ptr_deref_616_addr_3 
    SplitOperatorGroup78: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_616_root_address;
      ptr_deref_616_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_616_addr_3_req_0,
          ackL => ptr_deref_616_addr_3_ack_0,
          reqR => ptr_deref_616_addr_3_req_1,
          ackR => ptr_deref_616_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 78
    -- shared split operator group (79) : ptr_deref_783_addr_0 
    SplitOperatorGroup79: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_783_root_address;
      ptr_deref_783_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_783_addr_0_req_0,
          ackL => ptr_deref_783_addr_0_ack_0,
          reqR => ptr_deref_783_addr_0_req_1,
          ackR => ptr_deref_783_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 79
    -- shared split operator group (80) : ptr_deref_783_addr_1 
    SplitOperatorGroup80: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_783_root_address;
      ptr_deref_783_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_783_addr_1_req_0,
          ackL => ptr_deref_783_addr_1_ack_0,
          reqR => ptr_deref_783_addr_1_req_1,
          ackR => ptr_deref_783_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : ptr_deref_939_addr_0 
    SplitOperatorGroup81: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_939_root_address;
      ptr_deref_939_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_939_addr_0_req_0,
          ackL => ptr_deref_939_addr_0_ack_0,
          reqR => ptr_deref_939_addr_0_req_1,
          ackR => ptr_deref_939_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- shared split operator group (82) : ptr_deref_939_addr_1 
    SplitOperatorGroup82: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_939_root_address;
      ptr_deref_939_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_939_addr_1_req_0,
          ackL => ptr_deref_939_addr_1_ack_0,
          reqR => ptr_deref_939_addr_1_req_1,
          ackR => ptr_deref_939_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- shared split operator group (83) : ptr_deref_939_addr_2 
    SplitOperatorGroup83: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_939_root_address;
      ptr_deref_939_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_939_addr_2_req_0,
          ackL => ptr_deref_939_addr_2_ack_0,
          reqR => ptr_deref_939_addr_2_req_1,
          ackR => ptr_deref_939_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- shared split operator group (84) : ptr_deref_939_addr_3 
    SplitOperatorGroup84: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_939_root_address;
      ptr_deref_939_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_939_addr_3_req_0,
          ackL => ptr_deref_939_addr_3_ack_0,
          reqR => ptr_deref_939_addr_3_req_1,
          ackR => ptr_deref_939_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared split operator group (85) : ptr_deref_960_addr_0 
    SplitOperatorGroup85: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_960_root_address;
      ptr_deref_960_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_960_addr_0_req_0,
          ackL => ptr_deref_960_addr_0_ack_0,
          reqR => ptr_deref_960_addr_0_req_1,
          ackR => ptr_deref_960_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- shared split operator group (86) : ptr_deref_960_addr_1 
    SplitOperatorGroup86: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_960_root_address;
      ptr_deref_960_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_960_addr_1_req_0,
          ackL => ptr_deref_960_addr_1_ack_0,
          reqR => ptr_deref_960_addr_1_req_1,
          ackR => ptr_deref_960_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 86
    -- shared split operator group (87) : ptr_deref_960_addr_2 
    SplitOperatorGroup87: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_960_root_address;
      ptr_deref_960_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_960_addr_2_req_0,
          ackL => ptr_deref_960_addr_2_ack_0,
          reqR => ptr_deref_960_addr_2_req_1,
          ackR => ptr_deref_960_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 87
    -- shared split operator group (88) : ptr_deref_960_addr_3 
    SplitOperatorGroup88: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_960_root_address;
      ptr_deref_960_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_960_addr_3_req_0,
          ackL => ptr_deref_960_addr_3_ack_0,
          reqR => ptr_deref_960_addr_3_req_1,
          ackR => ptr_deref_960_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 88
    -- shared load operator group (0) : ptr_deref_553_load_3 ptr_deref_553_load_0 ptr_deref_616_load_2 ptr_deref_553_load_1 ptr_deref_616_load_3 ptr_deref_569_load_0 ptr_deref_553_load_2 ptr_deref_569_load_1 ptr_deref_569_load_2 ptr_deref_569_load_3 ptr_deref_783_load_0 ptr_deref_783_load_1 ptr_deref_616_load_1 ptr_deref_616_load_0 ptr_deref_862_load_0 ptr_deref_1016_load_0 ptr_deref_1016_load_1 ptr_deref_1016_load_2 ptr_deref_1016_load_3 ptr_deref_1046_load_0 ptr_deref_1046_load_1 ptr_deref_1046_load_2 ptr_deref_1046_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(367 downto 0);
      signal data_out: std_logic_vector(183 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 22 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_553_load_3_req_0,
        ptr_deref_553_load_3_ack_0,
        ptr_deref_553_load_3_req_1,
        ptr_deref_553_load_3_ack_1,
        "ptr_deref_553_load_3",
        "memory_space_5" ,
        ptr_deref_553_data_3,
        ptr_deref_553_word_address_3,
        "ptr_deref_553_data_3",
        "ptr_deref_553_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_0_req_0,
        ptr_deref_553_load_0_ack_0,
        ptr_deref_553_load_0_req_1,
        ptr_deref_553_load_0_ack_1,
        "ptr_deref_553_load_0",
        "memory_space_5" ,
        ptr_deref_553_data_0,
        ptr_deref_553_word_address_0,
        "ptr_deref_553_data_0",
        "ptr_deref_553_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_616_load_2_req_0,
        ptr_deref_616_load_2_ack_0,
        ptr_deref_616_load_2_req_1,
        ptr_deref_616_load_2_ack_1,
        "ptr_deref_616_load_2",
        "memory_space_5" ,
        ptr_deref_616_data_2,
        ptr_deref_616_word_address_2,
        "ptr_deref_616_data_2",
        "ptr_deref_616_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_1_req_0,
        ptr_deref_553_load_1_ack_0,
        ptr_deref_553_load_1_req_1,
        ptr_deref_553_load_1_ack_1,
        "ptr_deref_553_load_1",
        "memory_space_5" ,
        ptr_deref_553_data_1,
        ptr_deref_553_word_address_1,
        "ptr_deref_553_data_1",
        "ptr_deref_553_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_616_load_3_req_0,
        ptr_deref_616_load_3_ack_0,
        ptr_deref_616_load_3_req_1,
        ptr_deref_616_load_3_ack_1,
        "ptr_deref_616_load_3",
        "memory_space_5" ,
        ptr_deref_616_data_3,
        ptr_deref_616_word_address_3,
        "ptr_deref_616_data_3",
        "ptr_deref_616_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_0_req_0,
        ptr_deref_569_load_0_ack_0,
        ptr_deref_569_load_0_req_1,
        ptr_deref_569_load_0_ack_1,
        "ptr_deref_569_load_0",
        "memory_space_5" ,
        ptr_deref_569_data_0,
        ptr_deref_569_word_address_0,
        "ptr_deref_569_data_0",
        "ptr_deref_569_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_2_req_0,
        ptr_deref_553_load_2_ack_0,
        ptr_deref_553_load_2_req_1,
        ptr_deref_553_load_2_ack_1,
        "ptr_deref_553_load_2",
        "memory_space_5" ,
        ptr_deref_553_data_2,
        ptr_deref_553_word_address_2,
        "ptr_deref_553_data_2",
        "ptr_deref_553_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_1_req_0,
        ptr_deref_569_load_1_ack_0,
        ptr_deref_569_load_1_req_1,
        ptr_deref_569_load_1_ack_1,
        "ptr_deref_569_load_1",
        "memory_space_5" ,
        ptr_deref_569_data_1,
        ptr_deref_569_word_address_1,
        "ptr_deref_569_data_1",
        "ptr_deref_569_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_2_req_0,
        ptr_deref_569_load_2_ack_0,
        ptr_deref_569_load_2_req_1,
        ptr_deref_569_load_2_ack_1,
        "ptr_deref_569_load_2",
        "memory_space_5" ,
        ptr_deref_569_data_2,
        ptr_deref_569_word_address_2,
        "ptr_deref_569_data_2",
        "ptr_deref_569_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_3_req_0,
        ptr_deref_569_load_3_ack_0,
        ptr_deref_569_load_3_req_1,
        ptr_deref_569_load_3_ack_1,
        "ptr_deref_569_load_3",
        "memory_space_5" ,
        ptr_deref_569_data_3,
        ptr_deref_569_word_address_3,
        "ptr_deref_569_data_3",
        "ptr_deref_569_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_783_load_0_req_0,
        ptr_deref_783_load_0_ack_0,
        ptr_deref_783_load_0_req_1,
        ptr_deref_783_load_0_ack_1,
        "ptr_deref_783_load_0",
        "memory_space_5" ,
        ptr_deref_783_data_0,
        ptr_deref_783_word_address_0,
        "ptr_deref_783_data_0",
        "ptr_deref_783_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_783_load_1_req_0,
        ptr_deref_783_load_1_ack_0,
        ptr_deref_783_load_1_req_1,
        ptr_deref_783_load_1_ack_1,
        "ptr_deref_783_load_1",
        "memory_space_5" ,
        ptr_deref_783_data_1,
        ptr_deref_783_word_address_1,
        "ptr_deref_783_data_1",
        "ptr_deref_783_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_616_load_1_req_0,
        ptr_deref_616_load_1_ack_0,
        ptr_deref_616_load_1_req_1,
        ptr_deref_616_load_1_ack_1,
        "ptr_deref_616_load_1",
        "memory_space_5" ,
        ptr_deref_616_data_1,
        ptr_deref_616_word_address_1,
        "ptr_deref_616_data_1",
        "ptr_deref_616_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_616_load_0_req_0,
        ptr_deref_616_load_0_ack_0,
        ptr_deref_616_load_0_req_1,
        ptr_deref_616_load_0_ack_1,
        "ptr_deref_616_load_0",
        "memory_space_5" ,
        ptr_deref_616_data_0,
        ptr_deref_616_word_address_0,
        "ptr_deref_616_data_0",
        "ptr_deref_616_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_862_load_0_req_0,
        ptr_deref_862_load_0_ack_0,
        ptr_deref_862_load_0_req_1,
        ptr_deref_862_load_0_ack_1,
        "ptr_deref_862_load_0",
        "memory_space_5" ,
        ptr_deref_862_data_0,
        ptr_deref_862_word_address_0,
        "ptr_deref_862_data_0",
        "ptr_deref_862_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1016_load_0_req_0,
        ptr_deref_1016_load_0_ack_0,
        ptr_deref_1016_load_0_req_1,
        ptr_deref_1016_load_0_ack_1,
        "ptr_deref_1016_load_0",
        "memory_space_5" ,
        ptr_deref_1016_data_0,
        ptr_deref_1016_word_address_0,
        "ptr_deref_1016_data_0",
        "ptr_deref_1016_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1016_load_1_req_0,
        ptr_deref_1016_load_1_ack_0,
        ptr_deref_1016_load_1_req_1,
        ptr_deref_1016_load_1_ack_1,
        "ptr_deref_1016_load_1",
        "memory_space_5" ,
        ptr_deref_1016_data_1,
        ptr_deref_1016_word_address_1,
        "ptr_deref_1016_data_1",
        "ptr_deref_1016_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1016_load_2_req_0,
        ptr_deref_1016_load_2_ack_0,
        ptr_deref_1016_load_2_req_1,
        ptr_deref_1016_load_2_ack_1,
        "ptr_deref_1016_load_2",
        "memory_space_5" ,
        ptr_deref_1016_data_2,
        ptr_deref_1016_word_address_2,
        "ptr_deref_1016_data_2",
        "ptr_deref_1016_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1016_load_3_req_0,
        ptr_deref_1016_load_3_ack_0,
        ptr_deref_1016_load_3_req_1,
        ptr_deref_1016_load_3_ack_1,
        "ptr_deref_1016_load_3",
        "memory_space_5" ,
        ptr_deref_1016_data_3,
        ptr_deref_1016_word_address_3,
        "ptr_deref_1016_data_3",
        "ptr_deref_1016_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1046_load_0_req_0,
        ptr_deref_1046_load_0_ack_0,
        ptr_deref_1046_load_0_req_1,
        ptr_deref_1046_load_0_ack_1,
        "ptr_deref_1046_load_0",
        "memory_space_5" ,
        ptr_deref_1046_data_0,
        ptr_deref_1046_word_address_0,
        "ptr_deref_1046_data_0",
        "ptr_deref_1046_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1046_load_1_req_0,
        ptr_deref_1046_load_1_ack_0,
        ptr_deref_1046_load_1_req_1,
        ptr_deref_1046_load_1_ack_1,
        "ptr_deref_1046_load_1",
        "memory_space_5" ,
        ptr_deref_1046_data_1,
        ptr_deref_1046_word_address_1,
        "ptr_deref_1046_data_1",
        "ptr_deref_1046_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1046_load_2_req_0,
        ptr_deref_1046_load_2_ack_0,
        ptr_deref_1046_load_2_req_1,
        ptr_deref_1046_load_2_ack_1,
        "ptr_deref_1046_load_2",
        "memory_space_5" ,
        ptr_deref_1046_data_2,
        ptr_deref_1046_word_address_2,
        "ptr_deref_1046_data_2",
        "ptr_deref_1046_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1046_load_3_req_0,
        ptr_deref_1046_load_3_ack_0,
        ptr_deref_1046_load_3_req_1,
        ptr_deref_1046_load_3_ack_1,
        "ptr_deref_1046_load_3",
        "memory_space_5" ,
        ptr_deref_1046_data_3,
        ptr_deref_1046_word_address_3,
        "ptr_deref_1046_data_3",
        "ptr_deref_1046_word_address_3" -- 
      );
      reqL(22) <= ptr_deref_553_load_3_req_0;
      reqL(21) <= ptr_deref_553_load_0_req_0;
      reqL(20) <= ptr_deref_616_load_2_req_0;
      reqL(19) <= ptr_deref_553_load_1_req_0;
      reqL(18) <= ptr_deref_616_load_3_req_0;
      reqL(17) <= ptr_deref_569_load_0_req_0;
      reqL(16) <= ptr_deref_553_load_2_req_0;
      reqL(15) <= ptr_deref_569_load_1_req_0;
      reqL(14) <= ptr_deref_569_load_2_req_0;
      reqL(13) <= ptr_deref_569_load_3_req_0;
      reqL(12) <= ptr_deref_783_load_0_req_0;
      reqL(11) <= ptr_deref_783_load_1_req_0;
      reqL(10) <= ptr_deref_616_load_1_req_0;
      reqL(9) <= ptr_deref_616_load_0_req_0;
      reqL(8) <= ptr_deref_862_load_0_req_0;
      reqL(7) <= ptr_deref_1016_load_0_req_0;
      reqL(6) <= ptr_deref_1016_load_1_req_0;
      reqL(5) <= ptr_deref_1016_load_2_req_0;
      reqL(4) <= ptr_deref_1016_load_3_req_0;
      reqL(3) <= ptr_deref_1046_load_0_req_0;
      reqL(2) <= ptr_deref_1046_load_1_req_0;
      reqL(1) <= ptr_deref_1046_load_2_req_0;
      reqL(0) <= ptr_deref_1046_load_3_req_0;
      ptr_deref_553_load_3_ack_0 <= ackL(22);
      ptr_deref_553_load_0_ack_0 <= ackL(21);
      ptr_deref_616_load_2_ack_0 <= ackL(20);
      ptr_deref_553_load_1_ack_0 <= ackL(19);
      ptr_deref_616_load_3_ack_0 <= ackL(18);
      ptr_deref_569_load_0_ack_0 <= ackL(17);
      ptr_deref_553_load_2_ack_0 <= ackL(16);
      ptr_deref_569_load_1_ack_0 <= ackL(15);
      ptr_deref_569_load_2_ack_0 <= ackL(14);
      ptr_deref_569_load_3_ack_0 <= ackL(13);
      ptr_deref_783_load_0_ack_0 <= ackL(12);
      ptr_deref_783_load_1_ack_0 <= ackL(11);
      ptr_deref_616_load_1_ack_0 <= ackL(10);
      ptr_deref_616_load_0_ack_0 <= ackL(9);
      ptr_deref_862_load_0_ack_0 <= ackL(8);
      ptr_deref_1016_load_0_ack_0 <= ackL(7);
      ptr_deref_1016_load_1_ack_0 <= ackL(6);
      ptr_deref_1016_load_2_ack_0 <= ackL(5);
      ptr_deref_1016_load_3_ack_0 <= ackL(4);
      ptr_deref_1046_load_0_ack_0 <= ackL(3);
      ptr_deref_1046_load_1_ack_0 <= ackL(2);
      ptr_deref_1046_load_2_ack_0 <= ackL(1);
      ptr_deref_1046_load_3_ack_0 <= ackL(0);
      reqR(22) <= ptr_deref_553_load_3_req_1;
      reqR(21) <= ptr_deref_553_load_0_req_1;
      reqR(20) <= ptr_deref_616_load_2_req_1;
      reqR(19) <= ptr_deref_553_load_1_req_1;
      reqR(18) <= ptr_deref_616_load_3_req_1;
      reqR(17) <= ptr_deref_569_load_0_req_1;
      reqR(16) <= ptr_deref_553_load_2_req_1;
      reqR(15) <= ptr_deref_569_load_1_req_1;
      reqR(14) <= ptr_deref_569_load_2_req_1;
      reqR(13) <= ptr_deref_569_load_3_req_1;
      reqR(12) <= ptr_deref_783_load_0_req_1;
      reqR(11) <= ptr_deref_783_load_1_req_1;
      reqR(10) <= ptr_deref_616_load_1_req_1;
      reqR(9) <= ptr_deref_616_load_0_req_1;
      reqR(8) <= ptr_deref_862_load_0_req_1;
      reqR(7) <= ptr_deref_1016_load_0_req_1;
      reqR(6) <= ptr_deref_1016_load_1_req_1;
      reqR(5) <= ptr_deref_1016_load_2_req_1;
      reqR(4) <= ptr_deref_1016_load_3_req_1;
      reqR(3) <= ptr_deref_1046_load_0_req_1;
      reqR(2) <= ptr_deref_1046_load_1_req_1;
      reqR(1) <= ptr_deref_1046_load_2_req_1;
      reqR(0) <= ptr_deref_1046_load_3_req_1;
      ptr_deref_553_load_3_ack_1 <= ackR(22);
      ptr_deref_553_load_0_ack_1 <= ackR(21);
      ptr_deref_616_load_2_ack_1 <= ackR(20);
      ptr_deref_553_load_1_ack_1 <= ackR(19);
      ptr_deref_616_load_3_ack_1 <= ackR(18);
      ptr_deref_569_load_0_ack_1 <= ackR(17);
      ptr_deref_553_load_2_ack_1 <= ackR(16);
      ptr_deref_569_load_1_ack_1 <= ackR(15);
      ptr_deref_569_load_2_ack_1 <= ackR(14);
      ptr_deref_569_load_3_ack_1 <= ackR(13);
      ptr_deref_783_load_0_ack_1 <= ackR(12);
      ptr_deref_783_load_1_ack_1 <= ackR(11);
      ptr_deref_616_load_1_ack_1 <= ackR(10);
      ptr_deref_616_load_0_ack_1 <= ackR(9);
      ptr_deref_862_load_0_ack_1 <= ackR(8);
      ptr_deref_1016_load_0_ack_1 <= ackR(7);
      ptr_deref_1016_load_1_ack_1 <= ackR(6);
      ptr_deref_1016_load_2_ack_1 <= ackR(5);
      ptr_deref_1016_load_3_ack_1 <= ackR(4);
      ptr_deref_1046_load_0_ack_1 <= ackR(3);
      ptr_deref_1046_load_1_ack_1 <= ackR(2);
      ptr_deref_1046_load_2_ack_1 <= ackR(1);
      ptr_deref_1046_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_553_word_address_3 & ptr_deref_553_word_address_0 & ptr_deref_616_word_address_2 & ptr_deref_553_word_address_1 & ptr_deref_616_word_address_3 & ptr_deref_569_word_address_0 & ptr_deref_553_word_address_2 & ptr_deref_569_word_address_1 & ptr_deref_569_word_address_2 & ptr_deref_569_word_address_3 & ptr_deref_783_word_address_0 & ptr_deref_783_word_address_1 & ptr_deref_616_word_address_1 & ptr_deref_616_word_address_0 & ptr_deref_862_word_address_0 & ptr_deref_1016_word_address_0 & ptr_deref_1016_word_address_1 & ptr_deref_1016_word_address_2 & ptr_deref_1016_word_address_3 & ptr_deref_1046_word_address_0 & ptr_deref_1046_word_address_1 & ptr_deref_1046_word_address_2 & ptr_deref_1046_word_address_3;
      ptr_deref_553_data_3 <= data_out(183 downto 176);
      ptr_deref_553_data_0 <= data_out(175 downto 168);
      ptr_deref_616_data_2 <= data_out(167 downto 160);
      ptr_deref_553_data_1 <= data_out(159 downto 152);
      ptr_deref_616_data_3 <= data_out(151 downto 144);
      ptr_deref_569_data_0 <= data_out(143 downto 136);
      ptr_deref_553_data_2 <= data_out(135 downto 128);
      ptr_deref_569_data_1 <= data_out(127 downto 120);
      ptr_deref_569_data_2 <= data_out(119 downto 112);
      ptr_deref_569_data_3 <= data_out(111 downto 104);
      ptr_deref_783_data_0 <= data_out(103 downto 96);
      ptr_deref_783_data_1 <= data_out(95 downto 88);
      ptr_deref_616_data_1 <= data_out(87 downto 80);
      ptr_deref_616_data_0 <= data_out(79 downto 72);
      ptr_deref_862_data_0 <= data_out(71 downto 64);
      ptr_deref_1016_data_0 <= data_out(63 downto 56);
      ptr_deref_1016_data_1 <= data_out(55 downto 48);
      ptr_deref_1016_data_2 <= data_out(47 downto 40);
      ptr_deref_1016_data_3 <= data_out(39 downto 32);
      ptr_deref_1046_data_0 <= data_out(31 downto 24);
      ptr_deref_1046_data_1 <= data_out(23 downto 16);
      ptr_deref_1046_data_2 <= data_out(15 downto 8);
      ptr_deref_1046_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 23,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 23,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_939_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_939_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_939_word_address_0) &  " data ptr_deref_939_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_939_data_0) severity note; --
        end if;
        if ptr_deref_939_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_939_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_939_word_address_3) &  " data ptr_deref_939_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_939_data_3) severity note; --
        end if;
        if ptr_deref_939_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_939_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_939_word_address_1) &  " data ptr_deref_939_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_939_data_1) severity note; --
        end if;
        if ptr_deref_939_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_939_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_939_word_address_2) &  " data ptr_deref_939_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_939_data_2) severity note; --
        end if;
        if ptr_deref_960_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_960_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_960_word_address_0) &  " data ptr_deref_960_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_960_data_0) severity note; --
        end if;
        if ptr_deref_960_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_960_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_960_word_address_1) &  " data ptr_deref_960_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_960_data_1) severity note; --
        end if;
        if ptr_deref_960_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_960_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_960_word_address_2) &  " data ptr_deref_960_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_960_data_2) severity note; --
        end if;
        if ptr_deref_960_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_960_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_960_word_address_3) &  " data ptr_deref_960_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_960_data_3) severity note; --
        end if;
        if ptr_deref_1002_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1002_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1002_word_address_0) &  " data ptr_deref_1002_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1002_data_0) severity note; --
        end if;
        if ptr_deref_1002_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1002_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1002_word_address_1) &  " data ptr_deref_1002_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1002_data_1) severity note; --
        end if;
        if ptr_deref_1002_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1002_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1002_word_address_2) &  " data ptr_deref_1002_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1002_data_2) severity note; --
        end if;
        if ptr_deref_1002_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1002_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1002_word_address_3) &  " data ptr_deref_1002_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1002_data_3) severity note; --
        end if;
        if ptr_deref_1030_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1030_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1030_word_address_0) &  " data ptr_deref_1030_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1030_data_0) severity note; --
        end if;
        if ptr_deref_1030_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1030_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1030_word_address_1) &  " data ptr_deref_1030_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1030_data_1) severity note; --
        end if;
        if ptr_deref_1030_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1030_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1030_word_address_2) &  " data ptr_deref_1030_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1030_data_2) severity note; --
        end if;
        if ptr_deref_1030_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1030_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1030_word_address_3) &  " data ptr_deref_1030_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1030_data_3) severity note; --
        end if;
        if ptr_deref_1060_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1060_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1060_word_address_0) &  " data ptr_deref_1060_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1060_data_0) severity note; --
        end if;
        if ptr_deref_1060_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1060_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1060_word_address_1) &  " data ptr_deref_1060_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1060_data_1) severity note; --
        end if;
        if ptr_deref_1060_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1060_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1060_word_address_2) &  " data ptr_deref_1060_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1060_data_2) severity note; --
        end if;
        if ptr_deref_1060_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1060_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1060_word_address_3) &  " data ptr_deref_1060_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1060_data_3) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_939_store_0 ptr_deref_939_store_3 ptr_deref_939_store_1 ptr_deref_939_store_2 ptr_deref_960_store_0 ptr_deref_960_store_1 ptr_deref_960_store_2 ptr_deref_960_store_3 ptr_deref_1002_store_0 ptr_deref_1002_store_1 ptr_deref_1002_store_2 ptr_deref_1002_store_3 ptr_deref_1030_store_0 ptr_deref_1030_store_1 ptr_deref_1030_store_2 ptr_deref_1030_store_3 ptr_deref_1060_store_0 ptr_deref_1060_store_1 ptr_deref_1060_store_2 ptr_deref_1060_store_3 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(319 downto 0);
      signal data_in: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 19 downto 0);
      -- 
    begin -- 
      reqL(19) <= ptr_deref_939_store_0_req_0;
      reqL(18) <= ptr_deref_939_store_3_req_0;
      reqL(17) <= ptr_deref_939_store_1_req_0;
      reqL(16) <= ptr_deref_939_store_2_req_0;
      reqL(15) <= ptr_deref_960_store_0_req_0;
      reqL(14) <= ptr_deref_960_store_1_req_0;
      reqL(13) <= ptr_deref_960_store_2_req_0;
      reqL(12) <= ptr_deref_960_store_3_req_0;
      reqL(11) <= ptr_deref_1002_store_0_req_0;
      reqL(10) <= ptr_deref_1002_store_1_req_0;
      reqL(9) <= ptr_deref_1002_store_2_req_0;
      reqL(8) <= ptr_deref_1002_store_3_req_0;
      reqL(7) <= ptr_deref_1030_store_0_req_0;
      reqL(6) <= ptr_deref_1030_store_1_req_0;
      reqL(5) <= ptr_deref_1030_store_2_req_0;
      reqL(4) <= ptr_deref_1030_store_3_req_0;
      reqL(3) <= ptr_deref_1060_store_0_req_0;
      reqL(2) <= ptr_deref_1060_store_1_req_0;
      reqL(1) <= ptr_deref_1060_store_2_req_0;
      reqL(0) <= ptr_deref_1060_store_3_req_0;
      ptr_deref_939_store_0_ack_0 <= ackL(19);
      ptr_deref_939_store_3_ack_0 <= ackL(18);
      ptr_deref_939_store_1_ack_0 <= ackL(17);
      ptr_deref_939_store_2_ack_0 <= ackL(16);
      ptr_deref_960_store_0_ack_0 <= ackL(15);
      ptr_deref_960_store_1_ack_0 <= ackL(14);
      ptr_deref_960_store_2_ack_0 <= ackL(13);
      ptr_deref_960_store_3_ack_0 <= ackL(12);
      ptr_deref_1002_store_0_ack_0 <= ackL(11);
      ptr_deref_1002_store_1_ack_0 <= ackL(10);
      ptr_deref_1002_store_2_ack_0 <= ackL(9);
      ptr_deref_1002_store_3_ack_0 <= ackL(8);
      ptr_deref_1030_store_0_ack_0 <= ackL(7);
      ptr_deref_1030_store_1_ack_0 <= ackL(6);
      ptr_deref_1030_store_2_ack_0 <= ackL(5);
      ptr_deref_1030_store_3_ack_0 <= ackL(4);
      ptr_deref_1060_store_0_ack_0 <= ackL(3);
      ptr_deref_1060_store_1_ack_0 <= ackL(2);
      ptr_deref_1060_store_2_ack_0 <= ackL(1);
      ptr_deref_1060_store_3_ack_0 <= ackL(0);
      reqR(19) <= ptr_deref_939_store_0_req_1;
      reqR(18) <= ptr_deref_939_store_3_req_1;
      reqR(17) <= ptr_deref_939_store_1_req_1;
      reqR(16) <= ptr_deref_939_store_2_req_1;
      reqR(15) <= ptr_deref_960_store_0_req_1;
      reqR(14) <= ptr_deref_960_store_1_req_1;
      reqR(13) <= ptr_deref_960_store_2_req_1;
      reqR(12) <= ptr_deref_960_store_3_req_1;
      reqR(11) <= ptr_deref_1002_store_0_req_1;
      reqR(10) <= ptr_deref_1002_store_1_req_1;
      reqR(9) <= ptr_deref_1002_store_2_req_1;
      reqR(8) <= ptr_deref_1002_store_3_req_1;
      reqR(7) <= ptr_deref_1030_store_0_req_1;
      reqR(6) <= ptr_deref_1030_store_1_req_1;
      reqR(5) <= ptr_deref_1030_store_2_req_1;
      reqR(4) <= ptr_deref_1030_store_3_req_1;
      reqR(3) <= ptr_deref_1060_store_0_req_1;
      reqR(2) <= ptr_deref_1060_store_1_req_1;
      reqR(1) <= ptr_deref_1060_store_2_req_1;
      reqR(0) <= ptr_deref_1060_store_3_req_1;
      ptr_deref_939_store_0_ack_1 <= ackR(19);
      ptr_deref_939_store_3_ack_1 <= ackR(18);
      ptr_deref_939_store_1_ack_1 <= ackR(17);
      ptr_deref_939_store_2_ack_1 <= ackR(16);
      ptr_deref_960_store_0_ack_1 <= ackR(15);
      ptr_deref_960_store_1_ack_1 <= ackR(14);
      ptr_deref_960_store_2_ack_1 <= ackR(13);
      ptr_deref_960_store_3_ack_1 <= ackR(12);
      ptr_deref_1002_store_0_ack_1 <= ackR(11);
      ptr_deref_1002_store_1_ack_1 <= ackR(10);
      ptr_deref_1002_store_2_ack_1 <= ackR(9);
      ptr_deref_1002_store_3_ack_1 <= ackR(8);
      ptr_deref_1030_store_0_ack_1 <= ackR(7);
      ptr_deref_1030_store_1_ack_1 <= ackR(6);
      ptr_deref_1030_store_2_ack_1 <= ackR(5);
      ptr_deref_1030_store_3_ack_1 <= ackR(4);
      ptr_deref_1060_store_0_ack_1 <= ackR(3);
      ptr_deref_1060_store_1_ack_1 <= ackR(2);
      ptr_deref_1060_store_2_ack_1 <= ackR(1);
      ptr_deref_1060_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_939_word_address_0 & ptr_deref_939_word_address_3 & ptr_deref_939_word_address_1 & ptr_deref_939_word_address_2 & ptr_deref_960_word_address_0 & ptr_deref_960_word_address_1 & ptr_deref_960_word_address_2 & ptr_deref_960_word_address_3 & ptr_deref_1002_word_address_0 & ptr_deref_1002_word_address_1 & ptr_deref_1002_word_address_2 & ptr_deref_1002_word_address_3 & ptr_deref_1030_word_address_0 & ptr_deref_1030_word_address_1 & ptr_deref_1030_word_address_2 & ptr_deref_1030_word_address_3 & ptr_deref_1060_word_address_0 & ptr_deref_1060_word_address_1 & ptr_deref_1060_word_address_2 & ptr_deref_1060_word_address_3;
      data_in <= ptr_deref_939_data_0 & ptr_deref_939_data_3 & ptr_deref_939_data_1 & ptr_deref_939_data_2 & ptr_deref_960_data_0 & ptr_deref_960_data_1 & ptr_deref_960_data_2 & ptr_deref_960_data_3 & ptr_deref_1002_data_0 & ptr_deref_1002_data_1 & ptr_deref_1002_data_2 & ptr_deref_1002_data_3 & ptr_deref_1030_data_0 & ptr_deref_1030_data_1 & ptr_deref_1030_data_2 & ptr_deref_1030_data_3 & ptr_deref_1060_data_0 & ptr_deref_1060_data_1 & ptr_deref_1060_data_2 & ptr_deref_1060_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 20,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 20,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_537_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_537_inst_ack_0 then -- 
            assert false report " ReadPipe chk_in0 to wire simple_obj_ref_537_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_537_inst_req_0;
      simple_obj_ref_537_inst_ack_0 <= ack(0);
      simple_obj_ref_537_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => chk_in0_pipe_read_req(0),
          oack => chk_in0_pipe_read_ack(0),
          odata => chk_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1080_inst_ack_0 then -- 
          assert false report " WritePipe rtt_in0 from wire type_cast_1082_wire value="  &  convert_slv_to_hex_string(type_cast_1082_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_1080_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1080_inst_req_0;
      simple_obj_ref_1080_inst_ack_0 <= ack(0);
      data_in <= type_cast_1082_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => rtt_in0_pipe_write_req(0),
          oack => rtt_in0_pipe_write_ack(0),
          odata => rtt_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_710_call call_stmt_677_call call_stmt_648_call call_stmt_928_call call_stmt_607_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      reqL(4) <= call_stmt_710_call_req_0;
      reqL(3) <= call_stmt_677_call_req_0;
      reqL(2) <= call_stmt_648_call_req_0;
      reqL(1) <= call_stmt_928_call_req_0;
      reqL(0) <= call_stmt_607_call_req_0;
      call_stmt_710_call_ack_0 <= ackL(4);
      call_stmt_677_call_ack_0 <= ackL(3);
      call_stmt_648_call_ack_0 <= ackL(2);
      call_stmt_928_call_ack_0 <= ackL(1);
      call_stmt_607_call_ack_0 <= ackL(0);
      reqR(4) <= call_stmt_710_call_req_1;
      reqR(3) <= call_stmt_677_call_req_1;
      reqR(2) <= call_stmt_648_call_req_1;
      reqR(1) <= call_stmt_928_call_req_1;
      reqR(0) <= call_stmt_607_call_req_1;
      call_stmt_710_call_ack_1 <= ackR(4);
      call_stmt_677_call_ack_1 <= ackR(3);
      call_stmt_648_call_ack_1 <= ackR(2);
      call_stmt_928_call_ack_1 <= ackR(1);
      call_stmt_607_call_ack_1 <= ackR(0);
      data_in <= tmp13_539 & tmp13_539 & tmp13_539 & tmp13_539 & tmp13_539;
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 160,
        owidth => 32,
        twidth => 3,
        nreqs => 5,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_packet_free_call_reqs(0),
          ackR => ahir_packet_free_call_acks(0),
          dataR => ahir_packet_free_call_data(31 downto 0),
          tagR => ahir_packet_free_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 3, nreqs => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => ahir_packet_free_return_acks(0), -- cross-over
          ackL => ahir_packet_free_return_reqs(0), -- cross-over
          tagL => ahir_packet_free_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_682_call 
    CallGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_682_call_req_0;
      call_stmt_682_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_682_call_req_1;
      call_stmt_682_call_ack_1 <= ackR(0);
      data_in <= tmp35x_xi_639;
      tmp32_682 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 16,
        owidth => 16,
        twidth => 2,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 16, twidth => 2, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_rtt is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(4 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    rtt_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    rtt_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    rtt_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    to0_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to0_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to0_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    to1_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to1_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to1_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    to2_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to2_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to2_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    to3_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to3_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to3_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_packet_free_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_free_call_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_free_call_data : out  std_logic_vector(31 downto 0);
    ahir_packet_free_call_tag  :  out  std_logic_vector(2 downto 0);
    ahir_packet_free_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_free_return_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_free_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_rtt;
architecture Default of ahir_glue_rtt is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_rtt_CP_4152_start: Boolean;
  -- links between control-path and data-path
  signal binary_1157_inst_req_0 : boolean;
  signal binary_1203_inst_req_0 : boolean;
  signal if_stmt_1159_branch_ack_0 : boolean;
  signal binary_1203_inst_ack_1 : boolean;
  signal ptr_deref_1137_addr_0_req_0 : boolean;
  signal ptr_deref_1137_load_0_req_0 : boolean;
  signal binary_1157_inst_ack_0 : boolean;
  signal type_cast_1199_inst_ack_0 : boolean;
  signal ptr_deref_1141_gather_scatter_ack_0 : boolean;
  signal binary_1271_inst_req_0 : boolean;
  signal ptr_deref_1137_load_0_req_1 : boolean;
  signal if_stmt_1190_branch_ack_1 : boolean;
  signal ptr_deref_1137_load_0_ack_0 : boolean;
  signal addr_of_1261_final_reg_ack_0 : boolean;
  signal ptr_deref_1137_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1265_base_resize_ack_0 : boolean;
  signal binary_1151_inst_req_1 : boolean;
  signal binary_1203_inst_req_1 : boolean;
  signal if_stmt_1190_branch_ack_0 : boolean;
  signal binary_1203_inst_ack_0 : boolean;
  signal if_stmt_1190_branch_req_0 : boolean;
  signal binary_1151_inst_ack_0 : boolean;
  signal if_stmt_1205_branch_req_0 : boolean;
  signal ptr_deref_1265_root_address_inst_ack_0 : boolean;
  signal binary_1151_inst_req_0 : boolean;
  signal ptr_deref_1137_root_address_inst_req_0 : boolean;
  signal binary_1219_inst_req_1 : boolean;
  signal type_cast_1199_inst_req_0 : boolean;
  signal ptr_deref_1265_base_resize_req_0 : boolean;
  signal simple_obj_ref_1213_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1265_load_0_req_0 : boolean;
  signal addr_of_1261_final_reg_req_0 : boolean;
  signal ptr_deref_1265_load_0_ack_0 : boolean;
  signal array_obj_ref_1260_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1260_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_1213_gather_scatter_req_0 : boolean;
  signal ptr_deref_1265_root_address_inst_req_0 : boolean;
  signal binary_1188_inst_req_1 : boolean;
  signal ptr_deref_1141_load_0_ack_1 : boolean;
  signal addr_of_1285_final_reg_req_0 : boolean;
  signal ptr_deref_1265_gather_scatter_req_0 : boolean;
  signal type_cast_1184_inst_req_0 : boolean;
  signal ptr_deref_1141_gather_scatter_req_0 : boolean;
  signal binary_1271_inst_ack_0 : boolean;
  signal binary_1219_inst_ack_1 : boolean;
  signal ptr_deref_1265_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1213_load_0_ack_1 : boolean;
  signal addr_of_1285_final_reg_ack_0 : boolean;
  signal ptr_deref_1137_base_resize_ack_0 : boolean;
  signal array_obj_ref_1284_offset_inst_req_0 : boolean;
  signal ptr_deref_1141_load_0_req_1 : boolean;
  signal array_obj_ref_1260_offset_inst_ack_0 : boolean;
  signal simple_obj_ref_1213_load_0_req_1 : boolean;
  signal array_obj_ref_1284_offset_inst_ack_0 : boolean;
  signal binary_1151_inst_ack_1 : boolean;
  signal binary_1157_inst_req_1 : boolean;
  signal binary_1188_inst_ack_1 : boolean;
  signal array_obj_ref_1284_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1284_index_sum_1_ack_1 : boolean;
  signal binary_1146_inst_req_0 : boolean;
  signal binary_1146_inst_ack_0 : boolean;
  signal ptr_deref_1137_addr_0_ack_0 : boolean;
  signal ptr_deref_1137_base_resize_req_0 : boolean;
  signal addr_of_1133_final_reg_ack_0 : boolean;
  signal binary_1188_inst_ack_0 : boolean;
  signal ptr_deref_1137_load_0_ack_1 : boolean;
  signal binary_1146_inst_req_1 : boolean;
  signal array_obj_ref_1284_index_sum_1_req_0 : boolean;
  signal ptr_deref_1141_load_0_ack_0 : boolean;
  signal binary_1157_inst_ack_1 : boolean;
  signal array_obj_ref_1260_index_sum_1_req_0 : boolean;
  signal binary_1146_inst_ack_1 : boolean;
  signal array_obj_ref_1260_index_sum_1_ack_0 : boolean;
  signal binary_1271_inst_ack_1 : boolean;
  signal binary_1219_inst_ack_0 : boolean;
  signal array_obj_ref_1260_offset_inst_req_0 : boolean;
  signal ptr_deref_1141_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1260_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1260_index_sum_1_ack_1 : boolean;
  signal ptr_deref_1265_addr_0_req_0 : boolean;
  signal if_stmt_1159_branch_ack_1 : boolean;
  signal if_stmt_1273_branch_req_0 : boolean;
  signal ptr_deref_1137_gather_scatter_req_0 : boolean;
  signal binary_1219_inst_req_0 : boolean;
  signal binary_1300_inst_req_0 : boolean;
  signal array_obj_ref_1260_index_0_scale_ack_1 : boolean;
  signal binary_1300_inst_req_1 : boolean;
  signal binary_1188_inst_req_0 : boolean;
  signal ptr_deref_1141_load_0_req_0 : boolean;
  signal array_obj_ref_1260_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1260_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1260_index_0_scale_req_0 : boolean;
  signal ptr_deref_1137_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1213_load_0_ack_0 : boolean;
  signal type_cast_1184_inst_ack_0 : boolean;
  signal array_obj_ref_1260_index_0_resize_ack_0 : boolean;
  signal type_cast_1094_inst_ack_0 : boolean;
  signal array_obj_ref_1260_index_0_resize_req_0 : boolean;
  signal simple_obj_ref_1093_inst_req_0 : boolean;
  signal if_stmt_1273_branch_ack_1 : boolean;
  signal simple_obj_ref_1093_inst_ack_0 : boolean;
  signal array_obj_ref_1284_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1105_base_resize_req_0 : boolean;
  signal binary_1300_inst_ack_0 : boolean;
  signal if_stmt_1159_branch_req_0 : boolean;
  signal type_cast_1098_inst_ack_0 : boolean;
  signal addr_of_1133_final_reg_req_0 : boolean;
  signal array_obj_ref_1105_base_resize_ack_0 : boolean;
  signal array_obj_ref_1284_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1105_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1284_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1132_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_1213_load_0_req_0 : boolean;
  signal array_obj_ref_1105_final_reg_req_0 : boolean;
  signal array_obj_ref_1105_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1284_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1105_final_reg_ack_0 : boolean;
  signal ptr_deref_1265_load_0_ack_1 : boolean;
  signal type_cast_1094_inst_req_0 : boolean;
  signal array_obj_ref_1105_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1105_root_address_inst_ack_0 : boolean;
  signal type_cast_1098_inst_req_0 : boolean;
  signal ptr_deref_1458_root_address_inst_req_0 : boolean;
  signal ptr_deref_1458_root_address_inst_ack_0 : boolean;
  signal type_cast_1109_inst_req_0 : boolean;
  signal if_stmt_1232_branch_ack_0 : boolean;
  signal type_cast_1109_inst_ack_0 : boolean;
  signal ptr_deref_1265_load_0_req_1 : boolean;
  signal if_stmt_1321_branch_ack_0 : boolean;
  signal binary_1319_inst_req_0 : boolean;
  signal binary_1300_inst_ack_1 : boolean;
  signal if_stmt_1308_branch_req_0 : boolean;
  signal if_stmt_1205_branch_ack_0 : boolean;
  signal if_stmt_1308_branch_ack_1 : boolean;
  signal binary_1306_inst_req_0 : boolean;
  signal binary_1319_inst_ack_0 : boolean;
  signal binary_1319_inst_req_1 : boolean;
  signal binary_1319_inst_ack_1 : boolean;
  signal ptr_deref_1141_base_resize_req_0 : boolean;
  signal if_stmt_1205_branch_ack_1 : boolean;
  signal if_stmt_1308_branch_ack_0 : boolean;
  signal binary_1271_inst_req_1 : boolean;
  signal binary_1306_inst_req_1 : boolean;
  signal binary_1306_inst_ack_1 : boolean;
  signal if_stmt_1321_branch_ack_1 : boolean;
  signal ptr_deref_1141_base_resize_ack_0 : boolean;
  signal if_stmt_1321_branch_req_0 : boolean;
  signal ptr_deref_1141_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_1221_gather_scatter_req_0 : boolean;
  signal binary_1306_inst_ack_0 : boolean;
  signal simple_obj_ref_1221_gather_scatter_ack_0 : boolean;
  signal binary_1170_inst_ack_1 : boolean;
  signal binary_1170_inst_req_1 : boolean;
  signal if_stmt_1232_branch_ack_1 : boolean;
  signal binary_1170_inst_ack_0 : boolean;
  signal binary_1170_inst_req_0 : boolean;
  signal ptr_deref_1141_addr_0_ack_0 : boolean;
  signal if_stmt_1232_branch_req_0 : boolean;
  signal ptr_deref_1113_base_resize_req_0 : boolean;
  signal ptr_deref_1113_base_resize_ack_0 : boolean;
  signal ptr_deref_1141_addr_0_req_0 : boolean;
  signal ptr_deref_1113_root_address_inst_req_0 : boolean;
  signal ptr_deref_1113_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1284_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1284_index_0_scale_req_1 : boolean;
  signal ptr_deref_1113_addr_0_req_0 : boolean;
  signal ptr_deref_1113_addr_0_ack_0 : boolean;
  signal binary_1230_inst_ack_1 : boolean;
  signal ptr_deref_1113_addr_0_req_1 : boolean;
  signal array_obj_ref_1132_root_address_inst_req_0 : boolean;
  signal binary_1230_inst_req_1 : boolean;
  signal ptr_deref_1113_addr_0_ack_1 : boolean;
  signal binary_1230_inst_ack_0 : boolean;
  signal ptr_deref_1113_addr_1_req_0 : boolean;
  signal binary_1230_inst_req_0 : boolean;
  signal ptr_deref_1113_addr_1_ack_0 : boolean;
  signal ptr_deref_1113_addr_1_req_1 : boolean;
  signal ptr_deref_1113_addr_1_ack_1 : boolean;
  signal array_obj_ref_1284_index_0_scale_ack_0 : boolean;
  signal ptr_deref_1113_addr_2_req_0 : boolean;
  signal type_cast_1226_inst_ack_0 : boolean;
  signal ptr_deref_1113_addr_2_ack_0 : boolean;
  signal type_cast_1226_inst_req_0 : boolean;
  signal ptr_deref_1113_addr_2_req_1 : boolean;
  signal ptr_deref_1113_addr_2_ack_1 : boolean;
  signal ptr_deref_1113_addr_3_req_0 : boolean;
  signal ptr_deref_1113_addr_3_ack_0 : boolean;
  signal ptr_deref_1113_addr_3_req_1 : boolean;
  signal array_obj_ref_1132_offset_inst_ack_0 : boolean;
  signal ptr_deref_1113_addr_3_ack_1 : boolean;
  signal array_obj_ref_1284_index_0_scale_req_0 : boolean;
  signal ptr_deref_1113_load_0_req_0 : boolean;
  signal ptr_deref_1113_load_0_ack_0 : boolean;
  signal ptr_deref_1113_load_1_req_0 : boolean;
  signal ptr_deref_1113_load_1_ack_0 : boolean;
  signal ptr_deref_1113_load_2_req_0 : boolean;
  signal simple_obj_ref_1221_store_0_ack_1 : boolean;
  signal ptr_deref_1113_load_2_ack_0 : boolean;
  signal simple_obj_ref_1221_store_0_req_1 : boolean;
  signal ptr_deref_1113_load_3_req_0 : boolean;
  signal ptr_deref_1113_load_3_ack_0 : boolean;
  signal ptr_deref_1113_load_0_req_1 : boolean;
  signal ptr_deref_1113_load_0_ack_1 : boolean;
  signal array_obj_ref_1284_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1113_load_1_req_1 : boolean;
  signal ptr_deref_1113_load_1_ack_1 : boolean;
  signal ptr_deref_1113_load_2_req_1 : boolean;
  signal ptr_deref_1113_load_2_ack_1 : boolean;
  signal ptr_deref_1113_load_3_req_1 : boolean;
  signal ptr_deref_1113_load_3_ack_1 : boolean;
  signal if_stmt_1273_branch_ack_0 : boolean;
  signal simple_obj_ref_1221_store_0_ack_0 : boolean;
  signal ptr_deref_1113_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1221_store_0_req_0 : boolean;
  signal ptr_deref_1113_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1265_addr_0_ack_0 : boolean;
  signal ptr_deref_1442_load_3_req_1 : boolean;
  signal if_stmt_1449_branch_ack_1 : boolean;
  signal ptr_deref_1442_load_2_ack_1 : boolean;
  signal array_obj_ref_1123_index_0_resize_req_0 : boolean;
  signal ptr_deref_1442_load_3_ack_1 : boolean;
  signal array_obj_ref_1123_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1123_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1123_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1123_index_0_scale_req_1 : boolean;
  signal ptr_deref_1442_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1123_index_0_scale_ack_1 : boolean;
  signal binary_1447_inst_req_0 : boolean;
  signal ptr_deref_1442_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1123_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1123_index_sum_1_ack_0 : boolean;
  signal binary_1447_inst_ack_0 : boolean;
  signal if_stmt_1449_branch_ack_0 : boolean;
  signal array_obj_ref_1123_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1123_index_sum_1_ack_1 : boolean;
  signal binary_1447_inst_req_1 : boolean;
  signal array_obj_ref_1123_offset_inst_req_0 : boolean;
  signal array_obj_ref_1123_offset_inst_ack_0 : boolean;
  signal ptr_deref_1458_base_resize_req_0 : boolean;
  signal ptr_deref_1458_base_resize_ack_0 : boolean;
  signal array_obj_ref_1123_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1123_root_address_inst_ack_0 : boolean;
  signal binary_1447_inst_ack_1 : boolean;
  signal addr_of_1124_final_reg_req_0 : boolean;
  signal addr_of_1124_final_reg_ack_0 : boolean;
  signal array_obj_ref_1132_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1132_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1132_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1132_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1132_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1132_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1132_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1132_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1132_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1132_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1132_offset_inst_req_0 : boolean;
  signal array_obj_ref_1333_offset_inst_req_0 : boolean;
  signal array_obj_ref_1333_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1333_base_resize_req_0 : boolean;
  signal array_obj_ref_1333_base_resize_ack_0 : boolean;
  signal array_obj_ref_1333_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1333_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1333_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1333_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1333_final_reg_req_0 : boolean;
  signal array_obj_ref_1333_final_reg_ack_0 : boolean;
  signal ptr_deref_1336_base_resize_req_0 : boolean;
  signal ptr_deref_1336_base_resize_ack_0 : boolean;
  signal ptr_deref_1336_root_address_inst_req_0 : boolean;
  signal phi_stmt_1289_ack_0 : boolean;
  signal ptr_deref_1336_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1336_addr_0_req_0 : boolean;
  signal ptr_deref_1336_addr_0_ack_0 : boolean;
  signal ptr_deref_1336_gather_scatter_req_0 : boolean;
  signal ptr_deref_1336_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1336_store_0_req_0 : boolean;
  signal ptr_deref_1336_store_0_ack_0 : boolean;
  signal ptr_deref_1336_store_0_req_1 : boolean;
  signal phi_stmt_1248_req_1 : boolean;
  signal ptr_deref_1336_store_0_ack_1 : boolean;
  signal array_obj_ref_1343_base_resize_req_0 : boolean;
  signal array_obj_ref_1343_base_resize_ack_0 : boolean;
  signal array_obj_ref_1343_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1343_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1343_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1343_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1343_final_reg_req_0 : boolean;
  signal array_obj_ref_1343_final_reg_ack_0 : boolean;
  signal type_cast_1347_inst_req_0 : boolean;
  signal type_cast_1347_inst_ack_0 : boolean;
  signal ptr_deref_1350_base_resize_req_0 : boolean;
  signal ptr_deref_1350_base_resize_ack_0 : boolean;
  signal ptr_deref_1350_root_address_inst_req_0 : boolean;
  signal ptr_deref_1350_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1350_addr_0_req_0 : boolean;
  signal ptr_deref_1350_addr_0_ack_0 : boolean;
  signal ptr_deref_1350_addr_0_req_1 : boolean;
  signal phi_stmt_1241_req_1 : boolean;
  signal ptr_deref_1350_addr_0_ack_1 : boolean;
  signal ptr_deref_1350_addr_1_req_0 : boolean;
  signal ptr_deref_1350_addr_1_ack_0 : boolean;
  signal ptr_deref_1350_addr_1_req_1 : boolean;
  signal ptr_deref_1350_addr_1_ack_1 : boolean;
  signal ptr_deref_1350_addr_2_req_0 : boolean;
  signal ptr_deref_1350_addr_2_ack_0 : boolean;
  signal ptr_deref_1350_addr_2_req_1 : boolean;
  signal ptr_deref_1350_addr_2_ack_1 : boolean;
  signal ptr_deref_1350_addr_3_req_0 : boolean;
  signal ptr_deref_1350_addr_3_ack_0 : boolean;
  signal ptr_deref_1350_addr_3_req_1 : boolean;
  signal ptr_deref_1350_addr_3_ack_1 : boolean;
  signal ptr_deref_1350_gather_scatter_req_0 : boolean;
  signal ptr_deref_1350_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1350_store_0_req_0 : boolean;
  signal ptr_deref_1350_store_0_ack_0 : boolean;
  signal ptr_deref_1350_store_1_req_0 : boolean;
  signal ptr_deref_1350_store_1_ack_0 : boolean;
  signal ptr_deref_1350_store_2_req_0 : boolean;
  signal ptr_deref_1350_store_2_ack_0 : boolean;
  signal type_cast_1294_inst_req_0 : boolean;
  signal ptr_deref_1350_store_3_req_0 : boolean;
  signal ptr_deref_1350_store_3_ack_0 : boolean;
  signal ptr_deref_1350_store_0_req_1 : boolean;
  signal ptr_deref_1350_store_0_ack_1 : boolean;
  signal ptr_deref_1350_store_1_req_1 : boolean;
  signal ptr_deref_1350_store_1_ack_1 : boolean;
  signal ptr_deref_1350_store_2_req_1 : boolean;
  signal ptr_deref_1350_store_2_ack_1 : boolean;
  signal type_cast_1294_inst_ack_0 : boolean;
  signal ptr_deref_1350_store_3_req_1 : boolean;
  signal ptr_deref_1350_store_3_ack_1 : boolean;
  signal phi_stmt_1289_req_1 : boolean;
  signal array_obj_ref_1357_base_resize_req_0 : boolean;
  signal array_obj_ref_1357_base_resize_ack_0 : boolean;
  signal array_obj_ref_1357_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1357_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1357_root_address_inst_req_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal array_obj_ref_1357_root_address_inst_ack_1 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal array_obj_ref_1357_final_reg_req_0 : boolean;
  signal array_obj_ref_1357_final_reg_ack_0 : boolean;
  signal phi_stmt_1248_req_0 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_1292_inst_req_0 : boolean;
  signal type_cast_1365_inst_req_0 : boolean;
  signal type_cast_1365_inst_ack_0 : boolean;
  signal ptr_deref_1368_base_resize_req_0 : boolean;
  signal ptr_deref_1368_base_resize_ack_0 : boolean;
  signal ptr_deref_1368_root_address_inst_req_0 : boolean;
  signal ptr_deref_1368_root_address_inst_ack_0 : boolean;
  signal type_cast_1244_inst_req_0 : boolean;
  signal type_cast_1292_inst_ack_0 : boolean;
  signal ptr_deref_1368_addr_0_req_0 : boolean;
  signal ptr_deref_1368_addr_0_ack_0 : boolean;
  signal ptr_deref_1368_addr_0_req_1 : boolean;
  signal ptr_deref_1368_addr_0_ack_1 : boolean;
  signal ptr_deref_1368_addr_1_req_0 : boolean;
  signal ptr_deref_1368_addr_1_ack_0 : boolean;
  signal ptr_deref_1368_addr_1_req_1 : boolean;
  signal type_cast_1244_inst_ack_0 : boolean;
  signal ptr_deref_1368_addr_1_ack_1 : boolean;
  signal ptr_deref_1368_addr_2_req_0 : boolean;
  signal phi_stmt_1241_req_0 : boolean;
  signal ptr_deref_1368_addr_2_ack_0 : boolean;
  signal ptr_deref_1368_addr_2_req_1 : boolean;
  signal ptr_deref_1368_addr_2_ack_1 : boolean;
  signal ptr_deref_1368_addr_3_req_0 : boolean;
  signal ptr_deref_1368_addr_3_ack_0 : boolean;
  signal ptr_deref_1368_addr_3_req_1 : boolean;
  signal ptr_deref_1368_addr_3_ack_1 : boolean;
  signal ptr_deref_1368_gather_scatter_req_0 : boolean;
  signal ptr_deref_1368_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1368_store_0_req_0 : boolean;
  signal ptr_deref_1368_store_0_ack_0 : boolean;
  signal ptr_deref_1368_store_1_req_0 : boolean;
  signal ptr_deref_1368_store_1_ack_0 : boolean;
  signal ptr_deref_1368_store_2_req_0 : boolean;
  signal ptr_deref_1368_store_2_ack_0 : boolean;
  signal phi_stmt_1241_ack_0 : boolean;
  signal ptr_deref_1368_store_3_req_0 : boolean;
  signal ptr_deref_1368_store_3_ack_0 : boolean;
  signal phi_stmt_1248_ack_0 : boolean;
  signal ptr_deref_1368_store_0_req_1 : boolean;
  signal ptr_deref_1368_store_0_ack_1 : boolean;
  signal ptr_deref_1368_store_1_req_1 : boolean;
  signal ptr_deref_1368_store_1_ack_1 : boolean;
  signal ptr_deref_1368_store_2_req_1 : boolean;
  signal ptr_deref_1368_store_2_ack_1 : boolean;
  signal ptr_deref_1368_store_3_req_1 : boolean;
  signal ptr_deref_1368_store_3_ack_1 : boolean;
  signal type_cast_1374_inst_req_0 : boolean;
  signal type_cast_1374_inst_ack_0 : boolean;
  signal array_obj_ref_1383_base_resize_req_0 : boolean;
  signal phi_stmt_1289_req_0 : boolean;
  signal array_obj_ref_1383_base_resize_ack_0 : boolean;
  signal array_obj_ref_1383_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1383_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1383_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1383_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1383_final_reg_req_0 : boolean;
  signal array_obj_ref_1383_final_reg_ack_0 : boolean;
  signal binary_1389_inst_req_0 : boolean;
  signal binary_1389_inst_ack_0 : boolean;
  signal binary_1389_inst_req_1 : boolean;
  signal binary_1389_inst_ack_1 : boolean;
  signal if_stmt_1391_branch_req_0 : boolean;
  signal if_stmt_1391_branch_ack_1 : boolean;
  signal if_stmt_1391_branch_ack_0 : boolean;
  signal ptr_deref_1399_base_resize_req_0 : boolean;
  signal ptr_deref_1399_base_resize_ack_0 : boolean;
  signal ptr_deref_1399_root_address_inst_req_0 : boolean;
  signal ptr_deref_1399_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1399_addr_0_req_0 : boolean;
  signal ptr_deref_1399_addr_0_ack_0 : boolean;
  signal ptr_deref_1399_gather_scatter_req_0 : boolean;
  signal ptr_deref_1399_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1399_store_0_req_0 : boolean;
  signal ptr_deref_1399_store_0_ack_0 : boolean;
  signal ptr_deref_1399_store_0_req_1 : boolean;
  signal ptr_deref_1399_store_0_ack_1 : boolean;
  signal ptr_deref_1407_base_resize_req_0 : boolean;
  signal ptr_deref_1407_base_resize_ack_0 : boolean;
  signal ptr_deref_1407_root_address_inst_req_0 : boolean;
  signal ptr_deref_1407_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1407_addr_0_req_0 : boolean;
  signal ptr_deref_1407_addr_0_ack_0 : boolean;
  signal ptr_deref_1407_addr_0_req_1 : boolean;
  signal ptr_deref_1407_addr_0_ack_1 : boolean;
  signal ptr_deref_1407_addr_1_req_0 : boolean;
  signal ptr_deref_1407_addr_1_ack_0 : boolean;
  signal ptr_deref_1407_addr_1_req_1 : boolean;
  signal ptr_deref_1407_addr_1_ack_1 : boolean;
  signal ptr_deref_1407_addr_2_req_0 : boolean;
  signal ptr_deref_1407_addr_2_ack_0 : boolean;
  signal ptr_deref_1407_addr_2_req_1 : boolean;
  signal ptr_deref_1407_addr_2_ack_1 : boolean;
  signal ptr_deref_1407_addr_3_req_0 : boolean;
  signal ptr_deref_1407_addr_3_ack_0 : boolean;
  signal ptr_deref_1407_addr_3_req_1 : boolean;
  signal ptr_deref_1407_addr_3_ack_1 : boolean;
  signal ptr_deref_1407_load_0_req_0 : boolean;
  signal ptr_deref_1407_load_0_ack_0 : boolean;
  signal ptr_deref_1407_load_1_req_0 : boolean;
  signal ptr_deref_1407_load_1_ack_0 : boolean;
  signal ptr_deref_1407_load_2_req_0 : boolean;
  signal ptr_deref_1407_load_2_ack_0 : boolean;
  signal ptr_deref_1407_load_3_req_0 : boolean;
  signal ptr_deref_1407_load_3_ack_0 : boolean;
  signal ptr_deref_1407_load_0_req_1 : boolean;
  signal ptr_deref_1407_load_0_ack_1 : boolean;
  signal ptr_deref_1407_load_1_req_1 : boolean;
  signal ptr_deref_1407_load_1_ack_1 : boolean;
  signal ptr_deref_1407_load_2_req_1 : boolean;
  signal ptr_deref_1407_load_2_ack_1 : boolean;
  signal ptr_deref_1407_load_3_req_1 : boolean;
  signal ptr_deref_1407_load_3_ack_1 : boolean;
  signal ptr_deref_1407_gather_scatter_req_0 : boolean;
  signal ptr_deref_1407_gather_scatter_ack_0 : boolean;
  signal binary_1413_inst_req_0 : boolean;
  signal binary_1413_inst_ack_0 : boolean;
  signal binary_1413_inst_req_1 : boolean;
  signal binary_1413_inst_ack_1 : boolean;
  signal ptr_deref_1416_base_resize_req_0 : boolean;
  signal ptr_deref_1416_base_resize_ack_0 : boolean;
  signal ptr_deref_1416_root_address_inst_req_0 : boolean;
  signal ptr_deref_1416_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1416_addr_0_req_0 : boolean;
  signal ptr_deref_1416_addr_0_ack_0 : boolean;
  signal ptr_deref_1416_addr_0_req_1 : boolean;
  signal ptr_deref_1416_addr_0_ack_1 : boolean;
  signal ptr_deref_1416_addr_1_req_0 : boolean;
  signal ptr_deref_1416_addr_1_ack_0 : boolean;
  signal ptr_deref_1416_addr_1_req_1 : boolean;
  signal ptr_deref_1416_addr_1_ack_1 : boolean;
  signal ptr_deref_1416_addr_2_req_0 : boolean;
  signal ptr_deref_1416_addr_2_ack_0 : boolean;
  signal ptr_deref_1416_addr_2_req_1 : boolean;
  signal ptr_deref_1416_addr_2_ack_1 : boolean;
  signal ptr_deref_1416_addr_3_req_0 : boolean;
  signal ptr_deref_1416_addr_3_ack_0 : boolean;
  signal ptr_deref_1416_addr_3_req_1 : boolean;
  signal ptr_deref_1416_addr_3_ack_1 : boolean;
  signal ptr_deref_1416_gather_scatter_req_0 : boolean;
  signal ptr_deref_1416_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1416_store_0_req_0 : boolean;
  signal ptr_deref_1416_store_0_ack_0 : boolean;
  signal ptr_deref_1416_store_1_req_0 : boolean;
  signal ptr_deref_1416_store_1_ack_0 : boolean;
  signal ptr_deref_1416_store_2_req_0 : boolean;
  signal ptr_deref_1416_store_2_ack_0 : boolean;
  signal ptr_deref_1416_store_3_req_0 : boolean;
  signal ptr_deref_1416_store_3_ack_0 : boolean;
  signal ptr_deref_1416_store_0_req_1 : boolean;
  signal ptr_deref_1416_store_0_ack_1 : boolean;
  signal ptr_deref_1416_store_1_req_1 : boolean;
  signal ptr_deref_1416_store_1_ack_1 : boolean;
  signal ptr_deref_1416_store_2_req_1 : boolean;
  signal ptr_deref_1416_store_2_ack_1 : boolean;
  signal ptr_deref_1416_store_3_req_1 : boolean;
  signal ptr_deref_1416_store_3_ack_1 : boolean;
  signal ptr_deref_1421_base_resize_req_0 : boolean;
  signal ptr_deref_1421_base_resize_ack_0 : boolean;
  signal ptr_deref_1421_root_address_inst_req_0 : boolean;
  signal ptr_deref_1421_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1421_addr_0_req_0 : boolean;
  signal ptr_deref_1421_addr_0_ack_0 : boolean;
  signal ptr_deref_1421_addr_0_req_1 : boolean;
  signal ptr_deref_1421_addr_0_ack_1 : boolean;
  signal ptr_deref_1421_addr_1_req_0 : boolean;
  signal ptr_deref_1421_addr_1_ack_0 : boolean;
  signal ptr_deref_1421_addr_1_req_1 : boolean;
  signal ptr_deref_1421_addr_1_ack_1 : boolean;
  signal ptr_deref_1421_addr_2_req_0 : boolean;
  signal ptr_deref_1421_addr_2_ack_0 : boolean;
  signal ptr_deref_1421_addr_2_req_1 : boolean;
  signal ptr_deref_1421_addr_2_ack_1 : boolean;
  signal ptr_deref_1421_addr_3_req_0 : boolean;
  signal ptr_deref_1421_addr_3_ack_0 : boolean;
  signal ptr_deref_1421_addr_3_req_1 : boolean;
  signal ptr_deref_1421_addr_3_ack_1 : boolean;
  signal ptr_deref_1421_load_0_req_0 : boolean;
  signal ptr_deref_1421_load_0_ack_0 : boolean;
  signal ptr_deref_1421_load_1_req_0 : boolean;
  signal ptr_deref_1421_load_1_ack_0 : boolean;
  signal ptr_deref_1421_load_2_req_0 : boolean;
  signal ptr_deref_1421_load_2_ack_0 : boolean;
  signal ptr_deref_1421_load_3_req_0 : boolean;
  signal ptr_deref_1421_load_3_ack_0 : boolean;
  signal ptr_deref_1421_load_0_req_1 : boolean;
  signal ptr_deref_1421_load_0_ack_1 : boolean;
  signal ptr_deref_1421_load_1_req_1 : boolean;
  signal ptr_deref_1421_load_1_ack_1 : boolean;
  signal ptr_deref_1421_load_2_req_1 : boolean;
  signal ptr_deref_1421_load_2_ack_1 : boolean;
  signal ptr_deref_1421_load_3_req_1 : boolean;
  signal ptr_deref_1421_load_3_ack_1 : boolean;
  signal ptr_deref_1421_gather_scatter_req_0 : boolean;
  signal ptr_deref_1421_gather_scatter_ack_0 : boolean;
  signal binary_1427_inst_req_0 : boolean;
  signal binary_1427_inst_ack_0 : boolean;
  signal binary_1427_inst_req_1 : boolean;
  signal binary_1427_inst_ack_1 : boolean;
  signal if_stmt_1429_branch_req_0 : boolean;
  signal if_stmt_1429_branch_ack_1 : boolean;
  signal if_stmt_1429_branch_ack_0 : boolean;
  signal ptr_deref_1438_base_resize_req_0 : boolean;
  signal ptr_deref_1438_base_resize_ack_0 : boolean;
  signal ptr_deref_1438_root_address_inst_req_0 : boolean;
  signal ptr_deref_1438_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1438_addr_0_req_0 : boolean;
  signal ptr_deref_1438_addr_0_ack_0 : boolean;
  signal ptr_deref_1438_addr_0_req_1 : boolean;
  signal ptr_deref_1438_addr_0_ack_1 : boolean;
  signal ptr_deref_1438_addr_1_req_0 : boolean;
  signal ptr_deref_1438_addr_1_ack_0 : boolean;
  signal ptr_deref_1438_addr_1_req_1 : boolean;
  signal ptr_deref_1438_addr_1_ack_1 : boolean;
  signal ptr_deref_1438_addr_2_req_0 : boolean;
  signal ptr_deref_1438_addr_2_ack_0 : boolean;
  signal ptr_deref_1438_addr_2_req_1 : boolean;
  signal ptr_deref_1438_addr_2_ack_1 : boolean;
  signal ptr_deref_1438_addr_3_req_0 : boolean;
  signal ptr_deref_1438_addr_3_ack_0 : boolean;
  signal ptr_deref_1438_addr_3_req_1 : boolean;
  signal ptr_deref_1438_addr_3_ack_1 : boolean;
  signal ptr_deref_1438_load_0_req_0 : boolean;
  signal ptr_deref_1438_load_0_ack_0 : boolean;
  signal ptr_deref_1438_load_1_req_0 : boolean;
  signal ptr_deref_1438_load_1_ack_0 : boolean;
  signal ptr_deref_1438_load_2_req_0 : boolean;
  signal ptr_deref_1438_load_2_ack_0 : boolean;
  signal ptr_deref_1438_load_3_req_0 : boolean;
  signal ptr_deref_1438_load_3_ack_0 : boolean;
  signal ptr_deref_1438_load_0_req_1 : boolean;
  signal ptr_deref_1438_load_0_ack_1 : boolean;
  signal ptr_deref_1438_load_1_req_1 : boolean;
  signal ptr_deref_1438_load_1_ack_1 : boolean;
  signal ptr_deref_1438_load_2_req_1 : boolean;
  signal ptr_deref_1438_load_2_ack_1 : boolean;
  signal ptr_deref_1438_load_3_req_1 : boolean;
  signal ptr_deref_1438_load_3_ack_1 : boolean;
  signal ptr_deref_1438_gather_scatter_req_0 : boolean;
  signal ptr_deref_1438_gather_scatter_ack_0 : boolean;
  signal if_stmt_1449_branch_req_0 : boolean;
  signal ptr_deref_1442_base_resize_req_0 : boolean;
  signal ptr_deref_1442_base_resize_ack_0 : boolean;
  signal ptr_deref_1442_root_address_inst_req_0 : boolean;
  signal ptr_deref_1442_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1442_addr_0_req_0 : boolean;
  signal ptr_deref_1442_addr_0_ack_0 : boolean;
  signal ptr_deref_1442_addr_0_req_1 : boolean;
  signal ptr_deref_1442_addr_0_ack_1 : boolean;
  signal ptr_deref_1442_addr_1_req_0 : boolean;
  signal ptr_deref_1442_addr_1_ack_0 : boolean;
  signal ptr_deref_1442_addr_1_req_1 : boolean;
  signal ptr_deref_1442_addr_1_ack_1 : boolean;
  signal ptr_deref_1442_addr_2_req_0 : boolean;
  signal ptr_deref_1442_addr_2_ack_0 : boolean;
  signal ptr_deref_1442_addr_2_req_1 : boolean;
  signal ptr_deref_1442_addr_2_ack_1 : boolean;
  signal ptr_deref_1442_addr_3_req_0 : boolean;
  signal ptr_deref_1442_addr_3_ack_0 : boolean;
  signal ptr_deref_1442_addr_3_req_1 : boolean;
  signal ptr_deref_1442_addr_3_ack_1 : boolean;
  signal ptr_deref_1442_load_0_req_0 : boolean;
  signal ptr_deref_1442_load_0_ack_0 : boolean;
  signal ptr_deref_1442_load_1_req_0 : boolean;
  signal ptr_deref_1442_load_1_ack_0 : boolean;
  signal ptr_deref_1442_load_2_req_0 : boolean;
  signal ptr_deref_1442_load_2_ack_0 : boolean;
  signal ptr_deref_1442_load_3_req_0 : boolean;
  signal ptr_deref_1442_load_3_ack_0 : boolean;
  signal ptr_deref_1442_load_0_req_1 : boolean;
  signal ptr_deref_1442_load_0_ack_1 : boolean;
  signal ptr_deref_1442_load_1_req_1 : boolean;
  signal ptr_deref_1442_load_1_ack_1 : boolean;
  signal ptr_deref_1442_load_2_req_1 : boolean;
  signal ptr_deref_1458_addr_0_req_0 : boolean;
  signal ptr_deref_1458_addr_0_ack_0 : boolean;
  signal ptr_deref_1458_addr_0_req_1 : boolean;
  signal ptr_deref_1458_addr_0_ack_1 : boolean;
  signal ptr_deref_1458_addr_1_req_0 : boolean;
  signal ptr_deref_1458_addr_1_ack_0 : boolean;
  signal ptr_deref_1458_addr_1_req_1 : boolean;
  signal ptr_deref_1458_addr_1_ack_1 : boolean;
  signal ptr_deref_1458_addr_2_req_0 : boolean;
  signal ptr_deref_1458_addr_2_ack_0 : boolean;
  signal ptr_deref_1458_addr_2_req_1 : boolean;
  signal ptr_deref_1458_addr_2_ack_1 : boolean;
  signal ptr_deref_1458_addr_3_req_0 : boolean;
  signal ptr_deref_1458_addr_3_ack_0 : boolean;
  signal ptr_deref_1458_addr_3_req_1 : boolean;
  signal ptr_deref_1458_addr_3_ack_1 : boolean;
  signal ptr_deref_1458_load_0_req_0 : boolean;
  signal ptr_deref_1458_load_0_ack_0 : boolean;
  signal ptr_deref_1458_load_1_req_0 : boolean;
  signal ptr_deref_1458_load_1_ack_0 : boolean;
  signal ptr_deref_1458_load_2_req_0 : boolean;
  signal ptr_deref_1458_load_2_ack_0 : boolean;
  signal ptr_deref_1458_load_3_req_0 : boolean;
  signal ptr_deref_1458_load_3_ack_0 : boolean;
  signal ptr_deref_1458_load_0_req_1 : boolean;
  signal ptr_deref_1458_load_0_ack_1 : boolean;
  signal ptr_deref_1458_load_1_req_1 : boolean;
  signal ptr_deref_1458_load_1_ack_1 : boolean;
  signal ptr_deref_1458_load_2_req_1 : boolean;
  signal ptr_deref_1458_load_2_ack_1 : boolean;
  signal ptr_deref_1458_load_3_req_1 : boolean;
  signal ptr_deref_1458_load_3_ack_1 : boolean;
  signal ptr_deref_1458_gather_scatter_req_0 : boolean;
  signal ptr_deref_1458_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1463_base_resize_req_0 : boolean;
  signal ptr_deref_1463_base_resize_ack_0 : boolean;
  signal ptr_deref_1463_root_address_inst_req_0 : boolean;
  signal ptr_deref_1463_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1463_addr_0_req_0 : boolean;
  signal ptr_deref_1463_addr_0_ack_0 : boolean;
  signal ptr_deref_1463_gather_scatter_req_0 : boolean;
  signal ptr_deref_1463_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1463_store_0_req_0 : boolean;
  signal ptr_deref_1463_store_0_ack_0 : boolean;
  signal ptr_deref_1463_store_0_req_1 : boolean;
  signal ptr_deref_1463_store_0_ack_1 : boolean;
  signal call_stmt_1470_call_req_0 : boolean;
  signal call_stmt_1470_call_ack_0 : boolean;
  signal call_stmt_1470_call_req_1 : boolean;
  signal call_stmt_1470_call_ack_1 : boolean;
  signal array_obj_ref_1477_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1477_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1477_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1477_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1477_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1477_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1477_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1477_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1477_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1477_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1477_offset_inst_req_0 : boolean;
  signal array_obj_ref_1477_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1477_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1477_root_address_inst_ack_0 : boolean;
  signal addr_of_1478_final_reg_req_0 : boolean;
  signal addr_of_1478_final_reg_ack_0 : boolean;
  signal ptr_deref_1482_base_resize_req_0 : boolean;
  signal ptr_deref_1482_base_resize_ack_0 : boolean;
  signal ptr_deref_1482_root_address_inst_req_0 : boolean;
  signal ptr_deref_1482_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1482_addr_0_req_0 : boolean;
  signal ptr_deref_1482_addr_0_ack_0 : boolean;
  signal ptr_deref_1482_load_0_req_0 : boolean;
  signal ptr_deref_1482_load_0_ack_0 : boolean;
  signal ptr_deref_1482_load_0_req_1 : boolean;
  signal ptr_deref_1482_load_0_ack_1 : boolean;
  signal ptr_deref_1482_gather_scatter_req_0 : boolean;
  signal ptr_deref_1482_gather_scatter_ack_0 : boolean;
  signal binary_1488_inst_req_0 : boolean;
  signal binary_1488_inst_ack_0 : boolean;
  signal binary_1488_inst_req_1 : boolean;
  signal binary_1488_inst_ack_1 : boolean;
  signal array_obj_ref_1496_index_2_resize_req_0 : boolean;
  signal array_obj_ref_1496_index_2_resize_ack_0 : boolean;
  signal array_obj_ref_1496_index_2_rename_req_0 : boolean;
  signal array_obj_ref_1496_index_2_rename_ack_0 : boolean;
  signal array_obj_ref_1496_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1496_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1496_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1496_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1496_offset_inst_req_0 : boolean;
  signal array_obj_ref_1496_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1496_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1496_root_address_inst_ack_0 : boolean;
  signal addr_of_1497_final_reg_req_0 : boolean;
  signal addr_of_1497_final_reg_ack_0 : boolean;
  signal ptr_deref_1501_base_resize_req_0 : boolean;
  signal ptr_deref_1501_base_resize_ack_0 : boolean;
  signal ptr_deref_1501_root_address_inst_req_0 : boolean;
  signal ptr_deref_1501_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1501_addr_0_req_0 : boolean;
  signal ptr_deref_1501_addr_0_ack_0 : boolean;
  signal ptr_deref_1501_load_0_req_0 : boolean;
  signal ptr_deref_1501_load_0_ack_0 : boolean;
  signal ptr_deref_1501_load_0_req_1 : boolean;
  signal ptr_deref_1501_load_0_ack_1 : boolean;
  signal ptr_deref_1501_gather_scatter_req_0 : boolean;
  signal ptr_deref_1501_gather_scatter_ack_0 : boolean;
  signal binary_1507_inst_req_0 : boolean;
  signal binary_1507_inst_ack_0 : boolean;
  signal binary_1507_inst_req_1 : boolean;
  signal binary_1507_inst_ack_1 : boolean;
  signal if_stmt_1509_branch_req_0 : boolean;
  signal if_stmt_1509_branch_ack_1 : boolean;
  signal if_stmt_1509_branch_ack_0 : boolean;
  signal binary_1520_inst_req_0 : boolean;
  signal binary_1520_inst_ack_0 : boolean;
  signal binary_1520_inst_req_1 : boolean;
  signal binary_1520_inst_ack_1 : boolean;
  signal array_obj_ref_1528_index_2_resize_req_0 : boolean;
  signal array_obj_ref_1528_index_2_resize_ack_0 : boolean;
  signal array_obj_ref_1528_index_2_rename_req_0 : boolean;
  signal array_obj_ref_1528_index_2_rename_ack_0 : boolean;
  signal array_obj_ref_1528_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1528_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1528_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1528_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1528_offset_inst_req_0 : boolean;
  signal array_obj_ref_1528_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1528_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1528_root_address_inst_ack_0 : boolean;
  signal addr_of_1529_final_reg_req_0 : boolean;
  signal addr_of_1529_final_reg_ack_0 : boolean;
  signal ptr_deref_1533_base_resize_req_0 : boolean;
  signal ptr_deref_1533_base_resize_ack_0 : boolean;
  signal ptr_deref_1533_root_address_inst_req_0 : boolean;
  signal ptr_deref_1533_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1533_addr_0_req_0 : boolean;
  signal ptr_deref_1533_addr_0_ack_0 : boolean;
  signal ptr_deref_1533_load_0_req_0 : boolean;
  signal ptr_deref_1533_load_0_ack_0 : boolean;
  signal ptr_deref_1533_load_0_req_1 : boolean;
  signal ptr_deref_1533_load_0_ack_1 : boolean;
  signal ptr_deref_1533_gather_scatter_req_0 : boolean;
  signal ptr_deref_1533_gather_scatter_ack_0 : boolean;
  signal binary_1539_inst_req_0 : boolean;
  signal binary_1539_inst_ack_0 : boolean;
  signal binary_1539_inst_req_1 : boolean;
  signal binary_1539_inst_ack_1 : boolean;
  signal if_stmt_1541_branch_req_0 : boolean;
  signal if_stmt_1541_branch_ack_1 : boolean;
  signal if_stmt_1541_branch_ack_0 : boolean;
  signal binary_1552_inst_req_0 : boolean;
  signal binary_1552_inst_ack_0 : boolean;
  signal binary_1552_inst_req_1 : boolean;
  signal binary_1552_inst_ack_1 : boolean;
  signal array_obj_ref_1560_index_2_resize_req_0 : boolean;
  signal array_obj_ref_1560_index_2_resize_ack_0 : boolean;
  signal array_obj_ref_1560_index_2_rename_req_0 : boolean;
  signal array_obj_ref_1560_index_2_rename_ack_0 : boolean;
  signal array_obj_ref_1560_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1560_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1560_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1560_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1560_offset_inst_req_0 : boolean;
  signal array_obj_ref_1560_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1560_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1560_root_address_inst_ack_0 : boolean;
  signal addr_of_1561_final_reg_req_0 : boolean;
  signal addr_of_1561_final_reg_ack_0 : boolean;
  signal ptr_deref_1565_base_resize_req_0 : boolean;
  signal ptr_deref_1565_base_resize_ack_0 : boolean;
  signal ptr_deref_1565_root_address_inst_req_0 : boolean;
  signal ptr_deref_1565_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1565_addr_0_req_0 : boolean;
  signal ptr_deref_1565_addr_0_ack_0 : boolean;
  signal ptr_deref_1565_load_0_req_0 : boolean;
  signal ptr_deref_1565_load_0_ack_0 : boolean;
  signal ptr_deref_1565_load_0_req_1 : boolean;
  signal ptr_deref_1565_load_0_ack_1 : boolean;
  signal ptr_deref_1565_gather_scatter_req_0 : boolean;
  signal ptr_deref_1565_gather_scatter_ack_0 : boolean;
  signal type_cast_1570_inst_req_0 : boolean;
  signal type_cast_1570_inst_ack_0 : boolean;
  signal binary_1574_inst_req_0 : boolean;
  signal binary_1574_inst_ack_0 : boolean;
  signal binary_1574_inst_req_1 : boolean;
  signal binary_1574_inst_ack_1 : boolean;
  signal if_stmt_1576_branch_req_0 : boolean;
  signal if_stmt_1576_branch_ack_1 : boolean;
  signal if_stmt_1576_branch_ack_0 : boolean;
  signal type_cast_1585_inst_req_0 : boolean;
  signal type_cast_1585_inst_ack_0 : boolean;
  signal binary_1589_inst_req_0 : boolean;
  signal binary_1589_inst_ack_0 : boolean;
  signal binary_1589_inst_req_1 : boolean;
  signal binary_1589_inst_ack_1 : boolean;
  signal if_stmt_1591_branch_req_0 : boolean;
  signal if_stmt_1591_branch_ack_1 : boolean;
  signal if_stmt_1591_branch_ack_0 : boolean;
  signal binary_1602_inst_req_0 : boolean;
  signal binary_1602_inst_ack_0 : boolean;
  signal binary_1602_inst_req_1 : boolean;
  signal binary_1602_inst_ack_1 : boolean;
  signal if_stmt_1604_branch_req_0 : boolean;
  signal if_stmt_1604_branch_ack_1 : boolean;
  signal if_stmt_1604_branch_ack_0 : boolean;
  signal binary_1615_inst_req_0 : boolean;
  signal binary_1615_inst_ack_0 : boolean;
  signal binary_1615_inst_req_1 : boolean;
  signal binary_1615_inst_ack_1 : boolean;
  signal if_stmt_1617_branch_req_0 : boolean;
  signal if_stmt_1617_branch_ack_1 : boolean;
  signal if_stmt_1617_branch_ack_0 : boolean;
  signal type_cast_1626_inst_req_0 : boolean;
  signal type_cast_1626_inst_ack_0 : boolean;
  signal binary_1630_inst_req_0 : boolean;
  signal binary_1630_inst_ack_0 : boolean;
  signal binary_1630_inst_req_1 : boolean;
  signal binary_1630_inst_ack_1 : boolean;
  signal if_stmt_1632_branch_req_0 : boolean;
  signal if_stmt_1632_branch_ack_1 : boolean;
  signal if_stmt_1632_branch_ack_0 : boolean;
  signal binary_1643_inst_req_0 : boolean;
  signal binary_1643_inst_ack_0 : boolean;
  signal binary_1643_inst_req_1 : boolean;
  signal binary_1643_inst_ack_1 : boolean;
  signal if_stmt_1645_branch_req_0 : boolean;
  signal if_stmt_1645_branch_ack_1 : boolean;
  signal if_stmt_1645_branch_ack_0 : boolean;
  signal binary_1656_inst_req_0 : boolean;
  signal binary_1656_inst_ack_0 : boolean;
  signal binary_1656_inst_req_1 : boolean;
  signal binary_1656_inst_ack_1 : boolean;
  signal if_stmt_1658_branch_req_0 : boolean;
  signal if_stmt_1658_branch_ack_1 : boolean;
  signal if_stmt_1658_branch_ack_0 : boolean;
  signal type_cast_1667_inst_req_0 : boolean;
  signal type_cast_1667_inst_ack_0 : boolean;
  signal simple_obj_ref_1665_inst_req_0 : boolean;
  signal simple_obj_ref_1665_inst_ack_0 : boolean;
  signal type_cast_1673_inst_req_0 : boolean;
  signal type_cast_1673_inst_ack_0 : boolean;
  signal simple_obj_ref_1671_inst_req_0 : boolean;
  signal simple_obj_ref_1671_inst_ack_0 : boolean;
  signal type_cast_1679_inst_req_0 : boolean;
  signal type_cast_1679_inst_ack_0 : boolean;
  signal simple_obj_ref_1677_inst_req_0 : boolean;
  signal simple_obj_ref_1677_inst_ack_0 : boolean;
  signal type_cast_1685_inst_req_0 : boolean;
  signal type_cast_1685_inst_ack_0 : boolean;
  signal simple_obj_ref_1683_inst_req_0 : boolean;
  signal simple_obj_ref_1683_inst_ack_0 : boolean;
  signal type_cast_1691_inst_req_0 : boolean;
  signal type_cast_1691_inst_ack_0 : boolean;
  signal simple_obj_ref_1689_inst_req_0 : boolean;
  signal simple_obj_ref_1689_inst_ack_0 : boolean;
  signal phi_stmt_1174_req_1 : boolean;
  signal type_cast_1177_inst_req_0 : boolean;
  signal type_cast_1177_inst_ack_0 : boolean;
  signal phi_stmt_1174_req_0 : boolean;
  signal phi_stmt_1174_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_rtt_CP_4152: Block -- control-path 
    signal cp_elements: BooleanArray(1054 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1054);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(1054), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(140) & cp_elements(976));
    cp_elements(2) <= OrReduce(cp_elements(138) & cp_elements(982));
    cp_elements(3) <= OrReduce(cp_elements(984) & cp_elements(986));
    cp_elements(4) <= cp_elements(207);
    cp_elements(5) <= OrReduce(cp_elements(214) & cp_elements(988));
    cp_elements(6) <= cp_elements(1003);
    cp_elements(7) <= OrReduce(cp_elements(247) & cp_elements(1005));
    cp_elements(8) <= OrReduce(cp_elements(278) & cp_elements(1018));
    cp_elements(9) <= OrReduce(cp_elements(293) & cp_elements(1020));
    cp_elements(10) <= cp_elements(430);
    cp_elements(11) <= OrReduce(cp_elements(439) & cp_elements(1022));
    cp_elements(12) <= cp_elements(573);
    cp_elements(13) <= OrReduce(cp_elements(580) & cp_elements(1026));
    cpelement_group_14 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(668) & cp_elements(1028));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(14),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(15) <= OrReduce(cp_elements(771) & cp_elements(1034));
    cp_elements(16) <= OrReduce(cp_elements(807) & cp_elements(1036));
    cp_elements(17) <= OrReduce(cp_elements(848) & cp_elements(1038));
    cp_elements(18) <= OrReduce(cp_elements(866) & cp_elements(1040));
    cp_elements(19) <= OrReduce(cp_elements(864) & cp_elements(1042));
    cp_elements(20) <= OrReduce(cp_elements(846) & cp_elements(1044));
    cp_elements(21) <= OrReduce(cp_elements(914) & cp_elements(1046));
    cp_elements(22) <= OrReduce(cp_elements(912) & cp_elements(1048));
    cp_elements(23) <= OrReduce(cp_elements(942) & cp_elements(1050));
    cp_elements(24) <= cp_elements(0);
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(26) & cp_elements(28));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => type_cast_1094_inst_req_0); -- 
    cp_elements(26) <= cp_elements(24);
    cp_elements(27) <= cp_elements(24);
    req_4341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => simple_obj_ref_1093_inst_req_0); -- 
    ack_4342_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1093_inst_ack_0, ack => cp_elements(28)); -- 
    ack_4347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1094_inst_ack_0, ack => cp_elements(29)); -- 
    cp_elements(30) <= cp_elements(29);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(33));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => type_cast_1098_inst_req_0); -- 
    cp_elements(32) <= cp_elements(30);
    cp_elements(33) <= cp_elements(30);
    ack_4360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_0, ack => cp_elements(34)); -- 
    base_resize_req_4371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_1105_base_resize_req_0); -- 
    cp_elements(35) <= cp_elements(30);
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_1105_final_reg_req_0); -- 
    base_resize_ack_4372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_base_resize_ack_0, ack => cp_elements(37)); -- 
    plus_base_rr_4377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_1105_root_address_inst_req_0); -- 
    plus_base_ra_4378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_root_address_inst_ack_0, ack => cp_elements(38)); -- 
    plus_base_cr_4379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_1105_root_address_inst_req_1); -- 
    plus_base_ca_4380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_root_address_inst_ack_1, ack => cp_elements(39)); -- 
    final_reg_ack_4385_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_final_reg_ack_0, ack => cp_elements(40)); -- 
    cpelement_group_41 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(40) & cp_elements(42));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(41),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => type_cast_1109_inst_req_0); -- 
    cp_elements(42) <= cp_elements(30);
    cp_elements(43) <= type_cast_1109_inst_ack_0;
    cpelement_group_44 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(43) & cp_elements(60));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(44),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(45) <= cp_elements(43);
    base_resize_req_4408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_1113_base_resize_req_0); -- 
    base_resize_ack_4409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_base_resize_ack_0, ack => cp_elements(46)); -- 
    sum_rename_req_4413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_1113_root_address_inst_req_0); -- 
    cp_elements(47) <= ptr_deref_1113_root_address_inst_ack_0;
    cp_elements(48) <= cp_elements(47);
    rr_4421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_1113_addr_0_req_0); -- 
    ra_4422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_0_ack_0, ack => cp_elements(49)); -- 
    cr_4423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_1113_addr_0_req_1); -- 
    ca_4424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_0_ack_1, ack => cp_elements(50)); -- 
    cp_elements(51) <= cp_elements(47);
    rr_4428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => ptr_deref_1113_addr_1_req_0); -- 
    ra_4429_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_1_ack_0, ack => cp_elements(52)); -- 
    cr_4430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => ptr_deref_1113_addr_1_req_1); -- 
    ca_4431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_1_ack_1, ack => cp_elements(53)); -- 
    cp_elements(54) <= cp_elements(47);
    rr_4435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_1113_addr_2_req_0); -- 
    ra_4436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_2_ack_0, ack => cp_elements(55)); -- 
    cr_4437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => ptr_deref_1113_addr_2_req_1); -- 
    ca_4438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_2_ack_1, ack => cp_elements(56)); -- 
    cp_elements(57) <= cp_elements(47);
    rr_4442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => ptr_deref_1113_addr_3_req_0); -- 
    ra_4443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_3_ack_0, ack => cp_elements(58)); -- 
    cr_4444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_1113_addr_3_req_1); -- 
    ca_4445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_3_ack_1, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(53) & cp_elements(56) & cp_elements(59));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(61) <= cp_elements(44);
    rr_4455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_1113_load_0_req_0); -- 
    ra_4456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_0_ack_0, ack => cp_elements(62)); -- 
    cp_elements(63) <= cp_elements(44);
    rr_4460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_1113_load_1_req_0); -- 
    ra_4461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_1_ack_0, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(44);
    rr_4465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_1113_load_2_req_0); -- 
    ra_4466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_2_ack_0, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(44);
    rr_4470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => ptr_deref_1113_load_3_req_0); -- 
    ra_4471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_3_ack_0, ack => cp_elements(68)); -- 
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(62) & cp_elements(64) & cp_elements(66) & cp_elements(68));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(70) <= cp_elements(69);
    cr_4481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_1113_load_0_req_1); -- 
    ca_4482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_0_ack_1, ack => cp_elements(71)); -- 
    cp_elements(72) <= cp_elements(69);
    cr_4486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_1113_load_1_req_1); -- 
    ca_4487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_1_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= cp_elements(69);
    cr_4491_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_1113_load_2_req_1); -- 
    ca_4492_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_2_ack_1, ack => cp_elements(75)); -- 
    cp_elements(76) <= cp_elements(69);
    cr_4496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_1113_load_3_req_1); -- 
    ca_4497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_3_ack_1, ack => cp_elements(77)); -- 
    cpelement_group_78 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(73) & cp_elements(75) & cp_elements(77));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(78),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_4498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => ptr_deref_1113_gather_scatter_req_0); -- 
    merge_ack_4499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_gather_scatter_ack_0, ack => cp_elements(79)); -- 
    phi_stmt_1174_req_7304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => phi_stmt_1174_req_1); -- 
    cp_elements(80) <= cp_elements(162);
    cpelement_group_81 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(81),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4542_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => addr_of_1124_final_reg_req_0); -- 
    cp_elements(82) <= cp_elements(80);
    cp_elements(83) <= cp_elements(80);
    index_resize_req_4516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => array_obj_ref_1123_index_0_resize_req_0); -- 
    index_resize_ack_4517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_index_0_resize_ack_0, ack => cp_elements(84)); -- 
    scale_rr_4521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => array_obj_ref_1123_index_0_scale_req_0); -- 
    scale_ra_4522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_index_0_scale_ack_0, ack => cp_elements(85)); -- 
    scale_cr_4523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => array_obj_ref_1123_index_0_scale_req_1); -- 
    scale_ca_4524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_index_0_scale_ack_1, ack => cp_elements(86)); -- 
    partial_sum_1_rr_4528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => array_obj_ref_1123_index_sum_1_req_0); -- 
    partial_sum_1_ra_4529_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_index_sum_1_ack_0, ack => cp_elements(87)); -- 
    partial_sum_1_cr_4530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => array_obj_ref_1123_index_sum_1_req_1); -- 
    partial_sum_1_ca_4531_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_index_sum_1_ack_1, ack => cp_elements(88)); -- 
    final_index_req_4532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => array_obj_ref_1123_offset_inst_req_0); -- 
    final_index_ack_4533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_offset_inst_ack_0, ack => cp_elements(89)); -- 
    sum_rename_req_4537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => array_obj_ref_1123_root_address_inst_req_0); -- 
    sum_rename_ack_4538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1123_root_address_inst_ack_0, ack => cp_elements(90)); -- 
    cp_elements(91) <= addr_of_1124_final_reg_ack_0;
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(101));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => addr_of_1133_final_reg_req_0); -- 
    cp_elements(93) <= cp_elements(80);
    cp_elements(94) <= cp_elements(80);
    index_resize_req_4557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => array_obj_ref_1132_index_0_resize_req_0); -- 
    index_resize_ack_4558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_index_0_resize_ack_0, ack => cp_elements(95)); -- 
    scale_rr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_1132_index_0_scale_req_0); -- 
    scale_ra_4563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_index_0_scale_ack_0, ack => cp_elements(96)); -- 
    scale_cr_4564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => array_obj_ref_1132_index_0_scale_req_1); -- 
    scale_ca_4565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_index_0_scale_ack_1, ack => cp_elements(97)); -- 
    partial_sum_1_rr_4569_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => array_obj_ref_1132_index_sum_1_req_0); -- 
    partial_sum_1_ra_4570_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_index_sum_1_ack_0, ack => cp_elements(98)); -- 
    partial_sum_1_cr_4571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_1132_index_sum_1_req_1); -- 
    partial_sum_1_ca_4572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_index_sum_1_ack_1, ack => cp_elements(99)); -- 
    final_index_req_4573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => array_obj_ref_1132_offset_inst_req_0); -- 
    final_index_ack_4574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_offset_inst_ack_0, ack => cp_elements(100)); -- 
    sum_rename_req_4578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => array_obj_ref_1132_root_address_inst_req_0); -- 
    sum_rename_ack_4579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_root_address_inst_ack_0, ack => cp_elements(101)); -- 
    cp_elements(102) <= addr_of_1133_final_reg_ack_0;
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(107));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_1137_load_0_req_0); -- 
    cp_elements(104) <= cp_elements(91);
    base_resize_req_4597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_1137_base_resize_req_0); -- 
    base_resize_ack_4598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1137_base_resize_ack_0, ack => cp_elements(105)); -- 
    sum_rename_req_4602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_1137_root_address_inst_req_0); -- 
    sum_rename_ack_4603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1137_root_address_inst_ack_0, ack => cp_elements(106)); -- 
    root_rename_req_4607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_1137_addr_0_req_0); -- 
    root_rename_ack_4608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1137_addr_0_ack_0, ack => cp_elements(107)); -- 
    ra_4619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1137_load_0_ack_0, ack => cp_elements(108)); -- 
    cr_4629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => ptr_deref_1137_load_0_req_1); -- 
    ca_4630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1137_load_0_ack_1, ack => cp_elements(109)); -- 
    merge_req_4631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_1137_gather_scatter_req_0); -- 
    merge_ack_4632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1137_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(115));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_1141_load_0_req_0); -- 
    cp_elements(112) <= cp_elements(102);
    base_resize_req_4645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => ptr_deref_1141_base_resize_req_0); -- 
    base_resize_ack_4646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_base_resize_ack_0, ack => cp_elements(113)); -- 
    sum_rename_req_4650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_1141_root_address_inst_req_0); -- 
    sum_rename_ack_4651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_root_address_inst_ack_0, ack => cp_elements(114)); -- 
    root_rename_req_4655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => ptr_deref_1141_addr_0_req_0); -- 
    root_rename_ack_4656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_addr_0_ack_0, ack => cp_elements(115)); -- 
    ra_4667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_load_0_ack_0, ack => cp_elements(116)); -- 
    cr_4677_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => ptr_deref_1141_load_0_req_1); -- 
    ca_4678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_load_0_ack_1, ack => cp_elements(117)); -- 
    merge_req_4679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_1141_gather_scatter_req_0); -- 
    merge_ack_4680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_gather_scatter_ack_0, ack => cp_elements(118)); -- 
    cpelement_group_119 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(120) & cp_elements(121));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => binary_1146_inst_req_0); -- 
    cp_elements(120) <= cp_elements(80);
    cp_elements(121) <= cp_elements(80);
    ra_4691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1146_inst_ack_0, ack => cp_elements(122)); -- 
    cr_4692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => binary_1146_inst_req_1); -- 
    ca_4693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1146_inst_ack_1, ack => cp_elements(123)); -- 
    cpelement_group_124 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(123) & cp_elements(125));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(124),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => binary_1151_inst_req_0); -- 
    cp_elements(125) <= cp_elements(80);
    ra_4704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1151_inst_ack_0, ack => cp_elements(126)); -- 
    cr_4705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => binary_1151_inst_req_1); -- 
    ca_4706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1151_inst_ack_1, ack => cp_elements(127)); -- 
    cpelement_group_128 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(129));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(128),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4715_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => binary_1157_inst_req_0); -- 
    cp_elements(129) <= cp_elements(80);
    ra_4716_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1157_inst_ack_0, ack => cp_elements(130)); -- 
    cr_4717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => binary_1157_inst_req_1); -- 
    ca_4718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1157_inst_ack_1, ack => cp_elements(131)); -- 
    cp_elements(132) <= cp_elements(131);
    cp_elements(133) <= false;
    cp_elements(134) <= cp_elements(133);
    cp_elements(135) <= cp_elements(131);
    branch_req_4726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => if_stmt_1159_branch_req_0); -- 
    cp_elements(136) <= cp_elements(135);
    cp_elements(137) <= cp_elements(136);
    if_choice_transition_4731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1159_branch_ack_1, ack => cp_elements(138)); -- 
    cp_elements(139) <= cp_elements(136);
    else_choice_transition_4735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1159_branch_ack_0, ack => cp_elements(140)); -- 
    cp_elements(141) <= cp_elements(1);
    cpelement_group_142 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(144));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(142),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => binary_1170_inst_req_0); -- 
    cp_elements(143) <= cp_elements(141);
    cp_elements(144) <= cp_elements(141);
    ra_4750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1170_inst_ack_0, ack => cp_elements(145)); -- 
    cr_4751_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => binary_1170_inst_req_1); -- 
    ca_4752_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1170_inst_ack_1, ack => cp_elements(146)); -- 
    req_7317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(146), ack => type_cast_1177_inst_req_0); -- 
    cp_elements(147) <= cp_elements(980);
    cpelement_group_148 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(153));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(148),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => binary_1188_inst_req_0); -- 
    cp_elements(149) <= cp_elements(147);
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(151) & cp_elements(152));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(150), ack => type_cast_1184_inst_req_0); -- 
    cp_elements(151) <= cp_elements(147);
    cp_elements(152) <= cp_elements(147);
    ack_4767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1184_inst_ack_0, ack => cp_elements(153)); -- 
    ra_4772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1188_inst_ack_0, ack => cp_elements(154)); -- 
    cr_4773_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => binary_1188_inst_req_1); -- 
    ca_4774_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1188_inst_ack_1, ack => cp_elements(155)); -- 
    cp_elements(156) <= cp_elements(155);
    cp_elements(157) <= false;
    cp_elements(158) <= cp_elements(157);
    cp_elements(159) <= cp_elements(155);
    branch_req_4782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(159), ack => if_stmt_1190_branch_req_0); -- 
    cp_elements(160) <= cp_elements(159);
    cp_elements(161) <= cp_elements(160);
    if_choice_transition_4787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1190_branch_ack_1, ack => cp_elements(162)); -- 
    cp_elements(163) <= cp_elements(160);
    else_choice_transition_4791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1190_branch_ack_0, ack => cp_elements(164)); -- 
    cp_elements(165) <= cp_elements(2);
    cpelement_group_166 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(167) & cp_elements(171));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => binary_1203_inst_req_0); -- 
    cp_elements(167) <= cp_elements(165);
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => type_cast_1199_inst_req_0); -- 
    cp_elements(169) <= cp_elements(165);
    cp_elements(170) <= cp_elements(165);
    ack_4808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_0, ack => cp_elements(171)); -- 
    ra_4813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1203_inst_ack_0, ack => cp_elements(172)); -- 
    cr_4814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(172), ack => binary_1203_inst_req_1); -- 
    ca_4815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1203_inst_ack_1, ack => cp_elements(173)); -- 
    cp_elements(174) <= cp_elements(173);
    cp_elements(175) <= false;
    cp_elements(176) <= cp_elements(175);
    cp_elements(177) <= cp_elements(173);
    branch_req_4823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => if_stmt_1205_branch_req_0); -- 
    cp_elements(178) <= cp_elements(177);
    cp_elements(179) <= cp_elements(178);
    if_choice_transition_4828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1205_branch_ack_1, ack => cp_elements(180)); -- 
    cp_elements(181) <= cp_elements(178);
    else_choice_transition_4832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1205_branch_ack_0, ack => cp_elements(182)); -- 
    cp_elements(183) <= cp_elements(3);
    cp_elements(184) <= cp_elements(183);
    rr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(184), ack => simple_obj_ref_1213_load_0_req_0); -- 
    cp_elements(185) <= simple_obj_ref_1213_load_0_ack_0;
    cp_elements(186) <= cp_elements(185);
    cr_4864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => simple_obj_ref_1213_load_0_req_1); -- 
    ca_4865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1213_load_0_ack_1, ack => cp_elements(187)); -- 
    merge_req_4866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => simple_obj_ref_1213_gather_scatter_req_0); -- 
    merge_ack_4867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1213_gather_scatter_ack_0, ack => cp_elements(188)); -- 
    cpelement_group_189 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(188) & cp_elements(190));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(189),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => binary_1219_inst_req_0); -- 
    cp_elements(190) <= cp_elements(183);
    ra_4877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1219_inst_ack_0, ack => cp_elements(191)); -- 
    cr_4878_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => binary_1219_inst_req_1); -- 
    cp_elements(192) <= binary_1219_inst_ack_1;
    cp_elements(193) <= cp_elements(192);
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(185) & cp_elements(193) & cp_elements(195));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_4890_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => simple_obj_ref_1221_gather_scatter_req_0); -- 
    cp_elements(195) <= cp_elements(183);
    split_ack_4891_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1221_gather_scatter_ack_0, ack => cp_elements(196)); -- 
    rr_4898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => simple_obj_ref_1221_store_0_req_0); -- 
    ra_4899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1221_store_0_ack_0, ack => cp_elements(197)); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => simple_obj_ref_1221_store_0_req_1); -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1221_store_0_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(200) & cp_elements(204));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => binary_1230_inst_req_0); -- 
    cp_elements(200) <= cp_elements(183);
    cpelement_group_201 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(202) & cp_elements(203));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(201),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4921_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => type_cast_1226_inst_req_0); -- 
    cp_elements(202) <= cp_elements(183);
    cp_elements(203) <= cp_elements(192);
    ack_4922_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_0, ack => cp_elements(204)); -- 
    ra_4927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1230_inst_ack_0, ack => cp_elements(205)); -- 
    cr_4928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => binary_1230_inst_req_1); -- 
    ca_4929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1230_inst_ack_1, ack => cp_elements(206)); -- 
    cpelement_group_207 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(198) & cp_elements(206));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(207),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(208) <= cp_elements(4);
    cp_elements(209) <= false;
    cp_elements(210) <= cp_elements(209);
    cp_elements(211) <= cp_elements(4);
    branch_req_4937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => if_stmt_1232_branch_req_0); -- 
    cp_elements(212) <= cp_elements(211);
    cp_elements(213) <= cp_elements(212);
    if_choice_transition_4942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1232_branch_ack_1, ack => cp_elements(214)); -- 
    cp_elements(215) <= cp_elements(212);
    else_choice_transition_4946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1232_branch_ack_0, ack => cp_elements(216)); -- 
    cp_elements(217) <= cp_elements(6);
    cpelement_group_218 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(219) & cp_elements(227));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(218),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(218), ack => addr_of_1261_final_reg_req_0); -- 
    cp_elements(219) <= cp_elements(217);
    cp_elements(220) <= cp_elements(217);
    index_resize_req_4965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(220), ack => array_obj_ref_1260_index_0_resize_req_0); -- 
    index_resize_ack_4966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_0_resize_ack_0, ack => cp_elements(221)); -- 
    scale_rr_4970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => array_obj_ref_1260_index_0_scale_req_0); -- 
    scale_ra_4971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_0_scale_ack_0, ack => cp_elements(222)); -- 
    scale_cr_4972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => array_obj_ref_1260_index_0_scale_req_1); -- 
    scale_ca_4973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_0_scale_ack_1, ack => cp_elements(223)); -- 
    partial_sum_1_rr_4977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => array_obj_ref_1260_index_sum_1_req_0); -- 
    partial_sum_1_ra_4978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_sum_1_ack_0, ack => cp_elements(224)); -- 
    partial_sum_1_cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => array_obj_ref_1260_index_sum_1_req_1); -- 
    partial_sum_1_ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_sum_1_ack_1, ack => cp_elements(225)); -- 
    final_index_req_4981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => array_obj_ref_1260_offset_inst_req_0); -- 
    final_index_ack_4982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_offset_inst_ack_0, ack => cp_elements(226)); -- 
    sum_rename_req_4986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => array_obj_ref_1260_root_address_inst_req_0); -- 
    sum_rename_ack_4987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_root_address_inst_ack_0, ack => cp_elements(227)); -- 
    cp_elements(228) <= addr_of_1261_final_reg_ack_0;
    cpelement_group_229 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(228) & cp_elements(233));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(229),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => ptr_deref_1265_load_0_req_0); -- 
    cp_elements(230) <= cp_elements(228);
    base_resize_req_5005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => ptr_deref_1265_base_resize_req_0); -- 
    base_resize_ack_5006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_base_resize_ack_0, ack => cp_elements(231)); -- 
    sum_rename_req_5010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_1265_root_address_inst_req_0); -- 
    sum_rename_ack_5011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_root_address_inst_ack_0, ack => cp_elements(232)); -- 
    root_rename_req_5015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(232), ack => ptr_deref_1265_addr_0_req_0); -- 
    root_rename_ack_5016_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_addr_0_ack_0, ack => cp_elements(233)); -- 
    ra_5027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_load_0_ack_0, ack => cp_elements(234)); -- 
    cr_5037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_1265_load_0_req_1); -- 
    ca_5038_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_load_0_ack_1, ack => cp_elements(235)); -- 
    merge_req_5039_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => ptr_deref_1265_gather_scatter_req_0); -- 
    merge_ack_5040_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_gather_scatter_ack_0, ack => cp_elements(236)); -- 
    cpelement_group_237 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(236) & cp_elements(238));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(237),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => binary_1271_inst_req_0); -- 
    cp_elements(238) <= cp_elements(217);
    ra_5050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1271_inst_ack_0, ack => cp_elements(239)); -- 
    cr_5051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => binary_1271_inst_req_1); -- 
    ca_5052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1271_inst_ack_1, ack => cp_elements(240)); -- 
    cp_elements(241) <= cp_elements(240);
    cp_elements(242) <= false;
    cp_elements(243) <= cp_elements(242);
    cp_elements(244) <= cp_elements(240);
    branch_req_5060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => if_stmt_1273_branch_req_0); -- 
    cp_elements(245) <= cp_elements(244);
    cp_elements(246) <= cp_elements(245);
    if_choice_transition_5065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1273_branch_ack_1, ack => cp_elements(247)); -- 
    cp_elements(248) <= cp_elements(245);
    cp_elements(249) <= if_stmt_1273_branch_ack_0;
    cp_elements(250) <= cp_elements(7);
    cpelement_group_251 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(252) & cp_elements(260));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(251),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => addr_of_1285_final_reg_req_0); -- 
    cp_elements(252) <= cp_elements(250);
    cp_elements(253) <= cp_elements(250);
    index_resize_req_5088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(253), ack => array_obj_ref_1284_index_0_resize_req_0); -- 
    index_resize_ack_5089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_index_0_resize_ack_0, ack => cp_elements(254)); -- 
    scale_rr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(254), ack => array_obj_ref_1284_index_0_scale_req_0); -- 
    scale_ra_5094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_index_0_scale_ack_0, ack => cp_elements(255)); -- 
    scale_cr_5095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => array_obj_ref_1284_index_0_scale_req_1); -- 
    scale_ca_5096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_index_0_scale_ack_1, ack => cp_elements(256)); -- 
    partial_sum_1_rr_5100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => array_obj_ref_1284_index_sum_1_req_0); -- 
    partial_sum_1_ra_5101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_index_sum_1_ack_0, ack => cp_elements(257)); -- 
    partial_sum_1_cr_5102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => array_obj_ref_1284_index_sum_1_req_1); -- 
    partial_sum_1_ca_5103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_index_sum_1_ack_1, ack => cp_elements(258)); -- 
    final_index_req_5104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => array_obj_ref_1284_offset_inst_req_0); -- 
    final_index_ack_5105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_offset_inst_ack_0, ack => cp_elements(259)); -- 
    sum_rename_req_5109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => array_obj_ref_1284_root_address_inst_req_0); -- 
    sum_rename_ack_5110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1284_root_address_inst_ack_0, ack => cp_elements(260)); -- 
    cp_elements(261) <= addr_of_1285_final_reg_ack_0;
    cp_elements(262) <= cp_elements(1016);
    cpelement_group_263 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(264) & cp_elements(265));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(263),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => binary_1300_inst_req_0); -- 
    cp_elements(264) <= cp_elements(262);
    cp_elements(265) <= cp_elements(262);
    ra_5128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1300_inst_ack_0, ack => cp_elements(266)); -- 
    cr_5129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => binary_1300_inst_req_1); -- 
    ca_5130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1300_inst_ack_1, ack => cp_elements(267)); -- 
    cpelement_group_268 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(267) & cp_elements(269));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(268),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => binary_1306_inst_req_0); -- 
    cp_elements(269) <= cp_elements(262);
    ra_5140_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1306_inst_ack_0, ack => cp_elements(270)); -- 
    cr_5141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => binary_1306_inst_req_1); -- 
    ca_5142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1306_inst_ack_1, ack => cp_elements(271)); -- 
    cp_elements(272) <= cp_elements(271);
    cp_elements(273) <= false;
    cp_elements(274) <= cp_elements(273);
    cp_elements(275) <= cp_elements(271);
    branch_req_5150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => if_stmt_1308_branch_req_0); -- 
    cp_elements(276) <= cp_elements(275);
    cp_elements(277) <= cp_elements(276);
    if_choice_transition_5155_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1308_branch_ack_1, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(276);
    else_choice_transition_5159_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1308_branch_ack_0, ack => cp_elements(280)); -- 
    cp_elements(281) <= cp_elements(8);
    cpelement_group_282 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(284));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(282),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => binary_1319_inst_req_0); -- 
    cp_elements(283) <= cp_elements(281);
    cp_elements(284) <= cp_elements(281);
    ra_5174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1319_inst_ack_0, ack => cp_elements(285)); -- 
    cr_5175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(285), ack => binary_1319_inst_req_1); -- 
    ca_5176_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1319_inst_ack_1, ack => cp_elements(286)); -- 
    cp_elements(287) <= cp_elements(286);
    cp_elements(288) <= false;
    cp_elements(289) <= cp_elements(288);
    cp_elements(290) <= cp_elements(286);
    branch_req_5184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => if_stmt_1321_branch_req_0); -- 
    cp_elements(291) <= cp_elements(290);
    cp_elements(292) <= cp_elements(291);
    if_choice_transition_5189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1321_branch_ack_1, ack => cp_elements(293)); -- 
    cp_elements(294) <= cp_elements(291);
    else_choice_transition_5193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1321_branch_ack_0, ack => cp_elements(295)); -- 
    cp_elements(296) <= cp_elements(295);
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(297) & cp_elements(305));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5229_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => array_obj_ref_1333_final_reg_req_0); -- 
    cp_elements(299) <= cp_elements(296);
    base_resize_req_5216_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(299), ack => array_obj_ref_1333_base_resize_req_0); -- 
    cp_elements(300) <= cp_elements(296);
    final_index_req_5210_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => array_obj_ref_1333_offset_inst_req_0); -- 
    final_index_ack_5211_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1333_offset_inst_ack_0, ack => cp_elements(301)); -- 
    base_resize_ack_5217_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1333_base_resize_ack_0, ack => cp_elements(302)); -- 
    cpelement_group_303 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(301) & cp_elements(302));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(303),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_5222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(303), ack => array_obj_ref_1333_root_address_inst_req_0); -- 
    plus_base_ra_5223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1333_root_address_inst_ack_0, ack => cp_elements(304)); -- 
    plus_base_cr_5224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(304), ack => array_obj_ref_1333_root_address_inst_req_1); -- 
    plus_base_ca_5225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1333_root_address_inst_ack_1, ack => cp_elements(305)); -- 
    cp_elements(306) <= array_obj_ref_1333_final_reg_ack_0;
    cp_elements(307) <= cp_elements(296);
    cpelement_group_308 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(306) & cp_elements(307) & cp_elements(312));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5258_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => ptr_deref_1336_gather_scatter_req_0); -- 
    cp_elements(309) <= cp_elements(306);
    base_resize_req_5243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(309), ack => ptr_deref_1336_base_resize_req_0); -- 
    base_resize_ack_5244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1336_base_resize_ack_0, ack => cp_elements(310)); -- 
    sum_rename_req_5248_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(310), ack => ptr_deref_1336_root_address_inst_req_0); -- 
    sum_rename_ack_5249_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1336_root_address_inst_ack_0, ack => cp_elements(311)); -- 
    root_rename_req_5253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(311), ack => ptr_deref_1336_addr_0_req_0); -- 
    root_rename_ack_5254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1336_addr_0_ack_0, ack => cp_elements(312)); -- 
    split_ack_5259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1336_gather_scatter_ack_0, ack => cp_elements(313)); -- 
    rr_5266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(313), ack => ptr_deref_1336_store_0_req_0); -- 
    cp_elements(314) <= ptr_deref_1336_store_0_ack_0;
    cp_elements(315) <= cp_elements(314);
    cr_5277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => ptr_deref_1336_store_0_req_1); -- 
    ca_5278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1336_store_0_ack_1, ack => cp_elements(316)); -- 
    cp_elements(317) <= cp_elements(296);
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(317) & cp_elements(322));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => array_obj_ref_1343_final_reg_req_0); -- 
    cp_elements(319) <= cp_elements(296);
    base_resize_req_5289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => array_obj_ref_1343_base_resize_req_0); -- 
    base_resize_ack_5290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1343_base_resize_ack_0, ack => cp_elements(320)); -- 
    plus_base_rr_5295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(320), ack => array_obj_ref_1343_root_address_inst_req_0); -- 
    plus_base_ra_5296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1343_root_address_inst_ack_0, ack => cp_elements(321)); -- 
    plus_base_cr_5297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => array_obj_ref_1343_root_address_inst_req_1); -- 
    plus_base_ca_5298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1343_root_address_inst_ack_1, ack => cp_elements(322)); -- 
    final_reg_ack_5303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1343_final_reg_ack_0, ack => cp_elements(323)); -- 
    cpelement_group_324 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(323) & cp_elements(325));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(324),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(324), ack => type_cast_1347_inst_req_0); -- 
    cp_elements(325) <= cp_elements(296);
    cp_elements(326) <= type_cast_1347_inst_ack_0;
    cp_elements(327) <= cp_elements(296);
    cpelement_group_328 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(314) & cp_elements(326) & cp_elements(327) & cp_elements(344));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => ptr_deref_1350_gather_scatter_req_0); -- 
    cp_elements(329) <= cp_elements(326);
    base_resize_req_5326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => ptr_deref_1350_base_resize_req_0); -- 
    base_resize_ack_5327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_base_resize_ack_0, ack => cp_elements(330)); -- 
    sum_rename_req_5331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => ptr_deref_1350_root_address_inst_req_0); -- 
    cp_elements(331) <= ptr_deref_1350_root_address_inst_ack_0;
    cp_elements(332) <= cp_elements(331);
    rr_5339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(332), ack => ptr_deref_1350_addr_0_req_0); -- 
    ra_5340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_0_ack_0, ack => cp_elements(333)); -- 
    cr_5341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => ptr_deref_1350_addr_0_req_1); -- 
    ca_5342_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_0_ack_1, ack => cp_elements(334)); -- 
    cp_elements(335) <= cp_elements(331);
    rr_5346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => ptr_deref_1350_addr_1_req_0); -- 
    ra_5347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_1_ack_0, ack => cp_elements(336)); -- 
    cr_5348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => ptr_deref_1350_addr_1_req_1); -- 
    ca_5349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_1_ack_1, ack => cp_elements(337)); -- 
    cp_elements(338) <= cp_elements(331);
    rr_5353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => ptr_deref_1350_addr_2_req_0); -- 
    ra_5354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_2_ack_0, ack => cp_elements(339)); -- 
    cr_5355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => ptr_deref_1350_addr_2_req_1); -- 
    ca_5356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_2_ack_1, ack => cp_elements(340)); -- 
    cp_elements(341) <= cp_elements(331);
    rr_5360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => ptr_deref_1350_addr_3_req_0); -- 
    ra_5361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_3_ack_0, ack => cp_elements(342)); -- 
    cr_5362_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(342), ack => ptr_deref_1350_addr_3_req_1); -- 
    ca_5363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_addr_3_ack_1, ack => cp_elements(343)); -- 
    cpelement_group_344 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(334) & cp_elements(337) & cp_elements(340) & cp_elements(343));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(344),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(345) <= ptr_deref_1350_gather_scatter_ack_0;
    cp_elements(346) <= cp_elements(345);
    rr_5375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(346), ack => ptr_deref_1350_store_0_req_0); -- 
    ra_5376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_0_ack_0, ack => cp_elements(347)); -- 
    cp_elements(348) <= cp_elements(345);
    rr_5380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => ptr_deref_1350_store_1_req_0); -- 
    ra_5381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_1_ack_0, ack => cp_elements(349)); -- 
    cp_elements(350) <= cp_elements(345);
    rr_5385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => ptr_deref_1350_store_2_req_0); -- 
    ra_5386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_2_ack_0, ack => cp_elements(351)); -- 
    cp_elements(352) <= cp_elements(345);
    rr_5390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(352), ack => ptr_deref_1350_store_3_req_0); -- 
    ra_5391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_3_ack_0, ack => cp_elements(353)); -- 
    cpelement_group_354 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(349) & cp_elements(351) & cp_elements(353));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(354),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(355) <= cp_elements(354);
    cp_elements(356) <= cp_elements(355);
    cr_5401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => ptr_deref_1350_store_0_req_1); -- 
    ca_5402_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_0_ack_1, ack => cp_elements(357)); -- 
    cp_elements(358) <= cp_elements(355);
    cr_5406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(358), ack => ptr_deref_1350_store_1_req_1); -- 
    ca_5407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_1_ack_1, ack => cp_elements(359)); -- 
    cp_elements(360) <= cp_elements(355);
    cr_5411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => ptr_deref_1350_store_2_req_1); -- 
    ca_5412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_2_ack_1, ack => cp_elements(361)); -- 
    cp_elements(362) <= cp_elements(355);
    cr_5416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(362), ack => ptr_deref_1350_store_3_req_1); -- 
    ca_5417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1350_store_3_ack_1, ack => cp_elements(363)); -- 
    cpelement_group_364 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(357) & cp_elements(359) & cp_elements(361) & cp_elements(363));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(365) <= cp_elements(296);
    cpelement_group_366 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(365) & cp_elements(370));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(366),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(366), ack => array_obj_ref_1357_final_reg_req_0); -- 
    cp_elements(367) <= cp_elements(296);
    base_resize_req_5428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(367), ack => array_obj_ref_1357_base_resize_req_0); -- 
    base_resize_ack_5429_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1357_base_resize_ack_0, ack => cp_elements(368)); -- 
    plus_base_rr_5434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(368), ack => array_obj_ref_1357_root_address_inst_req_0); -- 
    plus_base_ra_5435_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1357_root_address_inst_ack_0, ack => cp_elements(369)); -- 
    plus_base_cr_5436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(369), ack => array_obj_ref_1357_root_address_inst_req_1); -- 
    plus_base_ca_5437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1357_root_address_inst_ack_1, ack => cp_elements(370)); -- 
    final_reg_ack_5442_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1357_final_reg_ack_0, ack => cp_elements(371)); -- 
    cpelement_group_372 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(371) & cp_elements(373));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(372),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(372), ack => type_cast_1361_inst_req_0); -- 
    cp_elements(373) <= cp_elements(296);
    ack_5452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => cp_elements(374)); -- 
    cpelement_group_375 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(376) & cp_elements(377));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(375),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(375), ack => type_cast_1365_inst_req_0); -- 
    cp_elements(376) <= cp_elements(296);
    cp_elements(377) <= cp_elements(296);
    cp_elements(378) <= type_cast_1365_inst_ack_0;
    cp_elements(379) <= cp_elements(296);
    cpelement_group_380 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(354) & cp_elements(378) & cp_elements(379) & cp_elements(396));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(380),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => ptr_deref_1368_gather_scatter_req_0); -- 
    cp_elements(381) <= cp_elements(378);
    base_resize_req_5475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => ptr_deref_1368_base_resize_req_0); -- 
    base_resize_ack_5476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_base_resize_ack_0, ack => cp_elements(382)); -- 
    sum_rename_req_5480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(382), ack => ptr_deref_1368_root_address_inst_req_0); -- 
    cp_elements(383) <= ptr_deref_1368_root_address_inst_ack_0;
    cp_elements(384) <= cp_elements(383);
    rr_5488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => ptr_deref_1368_addr_0_req_0); -- 
    ra_5489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_0_ack_0, ack => cp_elements(385)); -- 
    cr_5490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(385), ack => ptr_deref_1368_addr_0_req_1); -- 
    ca_5491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_0_ack_1, ack => cp_elements(386)); -- 
    cp_elements(387) <= cp_elements(383);
    rr_5495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(387), ack => ptr_deref_1368_addr_1_req_0); -- 
    ra_5496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_1_ack_0, ack => cp_elements(388)); -- 
    cr_5497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(388), ack => ptr_deref_1368_addr_1_req_1); -- 
    ca_5498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_1_ack_1, ack => cp_elements(389)); -- 
    cp_elements(390) <= cp_elements(383);
    rr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(390), ack => ptr_deref_1368_addr_2_req_0); -- 
    ra_5503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_2_ack_0, ack => cp_elements(391)); -- 
    cr_5504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(391), ack => ptr_deref_1368_addr_2_req_1); -- 
    ca_5505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_2_ack_1, ack => cp_elements(392)); -- 
    cp_elements(393) <= cp_elements(383);
    rr_5509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(393), ack => ptr_deref_1368_addr_3_req_0); -- 
    ra_5510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_3_ack_0, ack => cp_elements(394)); -- 
    cr_5511_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(394), ack => ptr_deref_1368_addr_3_req_1); -- 
    ca_5512_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_addr_3_ack_1, ack => cp_elements(395)); -- 
    cpelement_group_396 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(386) & cp_elements(389) & cp_elements(392) & cp_elements(395));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(396),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(397) <= ptr_deref_1368_gather_scatter_ack_0;
    cp_elements(398) <= cp_elements(397);
    rr_5524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(398), ack => ptr_deref_1368_store_0_req_0); -- 
    ra_5525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_0_ack_0, ack => cp_elements(399)); -- 
    cp_elements(400) <= cp_elements(397);
    rr_5529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(400), ack => ptr_deref_1368_store_1_req_0); -- 
    ra_5530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_1_ack_0, ack => cp_elements(401)); -- 
    cp_elements(402) <= cp_elements(397);
    rr_5534_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => ptr_deref_1368_store_2_req_0); -- 
    ra_5535_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_2_ack_0, ack => cp_elements(403)); -- 
    cp_elements(404) <= cp_elements(397);
    rr_5539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(404), ack => ptr_deref_1368_store_3_req_0); -- 
    ra_5540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_3_ack_0, ack => cp_elements(405)); -- 
    cpelement_group_406 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(399) & cp_elements(401) & cp_elements(403) & cp_elements(405));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(406),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(407) <= cp_elements(406);
    cr_5550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(407), ack => ptr_deref_1368_store_0_req_1); -- 
    ca_5551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_0_ack_1, ack => cp_elements(408)); -- 
    cp_elements(409) <= cp_elements(406);
    cr_5555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(409), ack => ptr_deref_1368_store_1_req_1); -- 
    ca_5556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_1_ack_1, ack => cp_elements(410)); -- 
    cp_elements(411) <= cp_elements(406);
    cr_5560_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => ptr_deref_1368_store_2_req_1); -- 
    ca_5561_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_2_ack_1, ack => cp_elements(412)); -- 
    cp_elements(413) <= cp_elements(406);
    cr_5565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(413), ack => ptr_deref_1368_store_3_req_1); -- 
    ca_5566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1368_store_3_ack_1, ack => cp_elements(414)); -- 
    cpelement_group_415 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(408) & cp_elements(410) & cp_elements(412) & cp_elements(414));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(415),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_416 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(417) & cp_elements(418));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(416),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(416), ack => type_cast_1374_inst_req_0); -- 
    cp_elements(417) <= cp_elements(296);
    cp_elements(418) <= cp_elements(296);
    ack_5576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1374_inst_ack_0, ack => cp_elements(419)); -- 
    base_resize_req_5587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(419), ack => array_obj_ref_1383_base_resize_req_0); -- 
    cp_elements(420) <= cp_elements(296);
    cpelement_group_421 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(420) & cp_elements(424));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(421),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(421), ack => array_obj_ref_1383_final_reg_req_0); -- 
    base_resize_ack_5588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1383_base_resize_ack_0, ack => cp_elements(422)); -- 
    plus_base_rr_5593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(422), ack => array_obj_ref_1383_root_address_inst_req_0); -- 
    plus_base_ra_5594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1383_root_address_inst_ack_0, ack => cp_elements(423)); -- 
    plus_base_cr_5595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(423), ack => array_obj_ref_1383_root_address_inst_req_1); -- 
    plus_base_ca_5596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1383_root_address_inst_ack_1, ack => cp_elements(424)); -- 
    final_reg_ack_5601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1383_final_reg_ack_0, ack => cp_elements(425)); -- 
    cpelement_group_426 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(425) & cp_elements(427));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(426),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(426), ack => binary_1389_inst_req_0); -- 
    cp_elements(427) <= cp_elements(296);
    ra_5611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1389_inst_ack_0, ack => cp_elements(428)); -- 
    cr_5612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(428), ack => binary_1389_inst_req_1); -- 
    ca_5613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1389_inst_ack_1, ack => cp_elements(429)); -- 
    cpelement_group_430 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(316) & cp_elements(364) & cp_elements(374) & cp_elements(415) & cp_elements(429));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(430),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(431) <= cp_elements(10);
    cp_elements(432) <= false;
    cp_elements(433) <= cp_elements(432);
    cp_elements(434) <= cp_elements(10);
    branch_req_5621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(434), ack => if_stmt_1391_branch_req_0); -- 
    cp_elements(435) <= cp_elements(434);
    cp_elements(436) <= cp_elements(435);
    if_choice_transition_5626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1391_branch_ack_1, ack => cp_elements(437)); -- 
    cp_elements(438) <= cp_elements(435);
    else_choice_transition_5630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1391_branch_ack_0, ack => cp_elements(439)); -- 
    cp_elements(440) <= cp_elements(11);
    cp_elements(441) <= cp_elements(440);
    cpelement_group_442 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(441) & cp_elements(443) & cp_elements(447));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(442),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(442), ack => ptr_deref_1399_gather_scatter_req_0); -- 
    cp_elements(443) <= cp_elements(440);
    cp_elements(444) <= cp_elements(443);
    base_resize_req_5648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => ptr_deref_1399_base_resize_req_0); -- 
    base_resize_ack_5649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1399_base_resize_ack_0, ack => cp_elements(445)); -- 
    sum_rename_req_5653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(445), ack => ptr_deref_1399_root_address_inst_req_0); -- 
    sum_rename_ack_5654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1399_root_address_inst_ack_0, ack => cp_elements(446)); -- 
    root_rename_req_5658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(446), ack => ptr_deref_1399_addr_0_req_0); -- 
    root_rename_ack_5659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1399_addr_0_ack_0, ack => cp_elements(447)); -- 
    split_ack_5664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1399_gather_scatter_ack_0, ack => cp_elements(448)); -- 
    rr_5671_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(448), ack => ptr_deref_1399_store_0_req_0); -- 
    ra_5672_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1399_store_0_ack_0, ack => cp_elements(449)); -- 
    cr_5682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => ptr_deref_1399_store_0_req_1); -- 
    ca_5683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1399_store_0_ack_1, ack => cp_elements(450)); -- 
    cp_elements(451) <= cp_elements(1024);
    cpelement_group_452 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(453) & cp_elements(469));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(452),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(453) <= cp_elements(451);
    cp_elements(454) <= cp_elements(453);
    base_resize_req_5699_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(454), ack => ptr_deref_1407_base_resize_req_0); -- 
    base_resize_ack_5700_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_base_resize_ack_0, ack => cp_elements(455)); -- 
    sum_rename_req_5704_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(455), ack => ptr_deref_1407_root_address_inst_req_0); -- 
    cp_elements(456) <= ptr_deref_1407_root_address_inst_ack_0;
    cp_elements(457) <= cp_elements(456);
    rr_5712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(457), ack => ptr_deref_1407_addr_0_req_0); -- 
    ra_5713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_0_ack_0, ack => cp_elements(458)); -- 
    cr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => ptr_deref_1407_addr_0_req_1); -- 
    ca_5715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_0_ack_1, ack => cp_elements(459)); -- 
    cp_elements(460) <= cp_elements(456);
    rr_5719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(460), ack => ptr_deref_1407_addr_1_req_0); -- 
    ra_5720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_1_ack_0, ack => cp_elements(461)); -- 
    cr_5721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => ptr_deref_1407_addr_1_req_1); -- 
    ca_5722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_1_ack_1, ack => cp_elements(462)); -- 
    cp_elements(463) <= cp_elements(456);
    rr_5726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(463), ack => ptr_deref_1407_addr_2_req_0); -- 
    ra_5727_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_2_ack_0, ack => cp_elements(464)); -- 
    cr_5728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(464), ack => ptr_deref_1407_addr_2_req_1); -- 
    ca_5729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_2_ack_1, ack => cp_elements(465)); -- 
    cp_elements(466) <= cp_elements(456);
    rr_5733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(466), ack => ptr_deref_1407_addr_3_req_0); -- 
    ra_5734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_3_ack_0, ack => cp_elements(467)); -- 
    cr_5735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(467), ack => ptr_deref_1407_addr_3_req_1); -- 
    ca_5736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_addr_3_ack_1, ack => cp_elements(468)); -- 
    cpelement_group_469 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(459) & cp_elements(462) & cp_elements(465) & cp_elements(468));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(469),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(470) <= cp_elements(452);
    rr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(470), ack => ptr_deref_1407_load_0_req_0); -- 
    ra_5747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_0_ack_0, ack => cp_elements(471)); -- 
    cp_elements(472) <= cp_elements(452);
    rr_5751_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(472), ack => ptr_deref_1407_load_1_req_0); -- 
    ra_5752_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_1_ack_0, ack => cp_elements(473)); -- 
    cp_elements(474) <= cp_elements(452);
    rr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(474), ack => ptr_deref_1407_load_2_req_0); -- 
    ra_5757_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_2_ack_0, ack => cp_elements(475)); -- 
    cp_elements(476) <= cp_elements(452);
    rr_5761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(476), ack => ptr_deref_1407_load_3_req_0); -- 
    ra_5762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_3_ack_0, ack => cp_elements(477)); -- 
    cpelement_group_478 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(471) & cp_elements(473) & cp_elements(475) & cp_elements(477));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(478),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(479) <= cp_elements(478);
    cp_elements(480) <= cp_elements(479);
    cr_5772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(480), ack => ptr_deref_1407_load_0_req_1); -- 
    ca_5773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_0_ack_1, ack => cp_elements(481)); -- 
    cp_elements(482) <= cp_elements(479);
    cr_5777_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(482), ack => ptr_deref_1407_load_1_req_1); -- 
    ca_5778_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_1_ack_1, ack => cp_elements(483)); -- 
    cp_elements(484) <= cp_elements(479);
    cr_5782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(484), ack => ptr_deref_1407_load_2_req_1); -- 
    ca_5783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_2_ack_1, ack => cp_elements(485)); -- 
    cp_elements(486) <= cp_elements(479);
    cr_5787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(486), ack => ptr_deref_1407_load_3_req_1); -- 
    ca_5788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_load_3_ack_1, ack => cp_elements(487)); -- 
    cpelement_group_488 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(481) & cp_elements(483) & cp_elements(485) & cp_elements(487));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(488),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_5789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(488), ack => ptr_deref_1407_gather_scatter_req_0); -- 
    merge_ack_5790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1407_gather_scatter_ack_0, ack => cp_elements(489)); -- 
    cpelement_group_490 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(489) & cp_elements(491));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(490),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5799_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => binary_1413_inst_req_0); -- 
    cp_elements(491) <= cp_elements(451);
    ra_5800_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1413_inst_ack_0, ack => cp_elements(492)); -- 
    cr_5801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(492), ack => binary_1413_inst_req_1); -- 
    ca_5802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1413_inst_ack_1, ack => cp_elements(493)); -- 
    cpelement_group_494 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(478) & cp_elements(493) & cp_elements(495) & cp_elements(511));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(494),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(494), ack => ptr_deref_1416_gather_scatter_req_0); -- 
    cp_elements(495) <= cp_elements(451);
    cp_elements(496) <= cp_elements(495);
    base_resize_req_5816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => ptr_deref_1416_base_resize_req_0); -- 
    base_resize_ack_5817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_base_resize_ack_0, ack => cp_elements(497)); -- 
    sum_rename_req_5821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(497), ack => ptr_deref_1416_root_address_inst_req_0); -- 
    cp_elements(498) <= ptr_deref_1416_root_address_inst_ack_0;
    cp_elements(499) <= cp_elements(498);
    rr_5829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => ptr_deref_1416_addr_0_req_0); -- 
    ra_5830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_0_ack_0, ack => cp_elements(500)); -- 
    cr_5831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => ptr_deref_1416_addr_0_req_1); -- 
    ca_5832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_0_ack_1, ack => cp_elements(501)); -- 
    cp_elements(502) <= cp_elements(498);
    rr_5836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(502), ack => ptr_deref_1416_addr_1_req_0); -- 
    ra_5837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_1_ack_0, ack => cp_elements(503)); -- 
    cr_5838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => ptr_deref_1416_addr_1_req_1); -- 
    ca_5839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_1_ack_1, ack => cp_elements(504)); -- 
    cp_elements(505) <= cp_elements(498);
    rr_5843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(505), ack => ptr_deref_1416_addr_2_req_0); -- 
    ra_5844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_2_ack_0, ack => cp_elements(506)); -- 
    cr_5845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => ptr_deref_1416_addr_2_req_1); -- 
    ca_5846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_2_ack_1, ack => cp_elements(507)); -- 
    cp_elements(508) <= cp_elements(498);
    rr_5850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(508), ack => ptr_deref_1416_addr_3_req_0); -- 
    ra_5851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_3_ack_0, ack => cp_elements(509)); -- 
    cr_5852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => ptr_deref_1416_addr_3_req_1); -- 
    ca_5853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_addr_3_ack_1, ack => cp_elements(510)); -- 
    cpelement_group_511 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(501) & cp_elements(504) & cp_elements(507) & cp_elements(510));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(511),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(512) <= ptr_deref_1416_gather_scatter_ack_0;
    cp_elements(513) <= cp_elements(512);
    rr_5865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(513), ack => ptr_deref_1416_store_0_req_0); -- 
    ra_5866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_0_ack_0, ack => cp_elements(514)); -- 
    cp_elements(515) <= cp_elements(512);
    rr_5870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => ptr_deref_1416_store_1_req_0); -- 
    ra_5871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_1_ack_0, ack => cp_elements(516)); -- 
    cp_elements(517) <= cp_elements(512);
    rr_5875_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => ptr_deref_1416_store_2_req_0); -- 
    ra_5876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_2_ack_0, ack => cp_elements(518)); -- 
    cp_elements(519) <= cp_elements(512);
    rr_5880_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => ptr_deref_1416_store_3_req_0); -- 
    ra_5881_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_3_ack_0, ack => cp_elements(520)); -- 
    cpelement_group_521 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(514) & cp_elements(516) & cp_elements(518) & cp_elements(520));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(521),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(522) <= cp_elements(521);
    cp_elements(523) <= cp_elements(522);
    cr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(523), ack => ptr_deref_1416_store_0_req_1); -- 
    ca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_0_ack_1, ack => cp_elements(524)); -- 
    cp_elements(525) <= cp_elements(522);
    cr_5896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(525), ack => ptr_deref_1416_store_1_req_1); -- 
    ca_5897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_1_ack_1, ack => cp_elements(526)); -- 
    cp_elements(527) <= cp_elements(522);
    cr_5901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(527), ack => ptr_deref_1416_store_2_req_1); -- 
    ca_5902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_2_ack_1, ack => cp_elements(528)); -- 
    cp_elements(529) <= cp_elements(522);
    cr_5906_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(529), ack => ptr_deref_1416_store_3_req_1); -- 
    ca_5907_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1416_store_3_ack_1, ack => cp_elements(530)); -- 
    cpelement_group_531 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(524) & cp_elements(526) & cp_elements(528) & cp_elements(530));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(531),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_532 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(521) & cp_elements(533) & cp_elements(549));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(532),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(533) <= cp_elements(451);
    cp_elements(534) <= cp_elements(533);
    base_resize_req_5920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(534), ack => ptr_deref_1421_base_resize_req_0); -- 
    base_resize_ack_5921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_base_resize_ack_0, ack => cp_elements(535)); -- 
    sum_rename_req_5925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(535), ack => ptr_deref_1421_root_address_inst_req_0); -- 
    cp_elements(536) <= ptr_deref_1421_root_address_inst_ack_0;
    cp_elements(537) <= cp_elements(536);
    rr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(537), ack => ptr_deref_1421_addr_0_req_0); -- 
    ra_5934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_0_ack_0, ack => cp_elements(538)); -- 
    cr_5935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => ptr_deref_1421_addr_0_req_1); -- 
    ca_5936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_0_ack_1, ack => cp_elements(539)); -- 
    cp_elements(540) <= cp_elements(536);
    rr_5940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(540), ack => ptr_deref_1421_addr_1_req_0); -- 
    ra_5941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_1_ack_0, ack => cp_elements(541)); -- 
    cr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => ptr_deref_1421_addr_1_req_1); -- 
    ca_5943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_1_ack_1, ack => cp_elements(542)); -- 
    cp_elements(543) <= cp_elements(536);
    rr_5947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(543), ack => ptr_deref_1421_addr_2_req_0); -- 
    ra_5948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_2_ack_0, ack => cp_elements(544)); -- 
    cr_5949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(544), ack => ptr_deref_1421_addr_2_req_1); -- 
    ca_5950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_2_ack_1, ack => cp_elements(545)); -- 
    cp_elements(546) <= cp_elements(536);
    rr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(546), ack => ptr_deref_1421_addr_3_req_0); -- 
    ra_5955_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_3_ack_0, ack => cp_elements(547)); -- 
    cr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(547), ack => ptr_deref_1421_addr_3_req_1); -- 
    ca_5957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_addr_3_ack_1, ack => cp_elements(548)); -- 
    cpelement_group_549 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(539) & cp_elements(542) & cp_elements(545) & cp_elements(548));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(549),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(550) <= cp_elements(532);
    rr_5967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => ptr_deref_1421_load_0_req_0); -- 
    ra_5968_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_0_ack_0, ack => cp_elements(551)); -- 
    cp_elements(552) <= cp_elements(532);
    rr_5972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => ptr_deref_1421_load_1_req_0); -- 
    ra_5973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_1_ack_0, ack => cp_elements(553)); -- 
    cp_elements(554) <= cp_elements(532);
    rr_5977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(554), ack => ptr_deref_1421_load_2_req_0); -- 
    ra_5978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_2_ack_0, ack => cp_elements(555)); -- 
    cp_elements(556) <= cp_elements(532);
    rr_5982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(556), ack => ptr_deref_1421_load_3_req_0); -- 
    ra_5983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_3_ack_0, ack => cp_elements(557)); -- 
    cpelement_group_558 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(551) & cp_elements(553) & cp_elements(555) & cp_elements(557));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(558),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(559) <= cp_elements(558);
    cr_5993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(559), ack => ptr_deref_1421_load_0_req_1); -- 
    ca_5994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_0_ack_1, ack => cp_elements(560)); -- 
    cp_elements(561) <= cp_elements(558);
    cr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => ptr_deref_1421_load_1_req_1); -- 
    ca_5999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_1_ack_1, ack => cp_elements(562)); -- 
    cp_elements(563) <= cp_elements(558);
    cr_6003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(563), ack => ptr_deref_1421_load_2_req_1); -- 
    ca_6004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_2_ack_1, ack => cp_elements(564)); -- 
    cp_elements(565) <= cp_elements(558);
    cr_6008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(565), ack => ptr_deref_1421_load_3_req_1); -- 
    ca_6009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_load_3_ack_1, ack => cp_elements(566)); -- 
    cpelement_group_567 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(560) & cp_elements(562) & cp_elements(564) & cp_elements(566));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(567),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_6010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(567), ack => ptr_deref_1421_gather_scatter_req_0); -- 
    merge_ack_6011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1421_gather_scatter_ack_0, ack => cp_elements(568)); -- 
    cpelement_group_569 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(568) & cp_elements(570));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(569),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(569), ack => binary_1427_inst_req_0); -- 
    cp_elements(570) <= cp_elements(451);
    ra_6021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1427_inst_ack_0, ack => cp_elements(571)); -- 
    cr_6022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => binary_1427_inst_req_1); -- 
    ca_6023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1427_inst_ack_1, ack => cp_elements(572)); -- 
    cpelement_group_573 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(531) & cp_elements(572));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(573),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(574) <= cp_elements(12);
    cp_elements(575) <= false;
    cp_elements(576) <= cp_elements(575);
    cp_elements(577) <= cp_elements(12);
    branch_req_6031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(577), ack => if_stmt_1429_branch_req_0); -- 
    cp_elements(578) <= cp_elements(577);
    cp_elements(579) <= cp_elements(578);
    if_choice_transition_6036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1429_branch_ack_1, ack => cp_elements(580)); -- 
    cp_elements(581) <= cp_elements(578);
    else_choice_transition_6040_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1429_branch_ack_0, ack => cp_elements(582)); -- 
    cp_elements(583) <= cp_elements(13);
    cpelement_group_584 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(585) & cp_elements(601));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(584),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(585) <= cp_elements(583);
    cp_elements(586) <= cp_elements(585);
    base_resize_req_6058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => ptr_deref_1438_base_resize_req_0); -- 
    base_resize_ack_6059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_base_resize_ack_0, ack => cp_elements(587)); -- 
    sum_rename_req_6063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(587), ack => ptr_deref_1438_root_address_inst_req_0); -- 
    cp_elements(588) <= ptr_deref_1438_root_address_inst_ack_0;
    cp_elements(589) <= cp_elements(588);
    rr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(589), ack => ptr_deref_1438_addr_0_req_0); -- 
    ra_6072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_0_ack_0, ack => cp_elements(590)); -- 
    cr_6073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(590), ack => ptr_deref_1438_addr_0_req_1); -- 
    ca_6074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_0_ack_1, ack => cp_elements(591)); -- 
    cp_elements(592) <= cp_elements(588);
    rr_6078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(592), ack => ptr_deref_1438_addr_1_req_0); -- 
    ra_6079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_1_ack_0, ack => cp_elements(593)); -- 
    cr_6080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => ptr_deref_1438_addr_1_req_1); -- 
    ca_6081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_1_ack_1, ack => cp_elements(594)); -- 
    cp_elements(595) <= cp_elements(588);
    rr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => ptr_deref_1438_addr_2_req_0); -- 
    ra_6086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_2_ack_0, ack => cp_elements(596)); -- 
    cr_6087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(596), ack => ptr_deref_1438_addr_2_req_1); -- 
    ca_6088_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_2_ack_1, ack => cp_elements(597)); -- 
    cp_elements(598) <= cp_elements(588);
    rr_6092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(598), ack => ptr_deref_1438_addr_3_req_0); -- 
    ra_6093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_3_ack_0, ack => cp_elements(599)); -- 
    cr_6094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(599), ack => ptr_deref_1438_addr_3_req_1); -- 
    ca_6095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_addr_3_ack_1, ack => cp_elements(600)); -- 
    cpelement_group_601 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(591) & cp_elements(594) & cp_elements(597) & cp_elements(600));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(601),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(602) <= cp_elements(584);
    rr_6105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(602), ack => ptr_deref_1438_load_0_req_0); -- 
    ra_6106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_0_ack_0, ack => cp_elements(603)); -- 
    cp_elements(604) <= cp_elements(584);
    rr_6110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(604), ack => ptr_deref_1438_load_1_req_0); -- 
    ra_6111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_1_ack_0, ack => cp_elements(605)); -- 
    cp_elements(606) <= cp_elements(584);
    rr_6115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(606), ack => ptr_deref_1438_load_2_req_0); -- 
    ra_6116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_2_ack_0, ack => cp_elements(607)); -- 
    cp_elements(608) <= cp_elements(584);
    rr_6120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(608), ack => ptr_deref_1438_load_3_req_0); -- 
    ra_6121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_3_ack_0, ack => cp_elements(609)); -- 
    cpelement_group_610 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(603) & cp_elements(605) & cp_elements(607) & cp_elements(609));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(610),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(611) <= cp_elements(610);
    cr_6131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(611), ack => ptr_deref_1438_load_0_req_1); -- 
    ca_6132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_0_ack_1, ack => cp_elements(612)); -- 
    cp_elements(613) <= cp_elements(610);
    cr_6136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(613), ack => ptr_deref_1438_load_1_req_1); -- 
    ca_6137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_1_ack_1, ack => cp_elements(614)); -- 
    cp_elements(615) <= cp_elements(610);
    cr_6141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(615), ack => ptr_deref_1438_load_2_req_1); -- 
    ca_6142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_2_ack_1, ack => cp_elements(616)); -- 
    cp_elements(617) <= cp_elements(610);
    cr_6146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(617), ack => ptr_deref_1438_load_3_req_1); -- 
    ca_6147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_load_3_ack_1, ack => cp_elements(618)); -- 
    cpelement_group_619 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(612) & cp_elements(614) & cp_elements(616) & cp_elements(618));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(619),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_6148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(619), ack => ptr_deref_1438_gather_scatter_req_0); -- 
    merge_ack_6149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1438_gather_scatter_ack_0, ack => cp_elements(620)); -- 
    cpelement_group_621 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(622) & cp_elements(638));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(622) <= cp_elements(583);
    cp_elements(623) <= cp_elements(622);
    base_resize_req_6162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(623), ack => ptr_deref_1442_base_resize_req_0); -- 
    base_resize_ack_6163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_base_resize_ack_0, ack => cp_elements(624)); -- 
    sum_rename_req_6167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(624), ack => ptr_deref_1442_root_address_inst_req_0); -- 
    cp_elements(625) <= ptr_deref_1442_root_address_inst_ack_0;
    cp_elements(626) <= cp_elements(625);
    rr_6175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(626), ack => ptr_deref_1442_addr_0_req_0); -- 
    ra_6176_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_0_ack_0, ack => cp_elements(627)); -- 
    cr_6177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(627), ack => ptr_deref_1442_addr_0_req_1); -- 
    ca_6178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_0_ack_1, ack => cp_elements(628)); -- 
    cp_elements(629) <= cp_elements(625);
    rr_6182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(629), ack => ptr_deref_1442_addr_1_req_0); -- 
    ra_6183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_1_ack_0, ack => cp_elements(630)); -- 
    cr_6184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => ptr_deref_1442_addr_1_req_1); -- 
    ca_6185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_1_ack_1, ack => cp_elements(631)); -- 
    cp_elements(632) <= cp_elements(625);
    rr_6189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(632), ack => ptr_deref_1442_addr_2_req_0); -- 
    ra_6190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_2_ack_0, ack => cp_elements(633)); -- 
    cr_6191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(633), ack => ptr_deref_1442_addr_2_req_1); -- 
    ca_6192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_2_ack_1, ack => cp_elements(634)); -- 
    cp_elements(635) <= cp_elements(625);
    rr_6196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(635), ack => ptr_deref_1442_addr_3_req_0); -- 
    ra_6197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_3_ack_0, ack => cp_elements(636)); -- 
    cr_6198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => ptr_deref_1442_addr_3_req_1); -- 
    ca_6199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_addr_3_ack_1, ack => cp_elements(637)); -- 
    cpelement_group_638 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(628) & cp_elements(631) & cp_elements(634) & cp_elements(637));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(638),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(639) <= cp_elements(621);
    rr_6209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => ptr_deref_1442_load_0_req_0); -- 
    ra_6210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_0_ack_0, ack => cp_elements(640)); -- 
    cp_elements(641) <= cp_elements(621);
    rr_6214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(641), ack => ptr_deref_1442_load_1_req_0); -- 
    ra_6215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_1_ack_0, ack => cp_elements(642)); -- 
    cp_elements(643) <= cp_elements(621);
    rr_6219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => ptr_deref_1442_load_2_req_0); -- 
    ra_6220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_2_ack_0, ack => cp_elements(644)); -- 
    cp_elements(645) <= cp_elements(621);
    rr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(645), ack => ptr_deref_1442_load_3_req_0); -- 
    ra_6225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_3_ack_0, ack => cp_elements(646)); -- 
    cpelement_group_647 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(640) & cp_elements(642) & cp_elements(644) & cp_elements(646));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(647),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(648) <= cp_elements(647);
    cr_6235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(648), ack => ptr_deref_1442_load_0_req_1); -- 
    ca_6236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_0_ack_1, ack => cp_elements(649)); -- 
    cp_elements(650) <= cp_elements(647);
    cr_6240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(650), ack => ptr_deref_1442_load_1_req_1); -- 
    ca_6241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_1_ack_1, ack => cp_elements(651)); -- 
    cp_elements(652) <= cp_elements(647);
    cr_6245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => ptr_deref_1442_load_2_req_1); -- 
    ca_6246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_2_ack_1, ack => cp_elements(653)); -- 
    cp_elements(654) <= cp_elements(647);
    cr_6250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ptr_deref_1442_load_3_req_1); -- 
    ca_6251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_load_3_ack_1, ack => cp_elements(655)); -- 
    cpelement_group_656 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(649) & cp_elements(651) & cp_elements(653) & cp_elements(655));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(656),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_6252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(656), ack => ptr_deref_1442_gather_scatter_req_0); -- 
    merge_ack_6253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1442_gather_scatter_ack_0, ack => cp_elements(657)); -- 
    cpelement_group_658 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(620) & cp_elements(657) & cp_elements(659));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(658),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(658), ack => binary_1447_inst_req_0); -- 
    cp_elements(659) <= cp_elements(583);
    ra_6264_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1447_inst_ack_0, ack => cp_elements(660)); -- 
    cr_6265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(660), ack => binary_1447_inst_req_1); -- 
    ca_6266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1447_inst_ack_1, ack => cp_elements(661)); -- 
    cp_elements(662) <= cp_elements(661);
    cp_elements(663) <= false;
    cp_elements(664) <= cp_elements(663);
    cp_elements(665) <= cp_elements(661);
    branch_req_6274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(665), ack => if_stmt_1449_branch_req_0); -- 
    cp_elements(666) <= cp_elements(665);
    cp_elements(667) <= cp_elements(666);
    if_choice_transition_6279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1449_branch_ack_1, ack => cp_elements(668)); -- 
    cp_elements(669) <= cp_elements(666);
    else_choice_transition_6283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1449_branch_ack_0, ack => cp_elements(670)); -- 
    cpelement_group_671 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(687));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(671),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(672) <= cp_elements(14);
    base_resize_req_6301_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(672), ack => ptr_deref_1458_base_resize_req_0); -- 
    base_resize_ack_6302_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_base_resize_ack_0, ack => cp_elements(673)); -- 
    sum_rename_req_6306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(673), ack => ptr_deref_1458_root_address_inst_req_0); -- 
    cp_elements(674) <= ptr_deref_1458_root_address_inst_ack_0;
    cp_elements(675) <= cp_elements(674);
    rr_6314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(675), ack => ptr_deref_1458_addr_0_req_0); -- 
    ra_6315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_0_ack_0, ack => cp_elements(676)); -- 
    cr_6316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(676), ack => ptr_deref_1458_addr_0_req_1); -- 
    ca_6317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_0_ack_1, ack => cp_elements(677)); -- 
    cp_elements(678) <= cp_elements(674);
    rr_6321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => ptr_deref_1458_addr_1_req_0); -- 
    ra_6322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_1_ack_0, ack => cp_elements(679)); -- 
    cr_6323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(679), ack => ptr_deref_1458_addr_1_req_1); -- 
    ca_6324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_1_ack_1, ack => cp_elements(680)); -- 
    cp_elements(681) <= cp_elements(674);
    rr_6328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(681), ack => ptr_deref_1458_addr_2_req_0); -- 
    ra_6329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_2_ack_0, ack => cp_elements(682)); -- 
    cr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => ptr_deref_1458_addr_2_req_1); -- 
    ca_6331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_2_ack_1, ack => cp_elements(683)); -- 
    cp_elements(684) <= cp_elements(674);
    rr_6335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(684), ack => ptr_deref_1458_addr_3_req_0); -- 
    ra_6336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_3_ack_0, ack => cp_elements(685)); -- 
    cr_6337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(685), ack => ptr_deref_1458_addr_3_req_1); -- 
    ca_6338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_addr_3_ack_1, ack => cp_elements(686)); -- 
    cpelement_group_687 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(677) & cp_elements(680) & cp_elements(683) & cp_elements(686));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(687),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(688) <= cp_elements(671);
    rr_6348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(688), ack => ptr_deref_1458_load_0_req_0); -- 
    ra_6349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_0_ack_0, ack => cp_elements(689)); -- 
    cp_elements(690) <= cp_elements(671);
    rr_6353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => ptr_deref_1458_load_1_req_0); -- 
    ra_6354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_1_ack_0, ack => cp_elements(691)); -- 
    cp_elements(692) <= cp_elements(671);
    rr_6358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(692), ack => ptr_deref_1458_load_2_req_0); -- 
    ra_6359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_2_ack_0, ack => cp_elements(693)); -- 
    cp_elements(694) <= cp_elements(671);
    rr_6363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => ptr_deref_1458_load_3_req_0); -- 
    ra_6364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_3_ack_0, ack => cp_elements(695)); -- 
    cpelement_group_696 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(689) & cp_elements(691) & cp_elements(693) & cp_elements(695));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(696),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(697) <= cp_elements(696);
    cr_6374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(697), ack => ptr_deref_1458_load_0_req_1); -- 
    ca_6375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_0_ack_1, ack => cp_elements(698)); -- 
    cp_elements(699) <= cp_elements(696);
    cr_6379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => ptr_deref_1458_load_1_req_1); -- 
    ca_6380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_1_ack_1, ack => cp_elements(700)); -- 
    cp_elements(701) <= cp_elements(696);
    cr_6384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => ptr_deref_1458_load_2_req_1); -- 
    ca_6385_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_2_ack_1, ack => cp_elements(702)); -- 
    cp_elements(703) <= cp_elements(696);
    cr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(703), ack => ptr_deref_1458_load_3_req_1); -- 
    ca_6390_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_load_3_ack_1, ack => cp_elements(704)); -- 
    cpelement_group_705 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(698) & cp_elements(700) & cp_elements(702) & cp_elements(704));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(705),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_6391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => ptr_deref_1458_gather_scatter_req_0); -- 
    merge_ack_6392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1458_gather_scatter_ack_0, ack => cp_elements(706)); -- 
    cp_elements(707) <= cp_elements(1030);
    cp_elements(708) <= cp_elements(707);
    cpelement_group_709 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(708) & cp_elements(710) & cp_elements(714));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(709),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(709), ack => ptr_deref_1463_gather_scatter_req_0); -- 
    cp_elements(710) <= cp_elements(707);
    cp_elements(711) <= cp_elements(710);
    base_resize_req_6408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => ptr_deref_1463_base_resize_req_0); -- 
    base_resize_ack_6409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_base_resize_ack_0, ack => cp_elements(712)); -- 
    sum_rename_req_6413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(712), ack => ptr_deref_1463_root_address_inst_req_0); -- 
    sum_rename_ack_6414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_root_address_inst_ack_0, ack => cp_elements(713)); -- 
    root_rename_req_6418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(713), ack => ptr_deref_1463_addr_0_req_0); -- 
    root_rename_ack_6419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_addr_0_ack_0, ack => cp_elements(714)); -- 
    split_ack_6424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_gather_scatter_ack_0, ack => cp_elements(715)); -- 
    rr_6431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(715), ack => ptr_deref_1463_store_0_req_0); -- 
    ra_6432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_store_0_ack_0, ack => cp_elements(716)); -- 
    cr_6442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(716), ack => ptr_deref_1463_store_0_req_1); -- 
    ca_6443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_store_0_ack_1, ack => cp_elements(717)); -- 
    cra_6454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1470_call_ack_0, ack => cp_elements(718)); -- 
    ccr_6458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(718), ack => call_stmt_1470_call_req_1); -- 
    cca_6459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1470_call_ack_1, ack => cp_elements(719)); -- 
    cp_elements(720) <= cp_elements(180);
    cpelement_group_721 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(722) & cp_elements(730));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(721),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(721), ack => addr_of_1478_final_reg_req_0); -- 
    cp_elements(722) <= cp_elements(720);
    cp_elements(723) <= cp_elements(720);
    index_resize_req_6478_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(723), ack => array_obj_ref_1477_index_0_resize_req_0); -- 
    index_resize_ack_6479_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_index_0_resize_ack_0, ack => cp_elements(724)); -- 
    scale_rr_6483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(724), ack => array_obj_ref_1477_index_0_scale_req_0); -- 
    scale_ra_6484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_index_0_scale_ack_0, ack => cp_elements(725)); -- 
    scale_cr_6485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(725), ack => array_obj_ref_1477_index_0_scale_req_1); -- 
    scale_ca_6486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_index_0_scale_ack_1, ack => cp_elements(726)); -- 
    partial_sum_1_rr_6490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(726), ack => array_obj_ref_1477_index_sum_1_req_0); -- 
    partial_sum_1_ra_6491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_index_sum_1_ack_0, ack => cp_elements(727)); -- 
    partial_sum_1_cr_6492_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => array_obj_ref_1477_index_sum_1_req_1); -- 
    partial_sum_1_ca_6493_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_index_sum_1_ack_1, ack => cp_elements(728)); -- 
    final_index_req_6494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => array_obj_ref_1477_offset_inst_req_0); -- 
    final_index_ack_6495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_offset_inst_ack_0, ack => cp_elements(729)); -- 
    sum_rename_req_6499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => array_obj_ref_1477_root_address_inst_req_0); -- 
    sum_rename_ack_6500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1477_root_address_inst_ack_0, ack => cp_elements(730)); -- 
    cp_elements(731) <= addr_of_1478_final_reg_ack_0;
    cpelement_group_732 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(731) & cp_elements(736));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(732),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(732), ack => ptr_deref_1482_load_0_req_0); -- 
    cp_elements(733) <= cp_elements(731);
    base_resize_req_6518_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(733), ack => ptr_deref_1482_base_resize_req_0); -- 
    base_resize_ack_6519_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1482_base_resize_ack_0, ack => cp_elements(734)); -- 
    sum_rename_req_6523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(734), ack => ptr_deref_1482_root_address_inst_req_0); -- 
    sum_rename_ack_6524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1482_root_address_inst_ack_0, ack => cp_elements(735)); -- 
    root_rename_req_6528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => ptr_deref_1482_addr_0_req_0); -- 
    root_rename_ack_6529_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1482_addr_0_ack_0, ack => cp_elements(736)); -- 
    ra_6540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1482_load_0_ack_0, ack => cp_elements(737)); -- 
    cr_6550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(737), ack => ptr_deref_1482_load_0_req_1); -- 
    ca_6551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1482_load_0_ack_1, ack => cp_elements(738)); -- 
    merge_req_6552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(738), ack => ptr_deref_1482_gather_scatter_req_0); -- 
    merge_ack_6553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1482_gather_scatter_ack_0, ack => cp_elements(739)); -- 
    cpelement_group_740 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(739) & cp_elements(741));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(740),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => binary_1488_inst_req_0); -- 
    cp_elements(741) <= cp_elements(720);
    ra_6563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1488_inst_ack_0, ack => cp_elements(742)); -- 
    cr_6564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(742), ack => binary_1488_inst_req_1); -- 
    ca_6565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1488_inst_ack_1, ack => cp_elements(743)); -- 
    index_resize_req_6579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => array_obj_ref_1496_index_2_resize_req_0); -- 
    cpelement_group_744 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(745) & cp_elements(751));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(744),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => addr_of_1497_final_reg_req_0); -- 
    cp_elements(745) <= cp_elements(720);
    index_resize_ack_6580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1496_index_2_resize_ack_0, ack => cp_elements(746)); -- 
    scale_rename_req_6584_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(746), ack => array_obj_ref_1496_index_2_rename_req_0); -- 
    scale_rename_ack_6585_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1496_index_2_rename_ack_0, ack => cp_elements(747)); -- 
    partial_sum_1_rr_6589_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(747), ack => array_obj_ref_1496_index_sum_1_req_0); -- 
    partial_sum_1_ra_6590_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1496_index_sum_1_ack_0, ack => cp_elements(748)); -- 
    partial_sum_1_cr_6591_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(748), ack => array_obj_ref_1496_index_sum_1_req_1); -- 
    partial_sum_1_ca_6592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1496_index_sum_1_ack_1, ack => cp_elements(749)); -- 
    final_index_req_6593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => array_obj_ref_1496_offset_inst_req_0); -- 
    final_index_ack_6594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1496_offset_inst_ack_0, ack => cp_elements(750)); -- 
    sum_rename_req_6598_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(750), ack => array_obj_ref_1496_root_address_inst_req_0); -- 
    sum_rename_ack_6599_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1496_root_address_inst_ack_0, ack => cp_elements(751)); -- 
    cp_elements(752) <= addr_of_1497_final_reg_ack_0;
    cpelement_group_753 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(752) & cp_elements(757));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(753),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => ptr_deref_1501_load_0_req_0); -- 
    cp_elements(754) <= cp_elements(752);
    base_resize_req_6617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(754), ack => ptr_deref_1501_base_resize_req_0); -- 
    base_resize_ack_6618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1501_base_resize_ack_0, ack => cp_elements(755)); -- 
    sum_rename_req_6622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(755), ack => ptr_deref_1501_root_address_inst_req_0); -- 
    sum_rename_ack_6623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1501_root_address_inst_ack_0, ack => cp_elements(756)); -- 
    root_rename_req_6627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => ptr_deref_1501_addr_0_req_0); -- 
    root_rename_ack_6628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1501_addr_0_ack_0, ack => cp_elements(757)); -- 
    ra_6639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1501_load_0_ack_0, ack => cp_elements(758)); -- 
    cr_6649_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(758), ack => ptr_deref_1501_load_0_req_1); -- 
    ca_6650_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1501_load_0_ack_1, ack => cp_elements(759)); -- 
    merge_req_6651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(759), ack => ptr_deref_1501_gather_scatter_req_0); -- 
    merge_ack_6652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1501_gather_scatter_ack_0, ack => cp_elements(760)); -- 
    cpelement_group_761 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(760) & cp_elements(762));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(761),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(761), ack => binary_1507_inst_req_0); -- 
    cp_elements(762) <= cp_elements(720);
    ra_6662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1507_inst_ack_0, ack => cp_elements(763)); -- 
    cr_6663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(763), ack => binary_1507_inst_req_1); -- 
    ca_6664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1507_inst_ack_1, ack => cp_elements(764)); -- 
    cp_elements(765) <= cp_elements(764);
    cp_elements(766) <= false;
    cp_elements(767) <= cp_elements(766);
    cp_elements(768) <= cp_elements(764);
    branch_req_6672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(768), ack => if_stmt_1509_branch_req_0); -- 
    cp_elements(769) <= cp_elements(768);
    cp_elements(770) <= cp_elements(769);
    if_choice_transition_6677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1509_branch_ack_1, ack => cp_elements(771)); -- 
    cp_elements(772) <= cp_elements(769);
    else_choice_transition_6681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1509_branch_ack_0, ack => cp_elements(773)); -- 
    cp_elements(774) <= cp_elements(15);
    cpelement_group_775 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(776) & cp_elements(777));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(775),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(775), ack => binary_1520_inst_req_0); -- 
    cp_elements(776) <= cp_elements(774);
    cp_elements(777) <= cp_elements(774);
    ra_6696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1520_inst_ack_0, ack => cp_elements(778)); -- 
    cr_6697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(778), ack => binary_1520_inst_req_1); -- 
    ca_6698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1520_inst_ack_1, ack => cp_elements(779)); -- 
    index_resize_req_6712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(779), ack => array_obj_ref_1528_index_2_resize_req_0); -- 
    cpelement_group_780 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(781) & cp_elements(787));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(780),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6736_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(780), ack => addr_of_1529_final_reg_req_0); -- 
    cp_elements(781) <= cp_elements(774);
    index_resize_ack_6713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1528_index_2_resize_ack_0, ack => cp_elements(782)); -- 
    scale_rename_req_6717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(782), ack => array_obj_ref_1528_index_2_rename_req_0); -- 
    scale_rename_ack_6718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1528_index_2_rename_ack_0, ack => cp_elements(783)); -- 
    partial_sum_1_rr_6722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => array_obj_ref_1528_index_sum_1_req_0); -- 
    partial_sum_1_ra_6723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1528_index_sum_1_ack_0, ack => cp_elements(784)); -- 
    partial_sum_1_cr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => array_obj_ref_1528_index_sum_1_req_1); -- 
    partial_sum_1_ca_6725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1528_index_sum_1_ack_1, ack => cp_elements(785)); -- 
    final_index_req_6726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => array_obj_ref_1528_offset_inst_req_0); -- 
    final_index_ack_6727_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1528_offset_inst_ack_0, ack => cp_elements(786)); -- 
    sum_rename_req_6731_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(786), ack => array_obj_ref_1528_root_address_inst_req_0); -- 
    sum_rename_ack_6732_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1528_root_address_inst_ack_0, ack => cp_elements(787)); -- 
    cp_elements(788) <= addr_of_1529_final_reg_ack_0;
    cpelement_group_789 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(788) & cp_elements(793));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(789),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(789), ack => ptr_deref_1533_load_0_req_0); -- 
    cp_elements(790) <= cp_elements(788);
    base_resize_req_6750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => ptr_deref_1533_base_resize_req_0); -- 
    base_resize_ack_6751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_base_resize_ack_0, ack => cp_elements(791)); -- 
    sum_rename_req_6755_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => ptr_deref_1533_root_address_inst_req_0); -- 
    sum_rename_ack_6756_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_root_address_inst_ack_0, ack => cp_elements(792)); -- 
    root_rename_req_6760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(792), ack => ptr_deref_1533_addr_0_req_0); -- 
    root_rename_ack_6761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_addr_0_ack_0, ack => cp_elements(793)); -- 
    ra_6772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_load_0_ack_0, ack => cp_elements(794)); -- 
    cr_6782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => ptr_deref_1533_load_0_req_1); -- 
    ca_6783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_load_0_ack_1, ack => cp_elements(795)); -- 
    merge_req_6784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(795), ack => ptr_deref_1533_gather_scatter_req_0); -- 
    merge_ack_6785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_gather_scatter_ack_0, ack => cp_elements(796)); -- 
    cpelement_group_797 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(796) & cp_elements(798));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(797),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => binary_1539_inst_req_0); -- 
    cp_elements(798) <= cp_elements(774);
    ra_6795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1539_inst_ack_0, ack => cp_elements(799)); -- 
    cr_6796_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => binary_1539_inst_req_1); -- 
    ca_6797_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1539_inst_ack_1, ack => cp_elements(800)); -- 
    cp_elements(801) <= cp_elements(800);
    cp_elements(802) <= false;
    cp_elements(803) <= cp_elements(802);
    cp_elements(804) <= cp_elements(800);
    branch_req_6805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(804), ack => if_stmt_1541_branch_req_0); -- 
    cp_elements(805) <= cp_elements(804);
    cp_elements(806) <= cp_elements(805);
    if_choice_transition_6810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1541_branch_ack_1, ack => cp_elements(807)); -- 
    cp_elements(808) <= cp_elements(805);
    else_choice_transition_6814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1541_branch_ack_0, ack => cp_elements(809)); -- 
    cp_elements(810) <= cp_elements(16);
    cpelement_group_811 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(812) & cp_elements(813));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(811),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(811), ack => binary_1552_inst_req_0); -- 
    cp_elements(812) <= cp_elements(810);
    cp_elements(813) <= cp_elements(810);
    ra_6829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1552_inst_ack_0, ack => cp_elements(814)); -- 
    cr_6830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(814), ack => binary_1552_inst_req_1); -- 
    ca_6831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1552_inst_ack_1, ack => cp_elements(815)); -- 
    index_resize_req_6845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => array_obj_ref_1560_index_2_resize_req_0); -- 
    cpelement_group_816 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(817) & cp_elements(823));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(816),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(816), ack => addr_of_1561_final_reg_req_0); -- 
    cp_elements(817) <= cp_elements(810);
    index_resize_ack_6846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1560_index_2_resize_ack_0, ack => cp_elements(818)); -- 
    scale_rename_req_6850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(818), ack => array_obj_ref_1560_index_2_rename_req_0); -- 
    scale_rename_ack_6851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1560_index_2_rename_ack_0, ack => cp_elements(819)); -- 
    partial_sum_1_rr_6855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(819), ack => array_obj_ref_1560_index_sum_1_req_0); -- 
    partial_sum_1_ra_6856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1560_index_sum_1_ack_0, ack => cp_elements(820)); -- 
    partial_sum_1_cr_6857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(820), ack => array_obj_ref_1560_index_sum_1_req_1); -- 
    partial_sum_1_ca_6858_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1560_index_sum_1_ack_1, ack => cp_elements(821)); -- 
    final_index_req_6859_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(821), ack => array_obj_ref_1560_offset_inst_req_0); -- 
    final_index_ack_6860_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1560_offset_inst_ack_0, ack => cp_elements(822)); -- 
    sum_rename_req_6864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(822), ack => array_obj_ref_1560_root_address_inst_req_0); -- 
    sum_rename_ack_6865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1560_root_address_inst_ack_0, ack => cp_elements(823)); -- 
    cp_elements(824) <= addr_of_1561_final_reg_ack_0;
    cpelement_group_825 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(824) & cp_elements(829));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(825),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(825), ack => ptr_deref_1565_load_0_req_0); -- 
    cp_elements(826) <= cp_elements(824);
    base_resize_req_6883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(826), ack => ptr_deref_1565_base_resize_req_0); -- 
    base_resize_ack_6884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1565_base_resize_ack_0, ack => cp_elements(827)); -- 
    sum_rename_req_6888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(827), ack => ptr_deref_1565_root_address_inst_req_0); -- 
    sum_rename_ack_6889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1565_root_address_inst_ack_0, ack => cp_elements(828)); -- 
    root_rename_req_6893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => ptr_deref_1565_addr_0_req_0); -- 
    root_rename_ack_6894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1565_addr_0_ack_0, ack => cp_elements(829)); -- 
    ra_6905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1565_load_0_ack_0, ack => cp_elements(830)); -- 
    cr_6915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(830), ack => ptr_deref_1565_load_0_req_1); -- 
    ca_6916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1565_load_0_ack_1, ack => cp_elements(831)); -- 
    merge_req_6917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(831), ack => ptr_deref_1565_gather_scatter_req_0); -- 
    merge_ack_6918_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1565_gather_scatter_ack_0, ack => cp_elements(832)); -- 
    cpelement_group_833 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(834) & cp_elements(837));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(833),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(833), ack => binary_1574_inst_req_0); -- 
    cp_elements(834) <= cp_elements(810);
    cpelement_group_835 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(832) & cp_elements(836));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(835),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => type_cast_1570_inst_req_0); -- 
    cp_elements(836) <= cp_elements(810);
    ack_6930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_0, ack => cp_elements(837)); -- 
    ra_6935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1574_inst_ack_0, ack => cp_elements(838)); -- 
    cr_6936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(838), ack => binary_1574_inst_req_1); -- 
    ca_6937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1574_inst_ack_1, ack => cp_elements(839)); -- 
    cp_elements(840) <= cp_elements(839);
    cp_elements(841) <= false;
    cp_elements(842) <= cp_elements(841);
    cp_elements(843) <= cp_elements(839);
    branch_req_6945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(843), ack => if_stmt_1576_branch_req_0); -- 
    cp_elements(844) <= cp_elements(843);
    cp_elements(845) <= cp_elements(844);
    if_choice_transition_6950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1576_branch_ack_1, ack => cp_elements(846)); -- 
    cp_elements(847) <= cp_elements(844);
    else_choice_transition_6954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1576_branch_ack_0, ack => cp_elements(848)); -- 
    cp_elements(849) <= cp_elements(17);
    cpelement_group_850 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(851) & cp_elements(855));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(850),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(850), ack => binary_1589_inst_req_0); -- 
    cp_elements(851) <= cp_elements(849);
    cpelement_group_852 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(853) & cp_elements(854));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(852),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(852), ack => type_cast_1585_inst_req_0); -- 
    cp_elements(853) <= cp_elements(849);
    cp_elements(854) <= cp_elements(849);
    ack_6971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_0, ack => cp_elements(855)); -- 
    ra_6976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1589_inst_ack_0, ack => cp_elements(856)); -- 
    cr_6977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(856), ack => binary_1589_inst_req_1); -- 
    ca_6978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1589_inst_ack_1, ack => cp_elements(857)); -- 
    cp_elements(858) <= cp_elements(857);
    cp_elements(859) <= false;
    cp_elements(860) <= cp_elements(859);
    cp_elements(861) <= cp_elements(857);
    branch_req_6986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(861), ack => if_stmt_1591_branch_req_0); -- 
    cp_elements(862) <= cp_elements(861);
    cp_elements(863) <= cp_elements(862);
    if_choice_transition_6991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1591_branch_ack_1, ack => cp_elements(864)); -- 
    cp_elements(865) <= cp_elements(862);
    else_choice_transition_6995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1591_branch_ack_0, ack => cp_elements(866)); -- 
    cp_elements(867) <= cp_elements(18);
    cpelement_group_868 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(869) & cp_elements(870));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(868),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => binary_1602_inst_req_0); -- 
    cp_elements(869) <= cp_elements(867);
    cp_elements(870) <= cp_elements(867);
    ra_7010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1602_inst_ack_0, ack => cp_elements(871)); -- 
    cr_7011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(871), ack => binary_1602_inst_req_1); -- 
    ca_7012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1602_inst_ack_1, ack => cp_elements(872)); -- 
    cp_elements(873) <= cp_elements(872);
    cp_elements(874) <= false;
    cp_elements(875) <= cp_elements(874);
    cp_elements(876) <= cp_elements(872);
    branch_req_7020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(876), ack => if_stmt_1604_branch_req_0); -- 
    cp_elements(877) <= cp_elements(876);
    cp_elements(878) <= cp_elements(877);
    if_choice_transition_7025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1604_branch_ack_1, ack => cp_elements(879)); -- 
    cp_elements(880) <= cp_elements(877);
    else_choice_transition_7029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1604_branch_ack_0, ack => cp_elements(881)); -- 
    cp_elements(882) <= cp_elements(19);
    cpelement_group_883 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(884) & cp_elements(885));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(883),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(883), ack => binary_1615_inst_req_0); -- 
    cp_elements(884) <= cp_elements(882);
    cp_elements(885) <= cp_elements(882);
    ra_7044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1615_inst_ack_0, ack => cp_elements(886)); -- 
    cr_7045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(886), ack => binary_1615_inst_req_1); -- 
    ca_7046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1615_inst_ack_1, ack => cp_elements(887)); -- 
    cp_elements(888) <= cp_elements(887);
    cp_elements(889) <= false;
    cp_elements(890) <= cp_elements(889);
    cp_elements(891) <= cp_elements(887);
    branch_req_7054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(891), ack => if_stmt_1617_branch_req_0); -- 
    cp_elements(892) <= cp_elements(891);
    cp_elements(893) <= cp_elements(892);
    if_choice_transition_7059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1617_branch_ack_1, ack => cp_elements(894)); -- 
    cp_elements(895) <= cp_elements(892);
    else_choice_transition_7063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1617_branch_ack_0, ack => cp_elements(896)); -- 
    cp_elements(897) <= cp_elements(20);
    cpelement_group_898 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(899) & cp_elements(903));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(898),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(898), ack => binary_1630_inst_req_0); -- 
    cp_elements(899) <= cp_elements(897);
    cpelement_group_900 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(901) & cp_elements(902));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(900),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7079_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(900), ack => type_cast_1626_inst_req_0); -- 
    cp_elements(901) <= cp_elements(897);
    cp_elements(902) <= cp_elements(897);
    ack_7080_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_0, ack => cp_elements(903)); -- 
    ra_7085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1630_inst_ack_0, ack => cp_elements(904)); -- 
    cr_7086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(904), ack => binary_1630_inst_req_1); -- 
    ca_7087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1630_inst_ack_1, ack => cp_elements(905)); -- 
    cp_elements(906) <= cp_elements(905);
    cp_elements(907) <= false;
    cp_elements(908) <= cp_elements(907);
    cp_elements(909) <= cp_elements(905);
    branch_req_7095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(909), ack => if_stmt_1632_branch_req_0); -- 
    cp_elements(910) <= cp_elements(909);
    cp_elements(911) <= cp_elements(910);
    if_choice_transition_7100_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1632_branch_ack_1, ack => cp_elements(912)); -- 
    cp_elements(913) <= cp_elements(910);
    else_choice_transition_7104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1632_branch_ack_0, ack => cp_elements(914)); -- 
    cp_elements(915) <= cp_elements(21);
    cpelement_group_916 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(917) & cp_elements(918));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(916),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(916), ack => binary_1643_inst_req_0); -- 
    cp_elements(917) <= cp_elements(915);
    cp_elements(918) <= cp_elements(915);
    ra_7119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1643_inst_ack_0, ack => cp_elements(919)); -- 
    cr_7120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(919), ack => binary_1643_inst_req_1); -- 
    ca_7121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1643_inst_ack_1, ack => cp_elements(920)); -- 
    cp_elements(921) <= cp_elements(920);
    cp_elements(922) <= false;
    cp_elements(923) <= cp_elements(922);
    cp_elements(924) <= cp_elements(920);
    branch_req_7129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(924), ack => if_stmt_1645_branch_req_0); -- 
    cp_elements(925) <= cp_elements(924);
    cp_elements(926) <= cp_elements(925);
    if_choice_transition_7134_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1645_branch_ack_1, ack => cp_elements(927)); -- 
    cp_elements(928) <= cp_elements(925);
    else_choice_transition_7138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1645_branch_ack_0, ack => cp_elements(929)); -- 
    cp_elements(930) <= cp_elements(22);
    cpelement_group_931 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(932) & cp_elements(933));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(931),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(931), ack => binary_1656_inst_req_0); -- 
    cp_elements(932) <= cp_elements(930);
    cp_elements(933) <= cp_elements(930);
    ra_7153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1656_inst_ack_0, ack => cp_elements(934)); -- 
    cr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(934), ack => binary_1656_inst_req_1); -- 
    ca_7155_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1656_inst_ack_1, ack => cp_elements(935)); -- 
    cp_elements(936) <= cp_elements(935);
    cp_elements(937) <= false;
    cp_elements(938) <= cp_elements(937);
    cp_elements(939) <= cp_elements(935);
    branch_req_7163_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => if_stmt_1658_branch_req_0); -- 
    cp_elements(940) <= cp_elements(939);
    cp_elements(941) <= cp_elements(940);
    if_choice_transition_7168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1658_branch_ack_1, ack => cp_elements(942)); -- 
    cp_elements(943) <= cp_elements(940);
    else_choice_transition_7172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1658_branch_ack_0, ack => cp_elements(944)); -- 
    cp_elements(945) <= cp_elements(23);
    cpelement_group_946 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(947) & cp_elements(948));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(946),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(946), ack => type_cast_1667_inst_req_0); -- 
    cp_elements(947) <= cp_elements(945);
    cp_elements(948) <= cp_elements(945);
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_0, ack => cp_elements(949)); -- 
    pipe_wreq_7192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => simple_obj_ref_1665_inst_req_0); -- 
    pipe_wack_7193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1665_inst_ack_0, ack => cp_elements(950)); -- 
    cp_elements(951) <= cp_elements(927);
    cpelement_group_952 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(953) & cp_elements(954));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(952),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(952), ack => type_cast_1673_inst_req_0); -- 
    cp_elements(953) <= cp_elements(951);
    cp_elements(954) <= cp_elements(951);
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_0, ack => cp_elements(955)); -- 
    pipe_wreq_7211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(955), ack => simple_obj_ref_1671_inst_req_0); -- 
    pipe_wack_7212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1671_inst_ack_0, ack => cp_elements(956)); -- 
    cp_elements(957) <= cp_elements(894);
    cpelement_group_958 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(959) & cp_elements(960));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(958),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(958), ack => type_cast_1679_inst_req_0); -- 
    cp_elements(959) <= cp_elements(957);
    cp_elements(960) <= cp_elements(957);
    ack_7225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1679_inst_ack_0, ack => cp_elements(961)); -- 
    pipe_wreq_7230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(961), ack => simple_obj_ref_1677_inst_req_0); -- 
    pipe_wack_7231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1677_inst_ack_0, ack => cp_elements(962)); -- 
    cp_elements(963) <= cp_elements(879);
    cpelement_group_964 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(965) & cp_elements(966));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(964),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(964), ack => type_cast_1685_inst_req_0); -- 
    cp_elements(965) <= cp_elements(963);
    cp_elements(966) <= cp_elements(963);
    ack_7244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1685_inst_ack_0, ack => cp_elements(967)); -- 
    pipe_wreq_7249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(967), ack => simple_obj_ref_1683_inst_req_0); -- 
    pipe_wack_7250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1683_inst_ack_0, ack => cp_elements(968)); -- 
    cp_elements(969) <= cp_elements(1052);
    cpelement_group_970 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(971) & cp_elements(972));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(970),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(970), ack => type_cast_1691_inst_req_0); -- 
    cp_elements(971) <= cp_elements(969);
    cp_elements(972) <= cp_elements(969);
    ack_7263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1691_inst_ack_0, ack => cp_elements(973)); -- 
    pipe_wreq_7268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(973), ack => simple_obj_ref_1689_inst_req_0); -- 
    pipe_wack_7269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1689_inst_ack_0, ack => cp_elements(974)); -- 
    cp_elements(975) <= false;
    cp_elements(976) <= cp_elements(975);
    ack_7318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_0, ack => cp_elements(977)); -- 
    phi_stmt_1174_req_7319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(977), ack => phi_stmt_1174_req_0); -- 
    cp_elements(978) <= OrReduce(cp_elements(79) & cp_elements(977));
    cp_elements(979) <= cp_elements(978);
    phi_stmt_1174_ack_7324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1174_ack_0, ack => cp_elements(980)); -- 
    cp_elements(981) <= false;
    cp_elements(982) <= cp_elements(981);
    cp_elements(983) <= false;
    cp_elements(984) <= cp_elements(983);
    cp_elements(985) <= OrReduce(cp_elements(164) & cp_elements(182));
    cp_elements(986) <= cp_elements(985);
    cp_elements(987) <= false;
    cp_elements(988) <= cp_elements(987);
    cp_elements(989) <= cp_elements(5);
    cp_elements(990) <= cp_elements(989);
    phi_stmt_1248_req_7378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(990), ack => phi_stmt_1248_req_1); -- 
    cp_elements(991) <= cp_elements(989);
    phi_stmt_1241_req_7390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(991), ack => phi_stmt_1241_req_1); -- 
    cpelement_group_992 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(990) & cp_elements(991));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(992),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(993) <= cp_elements(280);
    cp_elements(994) <= cp_elements(993);
    req_7403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(994), ack => type_cast_1251_inst_req_0); -- 
    ack_7404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => cp_elements(995)); -- 
    phi_stmt_1248_req_7405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(995), ack => phi_stmt_1248_req_0); -- 
    cp_elements(996) <= cp_elements(993);
    req_7415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(996), ack => type_cast_1244_inst_req_0); -- 
    ack_7416_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1244_inst_ack_0, ack => cp_elements(997)); -- 
    phi_stmt_1241_req_7417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(997), ack => phi_stmt_1241_req_0); -- 
    cpelement_group_998 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(995) & cp_elements(997));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(998),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(999) <= OrReduce(cp_elements(992) & cp_elements(998));
    cp_elements(1000) <= cp_elements(999);
    phi_stmt_1241_ack_7422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1241_ack_0, ack => cp_elements(1001)); -- 
    phi_stmt_1248_ack_7423_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1248_ack_0, ack => cp_elements(1002)); -- 
    cpelement_group_1003 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(1001) & cp_elements(1002));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1003),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(1004) <= false;
    cp_elements(1005) <= cp_elements(1004);
    cp_elements(1006) <= cp_elements(249);
    cp_elements(1007) <= cp_elements(249);
    req_7453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1007), ack => type_cast_1294_inst_req_0); -- 
    ack_7454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_0, ack => cp_elements(1008)); -- 
    cpelement_group_1009 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(1006) & cp_elements(1008));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1009),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1289_req_7455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1009), ack => phi_stmt_1289_req_1); -- 
    cp_elements(1010) <= cp_elements(261);
    req_7468_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1010), ack => type_cast_1292_inst_req_0); -- 
    ack_7469_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1292_inst_ack_0, ack => cp_elements(1011)); -- 
    cp_elements(1012) <= cp_elements(261);
    cpelement_group_1013 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(1011) & cp_elements(1012));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1013),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1289_req_7475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1013), ack => phi_stmt_1289_req_0); -- 
    cp_elements(1014) <= OrReduce(cp_elements(1009) & cp_elements(1013));
    cp_elements(1015) <= cp_elements(1014);
    phi_stmt_1289_ack_7480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1289_ack_0, ack => cp_elements(1016)); -- 
    cp_elements(1017) <= false;
    cp_elements(1018) <= cp_elements(1017);
    cp_elements(1019) <= false;
    cp_elements(1020) <= cp_elements(1019);
    cp_elements(1021) <= false;
    cp_elements(1022) <= cp_elements(1021);
    cp_elements(1023) <= OrReduce(cp_elements(437) & cp_elements(450));
    cp_elements(1024) <= cp_elements(1023);
    cp_elements(1025) <= false;
    cp_elements(1026) <= cp_elements(1025);
    cp_elements(1027) <= false;
    cp_elements(1028) <= cp_elements(1027);
    cp_elements(1029) <= OrReduce(cp_elements(670) & cp_elements(706));
    cp_elements(1030) <= cp_elements(1029);
    cp_elements(1031) <= OrReduce(cp_elements(9) & cp_elements(216) & cp_elements(582) & cp_elements(717));
    cp_elements(1032) <= cp_elements(1031);
    crr_6453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1032), ack => call_stmt_1470_call_req_0); -- 
    cp_elements(1033) <= false;
    cp_elements(1034) <= cp_elements(1033);
    cp_elements(1035) <= false;
    cp_elements(1036) <= cp_elements(1035);
    cp_elements(1037) <= false;
    cp_elements(1038) <= cp_elements(1037);
    cp_elements(1039) <= false;
    cp_elements(1040) <= cp_elements(1039);
    cp_elements(1041) <= false;
    cp_elements(1042) <= cp_elements(1041);
    cp_elements(1043) <= false;
    cp_elements(1044) <= cp_elements(1043);
    cp_elements(1045) <= false;
    cp_elements(1046) <= cp_elements(1045);
    cp_elements(1047) <= false;
    cp_elements(1048) <= cp_elements(1047);
    cp_elements(1049) <= false;
    cp_elements(1050) <= cp_elements(1049);
    cp_elements(1051) <= OrReduce(cp_elements(773) & cp_elements(809) & cp_elements(881) & cp_elements(896) & cp_elements(929) & cp_elements(944));
    cp_elements(1052) <= cp_elements(1051);
    cp_elements(1053) <= OrReduce(cp_elements(719) & cp_elements(950) & cp_elements(956) & cp_elements(962) & cp_elements(968) & cp_elements(974));
    cp_elements(1054) <= cp_elements(1053);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal Pivot13_1590 : std_logic_vector(0 downto 0);
    signal Pivot15_1575 : std_logic_vector(0 downto 0);
    signal Pivot_1631 : std_logic_vector(0 downto 0);
    signal SwitchLeaf11_1603 : std_logic_vector(0 downto 0);
    signal SwitchLeaf7_1644 : std_logic_vector(0 downto 0);
    signal SwitchLeaf9_1616 : std_logic_vector(0 downto 0);
    signal SwitchLeaf_1657 : std_logic_vector(0 downto 0);
    signal array_obj_ref_1105_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1105_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1105_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1123_constant_part_of_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_index_partial_sum_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_offset_scale_factor_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_offset_scale_factor_2 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1123_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_constant_part_of_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_index_partial_sum_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_offset_scale_factor_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_offset_scale_factor_2 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1132_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1260_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_index_partial_sum_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_index_partial_sum_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1284_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1333_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1333_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1333_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1333_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1333_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1343_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1343_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1343_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1357_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1357_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1357_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1383_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1383_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1383_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1477_constant_part_of_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1477_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1477_index_partial_sum_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1477_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1477_offset_scale_factor_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1477_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1477_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1496_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_offset_scale_factor_2 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1496_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_offset_scale_factor_2 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1528_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_offset_scale_factor_2 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1560_root_address : std_logic_vector(8 downto 0);
    signal elt1x_xi5x_xix_xi_1134 : std_logic_vector(31 downto 0);
    signal eltx_xi3x_xix_xi_1125 : std_logic_vector(31 downto 0);
    signal exitcond_1307 : std_logic_vector(0 downto 0);
    signal ptr_deref_1113_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1113_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1113_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1113_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1113_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1113_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1137_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1137_resized_base_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1137_root_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1137_word_address_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1137_word_offset_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1141_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1141_resized_base_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1141_root_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1141_word_address_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1141_word_offset_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1265_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1265_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1336_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1336_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1336_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1336_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1336_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1336_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1350_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1350_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1350_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1350_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1350_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1350_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1368_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1368_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1368_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1368_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1368_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1368_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1399_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1399_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1399_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1399_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1399_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1399_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1407_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1407_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1407_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1407_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1407_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1416_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1416_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1416_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1416_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1416_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1416_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1421_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1421_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1421_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1421_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1421_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1438_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1438_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1438_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1438_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1438_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1442_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1442_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1442_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1442_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1442_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1458_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1458_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1458_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1458_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1458_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1463_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1463_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1463_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1463_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1463_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1463_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1482_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1482_resized_base_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1482_root_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1482_word_address_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1482_word_offset_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1501_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1501_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1501_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1501_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1501_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1533_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1565_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1565_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1565_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1565_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1565_word_offset_0 : std_logic_vector(8 downto 0);
    signal scevgep1x_xix_xix_xix_xix_xi_1286 : std_logic_vector(31 downto 0);
    signal scevgepx_xix_xix_xix_xix_xi_1262 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1093_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1118_resized : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1118_scaled : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1127_resized : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1127_scaled : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1213_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1213_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1221_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1221_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1257_resized : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1257_scaled : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1281_resized : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1281_scaled : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1474_resized : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1474_scaled : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1495_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1495_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1527_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1527_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1559_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1559_scaled : std_logic_vector(8 downto 0);
    signal tmp16_1099 : std_logic_vector(31 downto 0);
    signal tmp17_1106 : std_logic_vector(31 downto 0);
    signal tmp18_1110 : std_logic_vector(31 downto 0);
    signal tmp19_1114 : std_logic_vector(31 downto 0);
    signal tmp20_1147 : std_logic_vector(31 downto 0);
    signal tmp21_1152 : std_logic_vector(31 downto 0);
    signal tmp22_1158 : std_logic_vector(0 downto 0);
    signal tmp23_1171 : std_logic_vector(31 downto 0);
    signal tmp24_1174 : std_logic_vector(31 downto 0);
    signal tmp25_1189 : std_logic_vector(0 downto 0);
    signal tmp26_1204 : std_logic_vector(0 downto 0);
    signal tmp27_1214 : std_logic_vector(31 downto 0);
    signal tmp28_1220 : std_logic_vector(31 downto 0);
    signal tmp29_1231 : std_logic_vector(0 downto 0);
    signal tmp35_1241 : std_logic_vector(31 downto 0);
    signal tmp36_1248 : std_logic_vector(31 downto 0);
    signal tmp37_1266 : std_logic_vector(7 downto 0);
    signal tmp38_1272 : std_logic_vector(0 downto 0);
    signal tmp39_1289 : std_logic_vector(31 downto 0);
    signal tmp40_1301 : std_logic_vector(31 downto 0);
    signal tmp41_1320 : std_logic_vector(0 downto 0);
    signal tmp42_1334 : std_logic_vector(31 downto 0);
    signal tmp43_1344 : std_logic_vector(31 downto 0);
    signal tmp44_1348 : std_logic_vector(31 downto 0);
    signal tmp45_1358 : std_logic_vector(31 downto 0);
    signal tmp46_1362 : std_logic_vector(31 downto 0);
    signal tmp47_1366 : std_logic_vector(31 downto 0);
    signal tmp48_1375 : std_logic_vector(31 downto 0);
    signal tmp50_1384 : std_logic_vector(31 downto 0);
    signal tmp51_1390 : std_logic_vector(0 downto 0);
    signal tmp52_1408 : std_logic_vector(31 downto 0);
    signal tmp53_1414 : std_logic_vector(31 downto 0);
    signal tmp54_1422 : std_logic_vector(31 downto 0);
    signal tmp55_1428 : std_logic_vector(0 downto 0);
    signal tmp56_1439 : std_logic_vector(31 downto 0);
    signal tmp57_1443 : std_logic_vector(31 downto 0);
    signal tmp58_1448 : std_logic_vector(0 downto 0);
    signal tmp59_1459 : std_logic_vector(31 downto 0);
    signal tmp60_1479 : std_logic_vector(31 downto 0);
    signal tmp61_1483 : std_logic_vector(31 downto 0);
    signal tmp62_1489 : std_logic_vector(31 downto 0);
    signal tmp63_1498 : std_logic_vector(31 downto 0);
    signal tmp64_1502 : std_logic_vector(7 downto 0);
    signal tmp65_1508 : std_logic_vector(0 downto 0);
    signal tmp66_1530 : std_logic_vector(31 downto 0);
    signal tmp67_1534 : std_logic_vector(7 downto 0);
    signal tmp68_1540 : std_logic_vector(0 downto 0);
    signal tmp69_1562 : std_logic_vector(31 downto 0);
    signal tmp70_1566 : std_logic_vector(7 downto 0);
    signal tmp_1095 : std_logic_vector(31 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1177_wire : std_logic_vector(31 downto 0);
    signal type_cast_1180_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1184_wire : std_logic_vector(31 downto 0);
    signal type_cast_1187_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1199_wire : std_logic_vector(31 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1218_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1226_wire : std_logic_vector(31 downto 0);
    signal type_cast_1229_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1244_wire : std_logic_vector(31 downto 0);
    signal type_cast_1247_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1251_wire : std_logic_vector(31 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1270_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1292_wire : std_logic_vector(31 downto 0);
    signal type_cast_1294_wire : std_logic_vector(31 downto 0);
    signal type_cast_1299_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1318_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1352_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1370_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1426_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1465_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1487_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1538_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1551_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1570_wire : std_logic_vector(7 downto 0);
    signal type_cast_1573_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1585_wire : std_logic_vector(7 downto 0);
    signal type_cast_1588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1601_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1614_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1626_wire : std_logic_vector(7 downto 0);
    signal type_cast_1629_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1642_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1655_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1667_wire : std_logic_vector(31 downto 0);
    signal type_cast_1673_wire : std_logic_vector(31 downto 0);
    signal type_cast_1679_wire : std_logic_vector(31 downto 0);
    signal type_cast_1685_wire : std_logic_vector(31 downto 0);
    signal type_cast_1691_wire : std_logic_vector(31 downto 0);
    signal val2x_xi6x_xix_xi_1142 : std_logic_vector(31 downto 0);
    signal valx_xi4x_xix_xi_1138 : std_logic_vector(31 downto 0);
    signal xx_xsum26x_xi_1521 : std_logic_vector(31 downto 0);
    signal xx_xsum27x_xi_1553 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1105_final_offset <= "0000000000011100";
    array_obj_ref_1123_constant_part_of_offset <= "00000";
    array_obj_ref_1123_offset_scale_factor_0 <= "00101";
    array_obj_ref_1123_offset_scale_factor_1 <= "00001";
    array_obj_ref_1123_offset_scale_factor_2 <= "00001";
    array_obj_ref_1123_resized_base_address <= "00000";
    array_obj_ref_1132_constant_part_of_offset <= "00001";
    array_obj_ref_1132_offset_scale_factor_0 <= "00101";
    array_obj_ref_1132_offset_scale_factor_1 <= "00001";
    array_obj_ref_1132_offset_scale_factor_2 <= "00001";
    array_obj_ref_1132_resized_base_address <= "00000";
    array_obj_ref_1260_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1260_offset_scale_factor_0 <= "00000010000000";
    array_obj_ref_1260_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1260_resized_base_address <= "00000000000000";
    array_obj_ref_1284_constant_part_of_offset <= "00000000000001";
    array_obj_ref_1284_offset_scale_factor_0 <= "00000010000000";
    array_obj_ref_1284_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1284_resized_base_address <= "00000000000000";
    array_obj_ref_1333_constant_part_of_offset <= "11111111111111";
    array_obj_ref_1333_offset_scale_factor_0 <= "00000000000001";
    array_obj_ref_1343_final_offset <= "00000000000100";
    array_obj_ref_1357_final_offset <= "00000000001000";
    array_obj_ref_1383_final_offset <= "00000000001100";
    array_obj_ref_1477_constant_part_of_offset <= "00011";
    array_obj_ref_1477_offset_scale_factor_0 <= "00101";
    array_obj_ref_1477_offset_scale_factor_1 <= "00001";
    array_obj_ref_1477_resized_base_address <= "00000";
    array_obj_ref_1496_constant_part_of_offset <= "000000000";
    array_obj_ref_1496_offset_scale_factor_0 <= "001001000";
    array_obj_ref_1496_offset_scale_factor_1 <= "001000000";
    array_obj_ref_1496_offset_scale_factor_2 <= "000000001";
    array_obj_ref_1496_resized_base_address <= "000000000";
    array_obj_ref_1528_constant_part_of_offset <= "000000000";
    array_obj_ref_1528_offset_scale_factor_0 <= "001001000";
    array_obj_ref_1528_offset_scale_factor_1 <= "001000000";
    array_obj_ref_1528_offset_scale_factor_2 <= "000000001";
    array_obj_ref_1528_resized_base_address <= "000000000";
    array_obj_ref_1560_constant_part_of_offset <= "000000000";
    array_obj_ref_1560_offset_scale_factor_0 <= "001001000";
    array_obj_ref_1560_offset_scale_factor_1 <= "001000000";
    array_obj_ref_1560_offset_scale_factor_2 <= "000000001";
    array_obj_ref_1560_resized_base_address <= "000000000";
    ptr_deref_1113_word_offset_0 <= "0000000000000000";
    ptr_deref_1113_word_offset_1 <= "0000000000000001";
    ptr_deref_1113_word_offset_2 <= "0000000000000010";
    ptr_deref_1113_word_offset_3 <= "0000000000000011";
    ptr_deref_1137_word_offset_0 <= "00000";
    ptr_deref_1141_word_offset_0 <= "00000";
    ptr_deref_1265_word_offset_0 <= "00000000000000";
    ptr_deref_1336_word_offset_0 <= "00000000000000";
    ptr_deref_1350_word_offset_0 <= "00000000000000";
    ptr_deref_1350_word_offset_1 <= "00000000000001";
    ptr_deref_1350_word_offset_2 <= "00000000000010";
    ptr_deref_1350_word_offset_3 <= "00000000000011";
    ptr_deref_1368_word_offset_0 <= "00000000000000";
    ptr_deref_1368_word_offset_1 <= "00000000000001";
    ptr_deref_1368_word_offset_2 <= "00000000000010";
    ptr_deref_1368_word_offset_3 <= "00000000000011";
    ptr_deref_1399_word_offset_0 <= "00000000000000";
    ptr_deref_1407_word_offset_0 <= "00000000000000";
    ptr_deref_1407_word_offset_1 <= "00000000000001";
    ptr_deref_1407_word_offset_2 <= "00000000000010";
    ptr_deref_1407_word_offset_3 <= "00000000000011";
    ptr_deref_1416_word_offset_0 <= "00000000000000";
    ptr_deref_1416_word_offset_1 <= "00000000000001";
    ptr_deref_1416_word_offset_2 <= "00000000000010";
    ptr_deref_1416_word_offset_3 <= "00000000000011";
    ptr_deref_1421_word_offset_0 <= "00000000000000";
    ptr_deref_1421_word_offset_1 <= "00000000000001";
    ptr_deref_1421_word_offset_2 <= "00000000000010";
    ptr_deref_1421_word_offset_3 <= "00000000000011";
    ptr_deref_1438_word_offset_0 <= "00000000000000";
    ptr_deref_1438_word_offset_1 <= "00000000000001";
    ptr_deref_1438_word_offset_2 <= "00000000000010";
    ptr_deref_1438_word_offset_3 <= "00000000000011";
    ptr_deref_1442_word_offset_0 <= "00000000000000";
    ptr_deref_1442_word_offset_1 <= "00000000000001";
    ptr_deref_1442_word_offset_2 <= "00000000000010";
    ptr_deref_1442_word_offset_3 <= "00000000000011";
    ptr_deref_1458_word_offset_0 <= "00000000000000";
    ptr_deref_1458_word_offset_1 <= "00000000000001";
    ptr_deref_1458_word_offset_2 <= "00000000000010";
    ptr_deref_1458_word_offset_3 <= "00000000000011";
    ptr_deref_1463_word_offset_0 <= "00000000000000";
    ptr_deref_1482_word_offset_0 <= "00000";
    ptr_deref_1501_word_offset_0 <= "000000000";
    ptr_deref_1533_word_offset_0 <= "000000000";
    ptr_deref_1565_word_offset_0 <= "000000000";
    simple_obj_ref_1213_word_address_0 <= "0";
    simple_obj_ref_1221_word_address_0 <= "0";
    type_cast_1156_wire_constant <= "00000000000000000000000000000000";
    type_cast_1169_wire_constant <= "00000000000000000000000000000001";
    type_cast_1180_wire_constant <= "00000000000000000000000000000000";
    type_cast_1187_wire_constant <= "00000000000000000000000000000100";
    type_cast_1202_wire_constant <= "11111111111111111111111111111111";
    type_cast_1218_wire_constant <= "00000000000000000000000000000001";
    type_cast_1229_wire_constant <= "00000000000000000000000000000110";
    type_cast_1247_wire_constant <= "00000000000000000000000000000000";
    type_cast_1254_wire_constant <= "11111111111111111111111111111111";
    type_cast_1270_wire_constant <= "00000001";
    type_cast_1299_wire_constant <= "00000000000000000000000000000001";
    type_cast_1305_wire_constant <= "00000000000000000000000001000000";
    type_cast_1318_wire_constant <= "11111111111111111111111111111111";
    type_cast_1338_wire_constant <= "00010001";
    type_cast_1352_wire_constant <= "00000000000000000000011111110100";
    type_cast_1370_wire_constant <= "00000000000000000000000000000001";
    type_cast_1388_wire_constant <= "11111111111111111111111111111111";
    type_cast_1401_wire_constant <= "00000000";
    type_cast_1412_wire_constant <= "11111111111111111111111111111111";
    type_cast_1426_wire_constant <= "00000000000000000000000000000000";
    type_cast_1465_wire_constant <= "00000001";
    type_cast_1487_wire_constant <= "00000000000000000000000001001000";
    type_cast_1506_wire_constant <= "01110100";
    type_cast_1519_wire_constant <= "00000000000000000000000000000001";
    type_cast_1538_wire_constant <= "01101111";
    type_cast_1551_wire_constant <= "00000000000000000000000000000010";
    type_cast_1573_wire_constant <= "00110010";
    type_cast_1588_wire_constant <= "00110011";
    type_cast_1601_wire_constant <= "00110011";
    type_cast_1614_wire_constant <= "00110010";
    type_cast_1629_wire_constant <= "00110001";
    type_cast_1642_wire_constant <= "00110001";
    type_cast_1655_wire_constant <= "00110000";
    phi_stmt_1174: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1177_wire & type_cast_1180_wire_constant;
      req <= phi_stmt_1174_req_0 & phi_stmt_1174_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1174_ack_0,
          idata => idata,
          odata => tmp24_1174,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1174
    phi_stmt_1241: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1244_wire & type_cast_1247_wire_constant;
      req <= phi_stmt_1241_req_0 & phi_stmt_1241_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1241_ack_0,
          idata => idata,
          odata => tmp35_1241,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1241
    phi_stmt_1248: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1251_wire & type_cast_1254_wire_constant;
      req <= phi_stmt_1248_req_0 & phi_stmt_1248_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1248_ack_0,
          idata => idata,
          odata => tmp36_1248,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1248
    phi_stmt_1289: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1292_wire & type_cast_1294_wire;
      req <= phi_stmt_1289_req_0 & phi_stmt_1289_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1289_ack_0,
          idata => idata,
          odata => tmp39_1289,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1289
    addr_of_1124_final_reg: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1123_root_address, dout => eltx_xi3x_xix_xi_1125, req => addr_of_1124_final_reg_req_0, ack => addr_of_1124_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1133_final_reg: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1132_root_address, dout => elt1x_xi5x_xix_xi_1134, req => addr_of_1133_final_reg_req_0, ack => addr_of_1133_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1261_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1260_root_address, dout => scevgepx_xix_xix_xix_xix_xi_1262, req => addr_of_1261_final_reg_req_0, ack => addr_of_1261_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1285_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1284_root_address, dout => scevgep1x_xix_xix_xix_xix_xi_1286, req => addr_of_1285_final_reg_req_0, ack => addr_of_1285_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1478_final_reg: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1477_root_address, dout => tmp60_1479, req => addr_of_1478_final_reg_req_0, ack => addr_of_1478_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1497_final_reg: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1496_root_address, dout => tmp63_1498, req => addr_of_1497_final_reg_req_0, ack => addr_of_1497_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1529_final_reg: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1528_root_address, dout => tmp66_1530, req => addr_of_1529_final_reg_req_0, ack => addr_of_1529_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1561_final_reg: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1560_root_address, dout => tmp69_1562, req => addr_of_1561_final_reg_req_0, ack => addr_of_1561_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1105_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1099, dout => array_obj_ref_1105_resized_base_address, req => array_obj_ref_1105_base_resize_req_0, ack => array_obj_ref_1105_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1105_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1105_root_address, dout => tmp17_1106, req => array_obj_ref_1105_final_reg_req_0, ack => array_obj_ref_1105_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1123_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp24_1174, dout => simple_obj_ref_1118_resized, req => array_obj_ref_1123_index_0_resize_req_0, ack => array_obj_ref_1123_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1123_offset_inst: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 5, flow_through => true ) 
      port map( din => array_obj_ref_1123_index_partial_sum_1, dout => array_obj_ref_1123_final_offset, req => array_obj_ref_1123_offset_inst_req_0, ack => array_obj_ref_1123_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1132_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp24_1174, dout => simple_obj_ref_1127_resized, req => array_obj_ref_1132_index_0_resize_req_0, ack => array_obj_ref_1132_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1132_offset_inst: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 5, flow_through => true ) 
      port map( din => array_obj_ref_1132_index_partial_sum_1, dout => array_obj_ref_1132_final_offset, req => array_obj_ref_1132_offset_inst_req_0, ack => array_obj_ref_1132_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1260_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp35_1241, dout => simple_obj_ref_1257_resized, req => array_obj_ref_1260_index_0_resize_req_0, ack => array_obj_ref_1260_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1260_offset_inst: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 14, flow_through => true ) 
      port map( din => array_obj_ref_1260_index_partial_sum_1, dout => array_obj_ref_1260_final_offset, req => array_obj_ref_1260_offset_inst_req_0, ack => array_obj_ref_1260_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1284_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp35_1241, dout => simple_obj_ref_1281_resized, req => array_obj_ref_1284_index_0_resize_req_0, ack => array_obj_ref_1284_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1284_offset_inst: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 14, flow_through => true ) 
      port map( din => array_obj_ref_1284_index_partial_sum_1, dout => array_obj_ref_1284_final_offset, req => array_obj_ref_1284_offset_inst_req_0, ack => array_obj_ref_1284_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1333_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp39_1289, dout => array_obj_ref_1333_resized_base_address, req => array_obj_ref_1333_base_resize_req_0, ack => array_obj_ref_1333_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1333_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1333_root_address, dout => tmp42_1334, req => array_obj_ref_1333_final_reg_req_0, ack => array_obj_ref_1333_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1333_offset_inst: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 14, flow_through => true ) 
      port map( din => array_obj_ref_1333_constant_part_of_offset, dout => array_obj_ref_1333_final_offset, req => array_obj_ref_1333_offset_inst_req_0, ack => array_obj_ref_1333_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1343_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp39_1289, dout => array_obj_ref_1343_resized_base_address, req => array_obj_ref_1343_base_resize_req_0, ack => array_obj_ref_1343_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1343_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1343_root_address, dout => tmp43_1344, req => array_obj_ref_1343_final_reg_req_0, ack => array_obj_ref_1343_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1357_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp39_1289, dout => array_obj_ref_1357_resized_base_address, req => array_obj_ref_1357_base_resize_req_0, ack => array_obj_ref_1357_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1357_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1357_root_address, dout => tmp45_1358, req => array_obj_ref_1357_final_reg_req_0, ack => array_obj_ref_1357_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1383_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp48_1375, dout => array_obj_ref_1383_resized_base_address, req => array_obj_ref_1383_base_resize_req_0, ack => array_obj_ref_1383_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1383_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1383_root_address, dout => tmp50_1384, req => array_obj_ref_1383_final_reg_req_0, ack => array_obj_ref_1383_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1477_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp24_1174, dout => simple_obj_ref_1474_resized, req => array_obj_ref_1477_index_0_resize_req_0, ack => array_obj_ref_1477_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1477_offset_inst: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 5, flow_through => true ) 
      port map( din => array_obj_ref_1477_index_partial_sum_1, dout => array_obj_ref_1477_final_offset, req => array_obj_ref_1477_offset_inst_req_0, ack => array_obj_ref_1477_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1496_index_2_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp62_1489, dout => simple_obj_ref_1495_resized, req => array_obj_ref_1496_index_2_resize_req_0, ack => array_obj_ref_1496_index_2_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1496_offset_inst: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 9, flow_through => true ) 
      port map( din => array_obj_ref_1496_index_partial_sum_1, dout => array_obj_ref_1496_final_offset, req => array_obj_ref_1496_offset_inst_req_0, ack => array_obj_ref_1496_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1528_index_2_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => xx_xsum26x_xi_1521, dout => simple_obj_ref_1527_resized, req => array_obj_ref_1528_index_2_resize_req_0, ack => array_obj_ref_1528_index_2_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1528_offset_inst: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 9, flow_through => true ) 
      port map( din => array_obj_ref_1528_index_partial_sum_1, dout => array_obj_ref_1528_final_offset, req => array_obj_ref_1528_offset_inst_req_0, ack => array_obj_ref_1528_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1560_index_2_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => xx_xsum27x_xi_1553, dout => simple_obj_ref_1559_resized, req => array_obj_ref_1560_index_2_resize_req_0, ack => array_obj_ref_1560_index_2_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1560_offset_inst: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 9, flow_through => true ) 
      port map( din => array_obj_ref_1560_index_partial_sum_1, dout => array_obj_ref_1560_final_offset, req => array_obj_ref_1560_offset_inst_req_0, ack => array_obj_ref_1560_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1113_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_1110, dout => ptr_deref_1113_resized_base_address, req => ptr_deref_1113_base_resize_req_0, ack => ptr_deref_1113_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1137_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => eltx_xi3x_xix_xi_1125, dout => ptr_deref_1137_resized_base_address, req => ptr_deref_1137_base_resize_req_0, ack => ptr_deref_1137_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1141_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => elt1x_xi5x_xix_xi_1134, dout => ptr_deref_1141_resized_base_address, req => ptr_deref_1141_base_resize_req_0, ack => ptr_deref_1141_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1265_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => scevgepx_xix_xix_xix_xix_xi_1262, dout => ptr_deref_1265_resized_base_address, req => ptr_deref_1265_base_resize_req_0, ack => ptr_deref_1265_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1336_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp42_1334, dout => ptr_deref_1336_resized_base_address, req => ptr_deref_1336_base_resize_req_0, ack => ptr_deref_1336_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1350_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp44_1348, dout => ptr_deref_1350_resized_base_address, req => ptr_deref_1350_base_resize_req_0, ack => ptr_deref_1350_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1368_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1366, dout => ptr_deref_1368_resized_base_address, req => ptr_deref_1368_base_resize_req_0, ack => ptr_deref_1368_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1399_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp50_1384, dout => ptr_deref_1399_resized_base_address, req => ptr_deref_1399_base_resize_req_0, ack => ptr_deref_1399_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1407_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1366, dout => ptr_deref_1407_resized_base_address, req => ptr_deref_1407_base_resize_req_0, ack => ptr_deref_1407_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1416_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1366, dout => ptr_deref_1416_resized_base_address, req => ptr_deref_1416_base_resize_req_0, ack => ptr_deref_1416_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1421_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1366, dout => ptr_deref_1421_resized_base_address, req => ptr_deref_1421_base_resize_req_0, ack => ptr_deref_1421_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1438_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp44_1348, dout => ptr_deref_1438_resized_base_address, req => ptr_deref_1438_base_resize_req_0, ack => ptr_deref_1438_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1442_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp46_1362, dout => ptr_deref_1442_resized_base_address, req => ptr_deref_1442_base_resize_req_0, ack => ptr_deref_1442_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1458_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp46_1362, dout => ptr_deref_1458_resized_base_address, req => ptr_deref_1458_base_resize_req_0, ack => ptr_deref_1458_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1463_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp42_1334, dout => ptr_deref_1463_resized_base_address, req => ptr_deref_1463_base_resize_req_0, ack => ptr_deref_1463_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1482_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp60_1479, dout => ptr_deref_1482_resized_base_address, req => ptr_deref_1482_base_resize_req_0, ack => ptr_deref_1482_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1501_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp63_1498, dout => ptr_deref_1501_resized_base_address, req => ptr_deref_1501_base_resize_req_0, ack => ptr_deref_1501_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1533_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp66_1530, dout => ptr_deref_1533_resized_base_address, req => ptr_deref_1533_base_resize_req_0, ack => ptr_deref_1533_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1565_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp69_1562, dout => ptr_deref_1565_resized_base_address, req => ptr_deref_1565_base_resize_req_0, ack => ptr_deref_1565_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1094_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_1093_wire, dout => tmp_1095, req => type_cast_1094_inst_req_0, ack => type_cast_1094_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1098_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_1095, dout => tmp16_1099, req => type_cast_1098_inst_req_0, ack => type_cast_1098_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1109_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_1106, dout => tmp18_1110, req => type_cast_1109_inst_req_0, ack => type_cast_1109_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1177_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp23_1171, dout => type_cast_1177_wire, req => type_cast_1177_inst_req_0, ack => type_cast_1177_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1184_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp24_1174, dout => type_cast_1184_wire, req => type_cast_1184_inst_req_0, ack => type_cast_1184_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1199_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp24_1174, dout => type_cast_1199_wire, req => type_cast_1199_inst_req_0, ack => type_cast_1199_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1226_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp28_1220, dout => type_cast_1226_wire, req => type_cast_1226_inst_req_0, ack => type_cast_1226_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1244_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_1301, dout => type_cast_1244_wire, req => type_cast_1244_inst_req_0, ack => type_cast_1244_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1251_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp39_1289, dout => type_cast_1251_wire, req => type_cast_1251_inst_req_0, ack => type_cast_1251_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1292_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => scevgep1x_xix_xix_xix_xix_xi_1286, dout => type_cast_1292_wire, req => type_cast_1292_inst_req_0, ack => type_cast_1292_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1294_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp36_1248, dout => type_cast_1294_wire, req => type_cast_1294_inst_req_0, ack => type_cast_1294_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1347_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp43_1344, dout => tmp44_1348, req => type_cast_1347_inst_req_0, ack => type_cast_1347_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1361_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp45_1358, dout => tmp46_1362, req => type_cast_1361_inst_req_0, ack => type_cast_1361_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1365_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp39_1289, dout => tmp47_1366, req => type_cast_1365_inst_req_0, ack => type_cast_1365_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1374_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp39_1289, dout => tmp48_1375, req => type_cast_1374_inst_req_0, ack => type_cast_1374_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1570_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => tmp70_1566, dout => type_cast_1570_wire, req => type_cast_1570_inst_req_0, ack => type_cast_1570_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1585_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => tmp70_1566, dout => type_cast_1585_wire, req => type_cast_1585_inst_req_0, ack => type_cast_1585_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1626_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => tmp70_1566, dout => type_cast_1626_wire, req => type_cast_1626_inst_req_0, ack => type_cast_1626_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1667_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1095, dout => type_cast_1667_wire, req => type_cast_1667_inst_req_0, ack => type_cast_1667_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1673_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1095, dout => type_cast_1673_wire, req => type_cast_1673_inst_req_0, ack => type_cast_1673_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1679_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1095, dout => type_cast_1679_wire, req => type_cast_1679_inst_req_0, ack => type_cast_1679_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1685_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1095, dout => type_cast_1685_wire, req => type_cast_1685_inst_req_0, ack => type_cast_1685_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1691_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1095, dout => type_cast_1691_wire, req => type_cast_1691_inst_req_0, ack => type_cast_1691_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1123_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      array_obj_ref_1123_root_address_inst_ack_0 <= array_obj_ref_1123_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1123_final_offset;
      array_obj_ref_1123_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    array_obj_ref_1132_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      array_obj_ref_1132_root_address_inst_ack_0 <= array_obj_ref_1132_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1132_final_offset;
      array_obj_ref_1132_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    array_obj_ref_1260_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      array_obj_ref_1260_root_address_inst_ack_0 <= array_obj_ref_1260_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1260_final_offset;
      array_obj_ref_1260_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    array_obj_ref_1284_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      array_obj_ref_1284_root_address_inst_ack_0 <= array_obj_ref_1284_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1284_final_offset;
      array_obj_ref_1284_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    array_obj_ref_1477_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      array_obj_ref_1477_root_address_inst_ack_0 <= array_obj_ref_1477_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1477_final_offset;
      array_obj_ref_1477_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    array_obj_ref_1496_index_2_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1496_index_2_rename_ack_0 <= array_obj_ref_1496_index_2_rename_req_0;
      aggregated_sig <= simple_obj_ref_1495_resized;
      simple_obj_ref_1495_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1496_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1496_root_address_inst_ack_0 <= array_obj_ref_1496_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1496_final_offset;
      array_obj_ref_1496_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1528_index_2_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1528_index_2_rename_ack_0 <= array_obj_ref_1528_index_2_rename_req_0;
      aggregated_sig <= simple_obj_ref_1527_resized;
      simple_obj_ref_1527_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1528_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1528_root_address_inst_ack_0 <= array_obj_ref_1528_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1528_final_offset;
      array_obj_ref_1528_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1560_index_2_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1560_index_2_rename_ack_0 <= array_obj_ref_1560_index_2_rename_req_0;
      aggregated_sig <= simple_obj_ref_1559_resized;
      simple_obj_ref_1559_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1560_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1560_root_address_inst_ack_0 <= array_obj_ref_1560_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1560_final_offset;
      array_obj_ref_1560_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1113_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1113_gather_scatter_ack_0 <= ptr_deref_1113_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1113_data_3 & ptr_deref_1113_data_2 & ptr_deref_1113_data_1 & ptr_deref_1113_data_0;
      tmp19_1114 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1113_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1113_root_address_inst_ack_0 <= ptr_deref_1113_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1113_resized_base_address;
      ptr_deref_1113_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1137_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1137_addr_0_ack_0 <= ptr_deref_1137_addr_0_req_0;
      aggregated_sig <= ptr_deref_1137_root_address;
      ptr_deref_1137_word_address_0 <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1137_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1137_gather_scatter_ack_0 <= ptr_deref_1137_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1137_data_0;
      valx_xi4x_xix_xi_1138 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1137_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1137_root_address_inst_ack_0 <= ptr_deref_1137_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1137_resized_base_address;
      ptr_deref_1137_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1141_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1141_addr_0_ack_0 <= ptr_deref_1141_addr_0_req_0;
      aggregated_sig <= ptr_deref_1141_root_address;
      ptr_deref_1141_word_address_0 <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1141_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1141_gather_scatter_ack_0 <= ptr_deref_1141_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1141_data_0;
      val2x_xi6x_xix_xi_1142 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1141_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1141_root_address_inst_ack_0 <= ptr_deref_1141_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1141_resized_base_address;
      ptr_deref_1141_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1265_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1265_addr_0_ack_0 <= ptr_deref_1265_addr_0_req_0;
      aggregated_sig <= ptr_deref_1265_root_address;
      ptr_deref_1265_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1265_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1265_gather_scatter_ack_0 <= ptr_deref_1265_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1265_data_0;
      tmp37_1266 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1265_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1265_root_address_inst_ack_0 <= ptr_deref_1265_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1265_resized_base_address;
      ptr_deref_1265_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1336_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1336_addr_0_ack_0 <= ptr_deref_1336_addr_0_req_0;
      aggregated_sig <= ptr_deref_1336_root_address;
      ptr_deref_1336_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1336_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1336_gather_scatter_ack_0 <= ptr_deref_1336_gather_scatter_req_0;
      aggregated_sig <= type_cast_1338_wire_constant;
      ptr_deref_1336_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1336_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1336_root_address_inst_ack_0 <= ptr_deref_1336_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1336_resized_base_address;
      ptr_deref_1336_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1350_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1350_gather_scatter_ack_0 <= ptr_deref_1350_gather_scatter_req_0;
      aggregated_sig <= type_cast_1352_wire_constant;
      ptr_deref_1350_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1350_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1350_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1350_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1350_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1350_root_address_inst_ack_0 <= ptr_deref_1350_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1350_resized_base_address;
      ptr_deref_1350_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1368_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1368_gather_scatter_ack_0 <= ptr_deref_1368_gather_scatter_req_0;
      aggregated_sig <= type_cast_1370_wire_constant;
      ptr_deref_1368_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1368_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1368_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1368_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1368_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1368_root_address_inst_ack_0 <= ptr_deref_1368_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1368_resized_base_address;
      ptr_deref_1368_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1399_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1399_addr_0_ack_0 <= ptr_deref_1399_addr_0_req_0;
      aggregated_sig <= ptr_deref_1399_root_address;
      ptr_deref_1399_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1399_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1399_gather_scatter_ack_0 <= ptr_deref_1399_gather_scatter_req_0;
      aggregated_sig <= type_cast_1401_wire_constant;
      ptr_deref_1399_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1399_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1399_root_address_inst_ack_0 <= ptr_deref_1399_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1399_resized_base_address;
      ptr_deref_1399_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1407_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1407_gather_scatter_ack_0 <= ptr_deref_1407_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1407_data_3 & ptr_deref_1407_data_2 & ptr_deref_1407_data_1 & ptr_deref_1407_data_0;
      tmp52_1408 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1407_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1407_root_address_inst_ack_0 <= ptr_deref_1407_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1407_resized_base_address;
      ptr_deref_1407_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1416_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1416_gather_scatter_ack_0 <= ptr_deref_1416_gather_scatter_req_0;
      aggregated_sig <= tmp53_1414;
      ptr_deref_1416_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1416_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1416_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1416_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1416_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1416_root_address_inst_ack_0 <= ptr_deref_1416_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1416_resized_base_address;
      ptr_deref_1416_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1421_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1421_gather_scatter_ack_0 <= ptr_deref_1421_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1421_data_3 & ptr_deref_1421_data_2 & ptr_deref_1421_data_1 & ptr_deref_1421_data_0;
      tmp54_1422 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1421_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1421_root_address_inst_ack_0 <= ptr_deref_1421_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1421_resized_base_address;
      ptr_deref_1421_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1438_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1438_gather_scatter_ack_0 <= ptr_deref_1438_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1438_data_3 & ptr_deref_1438_data_2 & ptr_deref_1438_data_1 & ptr_deref_1438_data_0;
      tmp56_1439 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1438_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1438_root_address_inst_ack_0 <= ptr_deref_1438_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1438_resized_base_address;
      ptr_deref_1438_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1442_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1442_gather_scatter_ack_0 <= ptr_deref_1442_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1442_data_3 & ptr_deref_1442_data_2 & ptr_deref_1442_data_1 & ptr_deref_1442_data_0;
      tmp57_1443 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1442_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1442_root_address_inst_ack_0 <= ptr_deref_1442_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1442_resized_base_address;
      ptr_deref_1442_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1458_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1458_gather_scatter_ack_0 <= ptr_deref_1458_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1458_data_3 & ptr_deref_1458_data_2 & ptr_deref_1458_data_1 & ptr_deref_1458_data_0;
      tmp59_1459 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1458_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1458_root_address_inst_ack_0 <= ptr_deref_1458_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1458_resized_base_address;
      ptr_deref_1458_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1463_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1463_addr_0_ack_0 <= ptr_deref_1463_addr_0_req_0;
      aggregated_sig <= ptr_deref_1463_root_address;
      ptr_deref_1463_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1463_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1463_gather_scatter_ack_0 <= ptr_deref_1463_gather_scatter_req_0;
      aggregated_sig <= type_cast_1465_wire_constant;
      ptr_deref_1463_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1463_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1463_root_address_inst_ack_0 <= ptr_deref_1463_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1463_resized_base_address;
      ptr_deref_1463_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1482_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1482_addr_0_ack_0 <= ptr_deref_1482_addr_0_req_0;
      aggregated_sig <= ptr_deref_1482_root_address;
      ptr_deref_1482_word_address_0 <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1482_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1482_gather_scatter_ack_0 <= ptr_deref_1482_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1482_data_0;
      tmp61_1483 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1482_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1482_root_address_inst_ack_0 <= ptr_deref_1482_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1482_resized_base_address;
      ptr_deref_1482_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1501_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1501_addr_0_ack_0 <= ptr_deref_1501_addr_0_req_0;
      aggregated_sig <= ptr_deref_1501_root_address;
      ptr_deref_1501_word_address_0 <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1501_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1501_gather_scatter_ack_0 <= ptr_deref_1501_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1501_data_0;
      tmp64_1502 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1501_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1501_root_address_inst_ack_0 <= ptr_deref_1501_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1501_resized_base_address;
      ptr_deref_1501_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1533_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1533_addr_0_ack_0 <= ptr_deref_1533_addr_0_req_0;
      aggregated_sig <= ptr_deref_1533_root_address;
      ptr_deref_1533_word_address_0 <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1533_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1533_gather_scatter_ack_0 <= ptr_deref_1533_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1533_data_0;
      tmp67_1534 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1533_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1533_root_address_inst_ack_0 <= ptr_deref_1533_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1533_resized_base_address;
      ptr_deref_1533_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1565_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1565_addr_0_ack_0 <= ptr_deref_1565_addr_0_req_0;
      aggregated_sig <= ptr_deref_1565_root_address;
      ptr_deref_1565_word_address_0 <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1565_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1565_gather_scatter_ack_0 <= ptr_deref_1565_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1565_data_0;
      tmp70_1566 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1565_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1565_root_address_inst_ack_0 <= ptr_deref_1565_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1565_resized_base_address;
      ptr_deref_1565_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    simple_obj_ref_1213_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1213_gather_scatter_ack_0 <= simple_obj_ref_1213_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_1213_data_0;
      tmp27_1214 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1221_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1221_gather_scatter_ack_0 <= simple_obj_ref_1221_gather_scatter_req_0;
      aggregated_sig <= tmp28_1220;
      simple_obj_ref_1221_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_1159_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp22_1158;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1159_branch_req_0,
          ack0 => if_stmt_1159_branch_ack_0,
          ack1 => if_stmt_1159_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1190_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp25_1189;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1190_branch_req_0,
          ack0 => if_stmt_1190_branch_ack_0,
          ack1 => if_stmt_1190_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1205_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp26_1204;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1205_branch_req_0,
          ack0 => if_stmt_1205_branch_ack_0,
          ack1 => if_stmt_1205_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1232_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp29_1231;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1232_branch_req_0,
          ack0 => if_stmt_1232_branch_ack_0,
          ack1 => if_stmt_1232_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1273_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp38_1272;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1273_branch_req_0,
          ack0 => if_stmt_1273_branch_ack_0,
          ack1 => if_stmt_1273_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1308_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1307;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1308_branch_req_0,
          ack0 => if_stmt_1308_branch_ack_0,
          ack1 => if_stmt_1308_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1321_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp41_1320;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1321_branch_req_0,
          ack0 => if_stmt_1321_branch_ack_0,
          ack1 => if_stmt_1321_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1391_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp51_1390;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1391_branch_req_0,
          ack0 => if_stmt_1391_branch_ack_0,
          ack1 => if_stmt_1391_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1429_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp55_1428;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1429_branch_req_0,
          ack0 => if_stmt_1429_branch_ack_0,
          ack1 => if_stmt_1429_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1449_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp58_1448;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1449_branch_req_0,
          ack0 => if_stmt_1449_branch_ack_0,
          ack1 => if_stmt_1449_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1509_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp65_1508;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1509_branch_req_0,
          ack0 => if_stmt_1509_branch_ack_0,
          ack1 => if_stmt_1509_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1541_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp68_1540;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1541_branch_req_0,
          ack0 => if_stmt_1541_branch_ack_0,
          ack1 => if_stmt_1541_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1576_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= Pivot15_1575;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1576_branch_req_0,
          ack0 => if_stmt_1576_branch_ack_0,
          ack1 => if_stmt_1576_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1591_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= Pivot13_1590;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1591_branch_req_0,
          ack0 => if_stmt_1591_branch_ack_0,
          ack1 => if_stmt_1591_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1604_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf11_1603;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1604_branch_req_0,
          ack0 => if_stmt_1604_branch_ack_0,
          ack1 => if_stmt_1604_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1617_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf9_1616;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1617_branch_req_0,
          ack0 => if_stmt_1617_branch_ack_0,
          ack1 => if_stmt_1617_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1632_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= Pivot_1631;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1632_branch_req_0,
          ack0 => if_stmt_1632_branch_ack_0,
          ack1 => if_stmt_1632_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1645_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf7_1644;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1645_branch_req_0,
          ack0 => if_stmt_1645_branch_ack_0,
          ack1 => if_stmt_1645_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1658_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf_1657;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1658_branch_req_0,
          ack0 => if_stmt_1658_branch_ack_0,
          ack1 => if_stmt_1658_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1105_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1105_resized_base_address;
      array_obj_ref_1105_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1105_root_address_inst_req_0,
          ackL => array_obj_ref_1105_root_address_inst_ack_0,
          reqR => array_obj_ref_1105_root_address_inst_req_1,
          ackR => array_obj_ref_1105_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1477_index_0_scale array_obj_ref_1123_index_0_scale array_obj_ref_1132_index_0_scale 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1474_resized & simple_obj_ref_1118_resized & simple_obj_ref_1127_resized;
      simple_obj_ref_1474_scaled <= data_out(14 downto 10);
      simple_obj_ref_1118_scaled <= data_out(9 downto 5);
      simple_obj_ref_1127_scaled <= data_out(4 downto 0);
      reqL(2) <= array_obj_ref_1477_index_0_scale_req_0;
      reqL(1) <= array_obj_ref_1123_index_0_scale_req_0;
      reqL(0) <= array_obj_ref_1132_index_0_scale_req_0;
      array_obj_ref_1477_index_0_scale_ack_0 <= ackL(2);
      array_obj_ref_1123_index_0_scale_ack_0 <= ackL(1);
      array_obj_ref_1132_index_0_scale_ack_0 <= ackL(0);
      reqR(2) <= array_obj_ref_1477_index_0_scale_req_1;
      reqR(1) <= array_obj_ref_1123_index_0_scale_req_1;
      reqR(0) <= array_obj_ref_1132_index_0_scale_req_1;
      array_obj_ref_1477_index_0_scale_ack_1 <= ackR(2);
      array_obj_ref_1123_index_0_scale_ack_1 <= ackR(1);
      array_obj_ref_1132_index_0_scale_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00101",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 3--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1123_index_sum_1 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(4 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1118_scaled;
      array_obj_ref_1123_index_partial_sum_1 <= data_out(4 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00000",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1123_index_sum_1_req_0,
          ackL => array_obj_ref_1123_index_sum_1_ack_0,
          reqR => array_obj_ref_1123_index_sum_1_req_1,
          ackR => array_obj_ref_1123_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1132_index_sum_1 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(4 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1127_scaled;
      array_obj_ref_1132_index_partial_sum_1 <= data_out(4 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00001",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1132_index_sum_1_req_0,
          ackL => array_obj_ref_1132_index_sum_1_ack_0,
          reqR => array_obj_ref_1132_index_sum_1_req_1,
          ackR => array_obj_ref_1132_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1260_index_0_scale array_obj_ref_1284_index_0_scale 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(27 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1257_resized & simple_obj_ref_1281_resized;
      simple_obj_ref_1257_scaled <= data_out(27 downto 14);
      simple_obj_ref_1281_scaled <= data_out(13 downto 0);
      reqL(1) <= array_obj_ref_1260_index_0_scale_req_0;
      reqL(0) <= array_obj_ref_1284_index_0_scale_req_0;
      array_obj_ref_1260_index_0_scale_ack_0 <= ackL(1);
      array_obj_ref_1284_index_0_scale_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1260_index_0_scale_req_1;
      reqR(0) <= array_obj_ref_1284_index_0_scale_req_1;
      array_obj_ref_1260_index_0_scale_ack_1 <= ackR(1);
      array_obj_ref_1284_index_0_scale_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000010000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1260_index_sum_1 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1257_scaled;
      array_obj_ref_1260_index_partial_sum_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1260_index_sum_1_req_0,
          ackL => array_obj_ref_1260_index_sum_1_ack_0,
          reqR => array_obj_ref_1260_index_sum_1_req_1,
          ackR => array_obj_ref_1260_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1284_index_sum_1 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1281_scaled;
      array_obj_ref_1284_index_partial_sum_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1284_index_sum_1_req_0,
          ackL => array_obj_ref_1284_index_sum_1_ack_0,
          reqR => array_obj_ref_1284_index_sum_1_req_1,
          ackR => array_obj_ref_1284_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1333_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1333_final_offset & array_obj_ref_1333_resized_base_address;
      array_obj_ref_1333_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 14, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1333_root_address_inst_req_0,
          ackL => array_obj_ref_1333_root_address_inst_ack_0,
          reqR => array_obj_ref_1333_root_address_inst_req_1,
          ackR => array_obj_ref_1333_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1343_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1343_resized_base_address;
      array_obj_ref_1343_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000100",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1343_root_address_inst_req_0,
          ackL => array_obj_ref_1343_root_address_inst_ack_0,
          reqR => array_obj_ref_1343_root_address_inst_req_1,
          ackR => array_obj_ref_1343_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1357_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1357_resized_base_address;
      array_obj_ref_1357_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000001000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1357_root_address_inst_req_0,
          ackL => array_obj_ref_1357_root_address_inst_ack_0,
          reqR => array_obj_ref_1357_root_address_inst_req_1,
          ackR => array_obj_ref_1357_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1383_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1383_resized_base_address;
      array_obj_ref_1383_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000001100",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1383_root_address_inst_req_0,
          ackL => array_obj_ref_1383_root_address_inst_ack_0,
          reqR => array_obj_ref_1383_root_address_inst_req_1,
          ackR => array_obj_ref_1383_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1477_index_sum_1 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(4 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1474_scaled;
      array_obj_ref_1477_index_partial_sum_1 <= data_out(4 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00011",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1477_index_sum_1_req_0,
          ackL => array_obj_ref_1477_index_sum_1_ack_0,
          reqR => array_obj_ref_1477_index_sum_1_req_1,
          ackR => array_obj_ref_1477_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1496_index_sum_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1495_scaled;
      array_obj_ref_1496_index_partial_sum_1 <= data_out(8 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1496_index_sum_1_req_0,
          ackL => array_obj_ref_1496_index_sum_1_ack_0,
          reqR => array_obj_ref_1496_index_sum_1_req_1,
          ackR => array_obj_ref_1496_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_1528_index_sum_1 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1527_scaled;
      array_obj_ref_1528_index_partial_sum_1 <= data_out(8 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1528_index_sum_1_req_0,
          ackL => array_obj_ref_1528_index_sum_1_ack_0,
          reqR => array_obj_ref_1528_index_sum_1_req_1,
          ackR => array_obj_ref_1528_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_1560_index_sum_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1559_scaled;
      array_obj_ref_1560_index_partial_sum_1 <= data_out(8 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1560_index_sum_1_req_0,
          ackL => array_obj_ref_1560_index_sum_1_ack_0,
          reqR => array_obj_ref_1560_index_sum_1_req_1,
          ackR => array_obj_ref_1560_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1146_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= valx_xi4x_xix_xi_1138 & tmp19_1114;
      tmp20_1147 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1146_inst_req_0,
          ackL => binary_1146_inst_ack_0,
          reqR => binary_1146_inst_req_1,
          ackR => binary_1146_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1151_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_1147 & val2x_xi6x_xix_xi_1142;
      tmp21_1152 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1151_inst_req_0,
          ackL => binary_1151_inst_ack_0,
          reqR => binary_1151_inst_req_1,
          ackR => binary_1151_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1427_inst binary_1157_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp54_1422 & tmp21_1152;
      tmp55_1428 <= data_out(1 downto 1);
      tmp22_1158 <= data_out(0 downto 0);
      reqL(1) <= binary_1427_inst_req_0;
      reqL(0) <= binary_1157_inst_req_0;
      binary_1427_inst_ack_0 <= ackL(1);
      binary_1157_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1427_inst_req_1;
      reqR(0) <= binary_1157_inst_req_1;
      binary_1427_inst_ack_1 <= ackR(1);
      binary_1157_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1170_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp24_1174;
      tmp23_1171 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1170_inst_req_0,
          ackL => binary_1170_inst_ack_0,
          reqR => binary_1170_inst_req_1,
          ackR => binary_1170_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1188_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1184_wire;
      tmp25_1189 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1188_inst_req_0,
          ackL => binary_1188_inst_ack_0,
          reqR => binary_1188_inst_req_1,
          ackR => binary_1188_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1203_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1199_wire;
      tmp26_1204 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1203_inst_req_0,
          ackL => binary_1203_inst_ack_0,
          reqR => binary_1203_inst_req_1,
          ackR => binary_1203_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1219_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp27_1214;
      tmp28_1220 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1219_inst_req_0,
          ackL => binary_1219_inst_ack_0,
          reqR => binary_1219_inst_req_1,
          ackR => binary_1219_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1230_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1226_wire;
      tmp29_1231 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1230_inst_req_0,
          ackL => binary_1230_inst_ack_0,
          reqR => binary_1230_inst_req_1,
          ackR => binary_1230_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1271_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp37_1266;
      tmp38_1272 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1271_inst_req_0,
          ackL => binary_1271_inst_ack_0,
          reqR => binary_1271_inst_req_1,
          ackR => binary_1271_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1300_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp35_1241;
      tmp40_1301 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1300_inst_req_0,
          ackL => binary_1300_inst_ack_0,
          reqR => binary_1300_inst_req_1,
          ackR => binary_1300_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1306_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp40_1301;
      exitcond_1307 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1306_inst_req_0,
          ackL => binary_1306_inst_ack_0,
          reqR => binary_1306_inst_req_1,
          ackR => binary_1306_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1319_inst binary_1389_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp39_1289 & tmp50_1384;
      tmp41_1320 <= data_out(1 downto 1);
      tmp51_1390 <= data_out(0 downto 0);
      reqL(1) <= binary_1319_inst_req_0;
      reqL(0) <= binary_1389_inst_req_0;
      binary_1319_inst_ack_0 <= ackL(1);
      binary_1389_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1319_inst_req_1;
      reqR(0) <= binary_1389_inst_req_1;
      binary_1319_inst_ack_1 <= ackR(1);
      binary_1389_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_1413_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp52_1408;
      tmp53_1414 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1413_inst_req_0,
          ackL => binary_1413_inst_ack_0,
          reqR => binary_1413_inst_req_1,
          ackR => binary_1413_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_1447_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp56_1439 & tmp57_1443;
      tmp58_1448 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1447_inst_req_0,
          ackL => binary_1447_inst_ack_0,
          reqR => binary_1447_inst_req_1,
          ackR => binary_1447_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_1488_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp61_1483;
      tmp62_1489 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000001001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1488_inst_req_0,
          ackL => binary_1488_inst_ack_0,
          reqR => binary_1488_inst_req_1,
          ackR => binary_1488_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_1507_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp64_1502;
      tmp65_1508 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01110100",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1507_inst_req_0,
          ackL => binary_1507_inst_ack_0,
          reqR => binary_1507_inst_req_1,
          ackR => binary_1507_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_1520_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp62_1489;
      xx_xsum26x_xi_1521 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1520_inst_req_0,
          ackL => binary_1520_inst_ack_0,
          reqR => binary_1520_inst_req_1,
          ackR => binary_1520_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_1539_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp67_1534;
      tmp68_1540 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01101111",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1539_inst_req_0,
          ackL => binary_1539_inst_ack_0,
          reqR => binary_1539_inst_req_1,
          ackR => binary_1539_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_1552_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp62_1489;
      xx_xsum27x_xi_1553 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1552_inst_req_0,
          ackL => binary_1552_inst_ack_0,
          reqR => binary_1552_inst_req_1,
          ackR => binary_1552_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_1574_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1570_wire;
      Pivot15_1575 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1574_inst_req_0,
          ackL => binary_1574_inst_ack_0,
          reqR => binary_1574_inst_req_1,
          ackR => binary_1574_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_1589_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1585_wire;
      Pivot13_1590 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1589_inst_req_0,
          ackL => binary_1589_inst_ack_0,
          reqR => binary_1589_inst_req_1,
          ackR => binary_1589_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_1602_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_1566;
      SwitchLeaf11_1603 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1602_inst_req_0,
          ackL => binary_1602_inst_ack_0,
          reqR => binary_1602_inst_req_1,
          ackR => binary_1602_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_1615_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_1566;
      SwitchLeaf9_1616 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1615_inst_req_0,
          ackL => binary_1615_inst_ack_0,
          reqR => binary_1615_inst_req_1,
          ackR => binary_1615_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_1630_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1626_wire;
      Pivot_1631 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1630_inst_req_0,
          ackL => binary_1630_inst_ack_0,
          reqR => binary_1630_inst_req_1,
          ackR => binary_1630_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_1643_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_1566;
      SwitchLeaf7_1644 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1643_inst_req_0,
          ackL => binary_1643_inst_ack_0,
          reqR => binary_1643_inst_req_1,
          ackR => binary_1643_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_1656_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_1566;
      SwitchLeaf_1657 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110000",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1656_inst_req_0,
          ackL => binary_1656_inst_ack_0,
          reqR => binary_1656_inst_req_1,
          ackR => binary_1656_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : ptr_deref_1113_addr_0 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1113_root_address;
      ptr_deref_1113_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1113_addr_0_req_0,
          ackL => ptr_deref_1113_addr_0_ack_0,
          reqR => ptr_deref_1113_addr_0_req_1,
          ackR => ptr_deref_1113_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : ptr_deref_1113_addr_1 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1113_root_address;
      ptr_deref_1113_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1113_addr_1_req_0,
          ackL => ptr_deref_1113_addr_1_ack_0,
          reqR => ptr_deref_1113_addr_1_req_1,
          ackR => ptr_deref_1113_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : ptr_deref_1113_addr_2 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1113_root_address;
      ptr_deref_1113_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1113_addr_2_req_0,
          ackL => ptr_deref_1113_addr_2_ack_0,
          reqR => ptr_deref_1113_addr_2_req_1,
          ackR => ptr_deref_1113_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : ptr_deref_1113_addr_3 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1113_root_address;
      ptr_deref_1113_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1113_addr_3_req_0,
          ackL => ptr_deref_1113_addr_3_ack_0,
          reqR => ptr_deref_1113_addr_3_req_1,
          ackR => ptr_deref_1113_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : ptr_deref_1350_addr_0 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1350_root_address;
      ptr_deref_1350_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1350_addr_0_req_0,
          ackL => ptr_deref_1350_addr_0_ack_0,
          reqR => ptr_deref_1350_addr_0_req_1,
          ackR => ptr_deref_1350_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : ptr_deref_1350_addr_1 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1350_root_address;
      ptr_deref_1350_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1350_addr_1_req_0,
          ackL => ptr_deref_1350_addr_1_ack_0,
          reqR => ptr_deref_1350_addr_1_req_1,
          ackR => ptr_deref_1350_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : ptr_deref_1350_addr_2 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1350_root_address;
      ptr_deref_1350_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1350_addr_2_req_0,
          ackL => ptr_deref_1350_addr_2_ack_0,
          reqR => ptr_deref_1350_addr_2_req_1,
          ackR => ptr_deref_1350_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : ptr_deref_1350_addr_3 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1350_root_address;
      ptr_deref_1350_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1350_addr_3_req_0,
          ackL => ptr_deref_1350_addr_3_ack_0,
          reqR => ptr_deref_1350_addr_3_req_1,
          ackR => ptr_deref_1350_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : ptr_deref_1368_addr_0 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1368_root_address;
      ptr_deref_1368_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1368_addr_0_req_0,
          ackL => ptr_deref_1368_addr_0_ack_0,
          reqR => ptr_deref_1368_addr_0_req_1,
          ackR => ptr_deref_1368_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : ptr_deref_1368_addr_1 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1368_root_address;
      ptr_deref_1368_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1368_addr_1_req_0,
          ackL => ptr_deref_1368_addr_1_ack_0,
          reqR => ptr_deref_1368_addr_1_req_1,
          ackR => ptr_deref_1368_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : ptr_deref_1368_addr_2 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1368_root_address;
      ptr_deref_1368_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1368_addr_2_req_0,
          ackL => ptr_deref_1368_addr_2_ack_0,
          reqR => ptr_deref_1368_addr_2_req_1,
          ackR => ptr_deref_1368_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_1368_addr_3 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1368_root_address;
      ptr_deref_1368_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1368_addr_3_req_0,
          ackL => ptr_deref_1368_addr_3_ack_0,
          reqR => ptr_deref_1368_addr_3_req_1,
          ackR => ptr_deref_1368_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_1407_addr_0 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1407_root_address;
      ptr_deref_1407_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1407_addr_0_req_0,
          ackL => ptr_deref_1407_addr_0_ack_0,
          reqR => ptr_deref_1407_addr_0_req_1,
          ackR => ptr_deref_1407_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_1407_addr_1 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1407_root_address;
      ptr_deref_1407_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1407_addr_1_req_0,
          ackL => ptr_deref_1407_addr_1_ack_0,
          reqR => ptr_deref_1407_addr_1_req_1,
          ackR => ptr_deref_1407_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_1407_addr_2 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1407_root_address;
      ptr_deref_1407_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1407_addr_2_req_0,
          ackL => ptr_deref_1407_addr_2_ack_0,
          reqR => ptr_deref_1407_addr_2_req_1,
          ackR => ptr_deref_1407_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_1407_addr_3 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1407_root_address;
      ptr_deref_1407_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1407_addr_3_req_0,
          ackL => ptr_deref_1407_addr_3_ack_0,
          reqR => ptr_deref_1407_addr_3_req_1,
          ackR => ptr_deref_1407_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_1416_addr_0 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1416_root_address;
      ptr_deref_1416_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1416_addr_0_req_0,
          ackL => ptr_deref_1416_addr_0_ack_0,
          reqR => ptr_deref_1416_addr_0_req_1,
          ackR => ptr_deref_1416_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_1416_addr_1 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1416_root_address;
      ptr_deref_1416_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1416_addr_1_req_0,
          ackL => ptr_deref_1416_addr_1_ack_0,
          reqR => ptr_deref_1416_addr_1_req_1,
          ackR => ptr_deref_1416_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : ptr_deref_1416_addr_2 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1416_root_address;
      ptr_deref_1416_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1416_addr_2_req_0,
          ackL => ptr_deref_1416_addr_2_ack_0,
          reqR => ptr_deref_1416_addr_2_req_1,
          ackR => ptr_deref_1416_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : ptr_deref_1416_addr_3 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1416_root_address;
      ptr_deref_1416_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1416_addr_3_req_0,
          ackL => ptr_deref_1416_addr_3_ack_0,
          reqR => ptr_deref_1416_addr_3_req_1,
          ackR => ptr_deref_1416_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : ptr_deref_1421_addr_0 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1421_root_address;
      ptr_deref_1421_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1421_addr_0_req_0,
          ackL => ptr_deref_1421_addr_0_ack_0,
          reqR => ptr_deref_1421_addr_0_req_1,
          ackR => ptr_deref_1421_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : ptr_deref_1421_addr_1 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1421_root_address;
      ptr_deref_1421_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1421_addr_1_req_0,
          ackL => ptr_deref_1421_addr_1_ack_0,
          reqR => ptr_deref_1421_addr_1_req_1,
          ackR => ptr_deref_1421_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : ptr_deref_1421_addr_2 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1421_root_address;
      ptr_deref_1421_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1421_addr_2_req_0,
          ackL => ptr_deref_1421_addr_2_ack_0,
          reqR => ptr_deref_1421_addr_2_req_1,
          ackR => ptr_deref_1421_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : ptr_deref_1421_addr_3 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1421_root_address;
      ptr_deref_1421_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1421_addr_3_req_0,
          ackL => ptr_deref_1421_addr_3_ack_0,
          reqR => ptr_deref_1421_addr_3_req_1,
          ackR => ptr_deref_1421_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : ptr_deref_1438_addr_0 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1438_root_address;
      ptr_deref_1438_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1438_addr_0_req_0,
          ackL => ptr_deref_1438_addr_0_ack_0,
          reqR => ptr_deref_1438_addr_0_req_1,
          ackR => ptr_deref_1438_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : ptr_deref_1438_addr_1 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1438_root_address;
      ptr_deref_1438_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1438_addr_1_req_0,
          ackL => ptr_deref_1438_addr_1_ack_0,
          reqR => ptr_deref_1438_addr_1_req_1,
          ackR => ptr_deref_1438_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : ptr_deref_1438_addr_2 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1438_root_address;
      ptr_deref_1438_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1438_addr_2_req_0,
          ackL => ptr_deref_1438_addr_2_ack_0,
          reqR => ptr_deref_1438_addr_2_req_1,
          ackR => ptr_deref_1438_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : ptr_deref_1438_addr_3 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1438_root_address;
      ptr_deref_1438_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1438_addr_3_req_0,
          ackL => ptr_deref_1438_addr_3_ack_0,
          reqR => ptr_deref_1438_addr_3_req_1,
          ackR => ptr_deref_1438_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : ptr_deref_1442_addr_0 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1442_root_address;
      ptr_deref_1442_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1442_addr_0_req_0,
          ackL => ptr_deref_1442_addr_0_ack_0,
          reqR => ptr_deref_1442_addr_0_req_1,
          ackR => ptr_deref_1442_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : ptr_deref_1442_addr_1 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1442_root_address;
      ptr_deref_1442_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1442_addr_1_req_0,
          ackL => ptr_deref_1442_addr_1_ack_0,
          reqR => ptr_deref_1442_addr_1_req_1,
          ackR => ptr_deref_1442_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : ptr_deref_1442_addr_2 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1442_root_address;
      ptr_deref_1442_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1442_addr_2_req_0,
          ackL => ptr_deref_1442_addr_2_ack_0,
          reqR => ptr_deref_1442_addr_2_req_1,
          ackR => ptr_deref_1442_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : ptr_deref_1442_addr_3 
    SplitOperatorGroup72: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1442_root_address;
      ptr_deref_1442_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1442_addr_3_req_0,
          ackL => ptr_deref_1442_addr_3_ack_0,
          reqR => ptr_deref_1442_addr_3_req_1,
          ackR => ptr_deref_1442_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : ptr_deref_1458_addr_0 
    SplitOperatorGroup73: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1458_root_address;
      ptr_deref_1458_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1458_addr_0_req_0,
          ackL => ptr_deref_1458_addr_0_ack_0,
          reqR => ptr_deref_1458_addr_0_req_1,
          ackR => ptr_deref_1458_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : ptr_deref_1458_addr_1 
    SplitOperatorGroup74: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1458_root_address;
      ptr_deref_1458_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1458_addr_1_req_0,
          ackL => ptr_deref_1458_addr_1_ack_0,
          reqR => ptr_deref_1458_addr_1_req_1,
          ackR => ptr_deref_1458_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : ptr_deref_1458_addr_2 
    SplitOperatorGroup75: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1458_root_address;
      ptr_deref_1458_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1458_addr_2_req_0,
          ackL => ptr_deref_1458_addr_2_ack_0,
          reqR => ptr_deref_1458_addr_2_req_1,
          ackR => ptr_deref_1458_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : ptr_deref_1458_addr_3 
    SplitOperatorGroup76: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1458_root_address;
      ptr_deref_1458_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1458_addr_3_req_0,
          ackL => ptr_deref_1458_addr_3_ack_0,
          reqR => ptr_deref_1458_addr_3_req_1,
          ackR => ptr_deref_1458_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared load operator group (0) : ptr_deref_1113_load_0 ptr_deref_1113_load_1 ptr_deref_1113_load_2 ptr_deref_1113_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1113_load_0_req_0,
        ptr_deref_1113_load_0_ack_0,
        ptr_deref_1113_load_0_req_1,
        ptr_deref_1113_load_0_ack_1,
        "ptr_deref_1113_load_0",
        "memory_space_5" ,
        ptr_deref_1113_data_0,
        ptr_deref_1113_word_address_0,
        "ptr_deref_1113_data_0",
        "ptr_deref_1113_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1113_load_1_req_0,
        ptr_deref_1113_load_1_ack_0,
        ptr_deref_1113_load_1_req_1,
        ptr_deref_1113_load_1_ack_1,
        "ptr_deref_1113_load_1",
        "memory_space_5" ,
        ptr_deref_1113_data_1,
        ptr_deref_1113_word_address_1,
        "ptr_deref_1113_data_1",
        "ptr_deref_1113_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1113_load_2_req_0,
        ptr_deref_1113_load_2_ack_0,
        ptr_deref_1113_load_2_req_1,
        ptr_deref_1113_load_2_ack_1,
        "ptr_deref_1113_load_2",
        "memory_space_5" ,
        ptr_deref_1113_data_2,
        ptr_deref_1113_word_address_2,
        "ptr_deref_1113_data_2",
        "ptr_deref_1113_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1113_load_3_req_0,
        ptr_deref_1113_load_3_ack_0,
        ptr_deref_1113_load_3_req_1,
        ptr_deref_1113_load_3_ack_1,
        "ptr_deref_1113_load_3",
        "memory_space_5" ,
        ptr_deref_1113_data_3,
        ptr_deref_1113_word_address_3,
        "ptr_deref_1113_data_3",
        "ptr_deref_1113_word_address_3" -- 
      );
      reqL(3) <= ptr_deref_1113_load_0_req_0;
      reqL(2) <= ptr_deref_1113_load_1_req_0;
      reqL(1) <= ptr_deref_1113_load_2_req_0;
      reqL(0) <= ptr_deref_1113_load_3_req_0;
      ptr_deref_1113_load_0_ack_0 <= ackL(3);
      ptr_deref_1113_load_1_ack_0 <= ackL(2);
      ptr_deref_1113_load_2_ack_0 <= ackL(1);
      ptr_deref_1113_load_3_ack_0 <= ackL(0);
      reqR(3) <= ptr_deref_1113_load_0_req_1;
      reqR(2) <= ptr_deref_1113_load_1_req_1;
      reqR(1) <= ptr_deref_1113_load_2_req_1;
      reqR(0) <= ptr_deref_1113_load_3_req_1;
      ptr_deref_1113_load_0_ack_1 <= ackR(3);
      ptr_deref_1113_load_1_ack_1 <= ackR(2);
      ptr_deref_1113_load_2_ack_1 <= ackR(1);
      ptr_deref_1113_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_1113_word_address_0 & ptr_deref_1113_word_address_1 & ptr_deref_1113_word_address_2 & ptr_deref_1113_word_address_3;
      ptr_deref_1113_data_0 <= data_out(31 downto 24);
      ptr_deref_1113_data_1 <= data_out(23 downto 16);
      ptr_deref_1113_data_2 <= data_out(15 downto 8);
      ptr_deref_1113_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 4,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 4,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1482_load_0 ptr_deref_1137_load_0 ptr_deref_1141_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1482_load_0_req_0,
        ptr_deref_1482_load_0_ack_0,
        ptr_deref_1482_load_0_req_1,
        ptr_deref_1482_load_0_ack_1,
        "ptr_deref_1482_load_0",
        "memory_space_2" ,
        ptr_deref_1482_data_0,
        ptr_deref_1482_word_address_0,
        "ptr_deref_1482_data_0",
        "ptr_deref_1482_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1137_load_0_req_0,
        ptr_deref_1137_load_0_ack_0,
        ptr_deref_1137_load_0_req_1,
        ptr_deref_1137_load_0_ack_1,
        "ptr_deref_1137_load_0",
        "memory_space_2" ,
        ptr_deref_1137_data_0,
        ptr_deref_1137_word_address_0,
        "ptr_deref_1137_data_0",
        "ptr_deref_1137_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1141_load_0_req_0,
        ptr_deref_1141_load_0_ack_0,
        ptr_deref_1141_load_0_req_1,
        ptr_deref_1141_load_0_ack_1,
        "ptr_deref_1141_load_0",
        "memory_space_2" ,
        ptr_deref_1141_data_0,
        ptr_deref_1141_word_address_0,
        "ptr_deref_1141_data_0",
        "ptr_deref_1141_word_address_0" -- 
      );
      reqL(2) <= ptr_deref_1482_load_0_req_0;
      reqL(1) <= ptr_deref_1137_load_0_req_0;
      reqL(0) <= ptr_deref_1141_load_0_req_0;
      ptr_deref_1482_load_0_ack_0 <= ackL(2);
      ptr_deref_1137_load_0_ack_0 <= ackL(1);
      ptr_deref_1141_load_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1482_load_0_req_1;
      reqR(1) <= ptr_deref_1137_load_0_req_1;
      reqR(0) <= ptr_deref_1141_load_0_req_1;
      ptr_deref_1482_load_0_ack_1 <= ackR(2);
      ptr_deref_1137_load_0_ack_1 <= ackR(1);
      ptr_deref_1141_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1482_word_address_0 & ptr_deref_1137_word_address_0 & ptr_deref_1141_word_address_0;
      ptr_deref_1482_data_0 <= data_out(95 downto 64);
      ptr_deref_1137_data_0 <= data_out(63 downto 32);
      ptr_deref_1141_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 5,
        num_reqs => 3,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(4 downto 0),
          mtag => memory_space_2_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1421_load_1 ptr_deref_1458_load_0 ptr_deref_1265_load_0 ptr_deref_1421_load_0 ptr_deref_1407_load_0 ptr_deref_1442_load_3 ptr_deref_1458_load_1 ptr_deref_1458_load_3 ptr_deref_1442_load_0 ptr_deref_1442_load_2 ptr_deref_1458_load_2 ptr_deref_1407_load_2 ptr_deref_1442_load_1 ptr_deref_1407_load_3 ptr_deref_1407_load_1 ptr_deref_1438_load_3 ptr_deref_1438_load_2 ptr_deref_1438_load_1 ptr_deref_1438_load_0 ptr_deref_1421_load_3 ptr_deref_1421_load_2 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(293 downto 0);
      signal data_out: std_logic_vector(167 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 20 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1421_load_1_req_0,
        ptr_deref_1421_load_1_ack_0,
        ptr_deref_1421_load_1_req_1,
        ptr_deref_1421_load_1_ack_1,
        "ptr_deref_1421_load_1",
        "memory_space_3" ,
        ptr_deref_1421_data_1,
        ptr_deref_1421_word_address_1,
        "ptr_deref_1421_data_1",
        "ptr_deref_1421_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1458_load_0_req_0,
        ptr_deref_1458_load_0_ack_0,
        ptr_deref_1458_load_0_req_1,
        ptr_deref_1458_load_0_ack_1,
        "ptr_deref_1458_load_0",
        "memory_space_3" ,
        ptr_deref_1458_data_0,
        ptr_deref_1458_word_address_0,
        "ptr_deref_1458_data_0",
        "ptr_deref_1458_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1265_load_0_req_0,
        ptr_deref_1265_load_0_ack_0,
        ptr_deref_1265_load_0_req_1,
        ptr_deref_1265_load_0_ack_1,
        "ptr_deref_1265_load_0",
        "memory_space_3" ,
        ptr_deref_1265_data_0,
        ptr_deref_1265_word_address_0,
        "ptr_deref_1265_data_0",
        "ptr_deref_1265_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1421_load_0_req_0,
        ptr_deref_1421_load_0_ack_0,
        ptr_deref_1421_load_0_req_1,
        ptr_deref_1421_load_0_ack_1,
        "ptr_deref_1421_load_0",
        "memory_space_3" ,
        ptr_deref_1421_data_0,
        ptr_deref_1421_word_address_0,
        "ptr_deref_1421_data_0",
        "ptr_deref_1421_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1407_load_0_req_0,
        ptr_deref_1407_load_0_ack_0,
        ptr_deref_1407_load_0_req_1,
        ptr_deref_1407_load_0_ack_1,
        "ptr_deref_1407_load_0",
        "memory_space_3" ,
        ptr_deref_1407_data_0,
        ptr_deref_1407_word_address_0,
        "ptr_deref_1407_data_0",
        "ptr_deref_1407_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1442_load_3_req_0,
        ptr_deref_1442_load_3_ack_0,
        ptr_deref_1442_load_3_req_1,
        ptr_deref_1442_load_3_ack_1,
        "ptr_deref_1442_load_3",
        "memory_space_3" ,
        ptr_deref_1442_data_3,
        ptr_deref_1442_word_address_3,
        "ptr_deref_1442_data_3",
        "ptr_deref_1442_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1458_load_1_req_0,
        ptr_deref_1458_load_1_ack_0,
        ptr_deref_1458_load_1_req_1,
        ptr_deref_1458_load_1_ack_1,
        "ptr_deref_1458_load_1",
        "memory_space_3" ,
        ptr_deref_1458_data_1,
        ptr_deref_1458_word_address_1,
        "ptr_deref_1458_data_1",
        "ptr_deref_1458_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1458_load_3_req_0,
        ptr_deref_1458_load_3_ack_0,
        ptr_deref_1458_load_3_req_1,
        ptr_deref_1458_load_3_ack_1,
        "ptr_deref_1458_load_3",
        "memory_space_3" ,
        ptr_deref_1458_data_3,
        ptr_deref_1458_word_address_3,
        "ptr_deref_1458_data_3",
        "ptr_deref_1458_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1442_load_0_req_0,
        ptr_deref_1442_load_0_ack_0,
        ptr_deref_1442_load_0_req_1,
        ptr_deref_1442_load_0_ack_1,
        "ptr_deref_1442_load_0",
        "memory_space_3" ,
        ptr_deref_1442_data_0,
        ptr_deref_1442_word_address_0,
        "ptr_deref_1442_data_0",
        "ptr_deref_1442_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1442_load_2_req_0,
        ptr_deref_1442_load_2_ack_0,
        ptr_deref_1442_load_2_req_1,
        ptr_deref_1442_load_2_ack_1,
        "ptr_deref_1442_load_2",
        "memory_space_3" ,
        ptr_deref_1442_data_2,
        ptr_deref_1442_word_address_2,
        "ptr_deref_1442_data_2",
        "ptr_deref_1442_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1458_load_2_req_0,
        ptr_deref_1458_load_2_ack_0,
        ptr_deref_1458_load_2_req_1,
        ptr_deref_1458_load_2_ack_1,
        "ptr_deref_1458_load_2",
        "memory_space_3" ,
        ptr_deref_1458_data_2,
        ptr_deref_1458_word_address_2,
        "ptr_deref_1458_data_2",
        "ptr_deref_1458_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1407_load_2_req_0,
        ptr_deref_1407_load_2_ack_0,
        ptr_deref_1407_load_2_req_1,
        ptr_deref_1407_load_2_ack_1,
        "ptr_deref_1407_load_2",
        "memory_space_3" ,
        ptr_deref_1407_data_2,
        ptr_deref_1407_word_address_2,
        "ptr_deref_1407_data_2",
        "ptr_deref_1407_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1442_load_1_req_0,
        ptr_deref_1442_load_1_ack_0,
        ptr_deref_1442_load_1_req_1,
        ptr_deref_1442_load_1_ack_1,
        "ptr_deref_1442_load_1",
        "memory_space_3" ,
        ptr_deref_1442_data_1,
        ptr_deref_1442_word_address_1,
        "ptr_deref_1442_data_1",
        "ptr_deref_1442_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1407_load_3_req_0,
        ptr_deref_1407_load_3_ack_0,
        ptr_deref_1407_load_3_req_1,
        ptr_deref_1407_load_3_ack_1,
        "ptr_deref_1407_load_3",
        "memory_space_3" ,
        ptr_deref_1407_data_3,
        ptr_deref_1407_word_address_3,
        "ptr_deref_1407_data_3",
        "ptr_deref_1407_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1407_load_1_req_0,
        ptr_deref_1407_load_1_ack_0,
        ptr_deref_1407_load_1_req_1,
        ptr_deref_1407_load_1_ack_1,
        "ptr_deref_1407_load_1",
        "memory_space_3" ,
        ptr_deref_1407_data_1,
        ptr_deref_1407_word_address_1,
        "ptr_deref_1407_data_1",
        "ptr_deref_1407_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1438_load_3_req_0,
        ptr_deref_1438_load_3_ack_0,
        ptr_deref_1438_load_3_req_1,
        ptr_deref_1438_load_3_ack_1,
        "ptr_deref_1438_load_3",
        "memory_space_3" ,
        ptr_deref_1438_data_3,
        ptr_deref_1438_word_address_3,
        "ptr_deref_1438_data_3",
        "ptr_deref_1438_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1438_load_2_req_0,
        ptr_deref_1438_load_2_ack_0,
        ptr_deref_1438_load_2_req_1,
        ptr_deref_1438_load_2_ack_1,
        "ptr_deref_1438_load_2",
        "memory_space_3" ,
        ptr_deref_1438_data_2,
        ptr_deref_1438_word_address_2,
        "ptr_deref_1438_data_2",
        "ptr_deref_1438_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1438_load_1_req_0,
        ptr_deref_1438_load_1_ack_0,
        ptr_deref_1438_load_1_req_1,
        ptr_deref_1438_load_1_ack_1,
        "ptr_deref_1438_load_1",
        "memory_space_3" ,
        ptr_deref_1438_data_1,
        ptr_deref_1438_word_address_1,
        "ptr_deref_1438_data_1",
        "ptr_deref_1438_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1438_load_0_req_0,
        ptr_deref_1438_load_0_ack_0,
        ptr_deref_1438_load_0_req_1,
        ptr_deref_1438_load_0_ack_1,
        "ptr_deref_1438_load_0",
        "memory_space_3" ,
        ptr_deref_1438_data_0,
        ptr_deref_1438_word_address_0,
        "ptr_deref_1438_data_0",
        "ptr_deref_1438_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1421_load_3_req_0,
        ptr_deref_1421_load_3_ack_0,
        ptr_deref_1421_load_3_req_1,
        ptr_deref_1421_load_3_ack_1,
        "ptr_deref_1421_load_3",
        "memory_space_3" ,
        ptr_deref_1421_data_3,
        ptr_deref_1421_word_address_3,
        "ptr_deref_1421_data_3",
        "ptr_deref_1421_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1421_load_2_req_0,
        ptr_deref_1421_load_2_ack_0,
        ptr_deref_1421_load_2_req_1,
        ptr_deref_1421_load_2_ack_1,
        "ptr_deref_1421_load_2",
        "memory_space_3" ,
        ptr_deref_1421_data_2,
        ptr_deref_1421_word_address_2,
        "ptr_deref_1421_data_2",
        "ptr_deref_1421_word_address_2" -- 
      );
      reqL(20) <= ptr_deref_1421_load_1_req_0;
      reqL(19) <= ptr_deref_1458_load_0_req_0;
      reqL(18) <= ptr_deref_1265_load_0_req_0;
      reqL(17) <= ptr_deref_1421_load_0_req_0;
      reqL(16) <= ptr_deref_1407_load_0_req_0;
      reqL(15) <= ptr_deref_1442_load_3_req_0;
      reqL(14) <= ptr_deref_1458_load_1_req_0;
      reqL(13) <= ptr_deref_1458_load_3_req_0;
      reqL(12) <= ptr_deref_1442_load_0_req_0;
      reqL(11) <= ptr_deref_1442_load_2_req_0;
      reqL(10) <= ptr_deref_1458_load_2_req_0;
      reqL(9) <= ptr_deref_1407_load_2_req_0;
      reqL(8) <= ptr_deref_1442_load_1_req_0;
      reqL(7) <= ptr_deref_1407_load_3_req_0;
      reqL(6) <= ptr_deref_1407_load_1_req_0;
      reqL(5) <= ptr_deref_1438_load_3_req_0;
      reqL(4) <= ptr_deref_1438_load_2_req_0;
      reqL(3) <= ptr_deref_1438_load_1_req_0;
      reqL(2) <= ptr_deref_1438_load_0_req_0;
      reqL(1) <= ptr_deref_1421_load_3_req_0;
      reqL(0) <= ptr_deref_1421_load_2_req_0;
      ptr_deref_1421_load_1_ack_0 <= ackL(20);
      ptr_deref_1458_load_0_ack_0 <= ackL(19);
      ptr_deref_1265_load_0_ack_0 <= ackL(18);
      ptr_deref_1421_load_0_ack_0 <= ackL(17);
      ptr_deref_1407_load_0_ack_0 <= ackL(16);
      ptr_deref_1442_load_3_ack_0 <= ackL(15);
      ptr_deref_1458_load_1_ack_0 <= ackL(14);
      ptr_deref_1458_load_3_ack_0 <= ackL(13);
      ptr_deref_1442_load_0_ack_0 <= ackL(12);
      ptr_deref_1442_load_2_ack_0 <= ackL(11);
      ptr_deref_1458_load_2_ack_0 <= ackL(10);
      ptr_deref_1407_load_2_ack_0 <= ackL(9);
      ptr_deref_1442_load_1_ack_0 <= ackL(8);
      ptr_deref_1407_load_3_ack_0 <= ackL(7);
      ptr_deref_1407_load_1_ack_0 <= ackL(6);
      ptr_deref_1438_load_3_ack_0 <= ackL(5);
      ptr_deref_1438_load_2_ack_0 <= ackL(4);
      ptr_deref_1438_load_1_ack_0 <= ackL(3);
      ptr_deref_1438_load_0_ack_0 <= ackL(2);
      ptr_deref_1421_load_3_ack_0 <= ackL(1);
      ptr_deref_1421_load_2_ack_0 <= ackL(0);
      reqR(20) <= ptr_deref_1421_load_1_req_1;
      reqR(19) <= ptr_deref_1458_load_0_req_1;
      reqR(18) <= ptr_deref_1265_load_0_req_1;
      reqR(17) <= ptr_deref_1421_load_0_req_1;
      reqR(16) <= ptr_deref_1407_load_0_req_1;
      reqR(15) <= ptr_deref_1442_load_3_req_1;
      reqR(14) <= ptr_deref_1458_load_1_req_1;
      reqR(13) <= ptr_deref_1458_load_3_req_1;
      reqR(12) <= ptr_deref_1442_load_0_req_1;
      reqR(11) <= ptr_deref_1442_load_2_req_1;
      reqR(10) <= ptr_deref_1458_load_2_req_1;
      reqR(9) <= ptr_deref_1407_load_2_req_1;
      reqR(8) <= ptr_deref_1442_load_1_req_1;
      reqR(7) <= ptr_deref_1407_load_3_req_1;
      reqR(6) <= ptr_deref_1407_load_1_req_1;
      reqR(5) <= ptr_deref_1438_load_3_req_1;
      reqR(4) <= ptr_deref_1438_load_2_req_1;
      reqR(3) <= ptr_deref_1438_load_1_req_1;
      reqR(2) <= ptr_deref_1438_load_0_req_1;
      reqR(1) <= ptr_deref_1421_load_3_req_1;
      reqR(0) <= ptr_deref_1421_load_2_req_1;
      ptr_deref_1421_load_1_ack_1 <= ackR(20);
      ptr_deref_1458_load_0_ack_1 <= ackR(19);
      ptr_deref_1265_load_0_ack_1 <= ackR(18);
      ptr_deref_1421_load_0_ack_1 <= ackR(17);
      ptr_deref_1407_load_0_ack_1 <= ackR(16);
      ptr_deref_1442_load_3_ack_1 <= ackR(15);
      ptr_deref_1458_load_1_ack_1 <= ackR(14);
      ptr_deref_1458_load_3_ack_1 <= ackR(13);
      ptr_deref_1442_load_0_ack_1 <= ackR(12);
      ptr_deref_1442_load_2_ack_1 <= ackR(11);
      ptr_deref_1458_load_2_ack_1 <= ackR(10);
      ptr_deref_1407_load_2_ack_1 <= ackR(9);
      ptr_deref_1442_load_1_ack_1 <= ackR(8);
      ptr_deref_1407_load_3_ack_1 <= ackR(7);
      ptr_deref_1407_load_1_ack_1 <= ackR(6);
      ptr_deref_1438_load_3_ack_1 <= ackR(5);
      ptr_deref_1438_load_2_ack_1 <= ackR(4);
      ptr_deref_1438_load_1_ack_1 <= ackR(3);
      ptr_deref_1438_load_0_ack_1 <= ackR(2);
      ptr_deref_1421_load_3_ack_1 <= ackR(1);
      ptr_deref_1421_load_2_ack_1 <= ackR(0);
      data_in <= ptr_deref_1421_word_address_1 & ptr_deref_1458_word_address_0 & ptr_deref_1265_word_address_0 & ptr_deref_1421_word_address_0 & ptr_deref_1407_word_address_0 & ptr_deref_1442_word_address_3 & ptr_deref_1458_word_address_1 & ptr_deref_1458_word_address_3 & ptr_deref_1442_word_address_0 & ptr_deref_1442_word_address_2 & ptr_deref_1458_word_address_2 & ptr_deref_1407_word_address_2 & ptr_deref_1442_word_address_1 & ptr_deref_1407_word_address_3 & ptr_deref_1407_word_address_1 & ptr_deref_1438_word_address_3 & ptr_deref_1438_word_address_2 & ptr_deref_1438_word_address_1 & ptr_deref_1438_word_address_0 & ptr_deref_1421_word_address_3 & ptr_deref_1421_word_address_2;
      ptr_deref_1421_data_1 <= data_out(167 downto 160);
      ptr_deref_1458_data_0 <= data_out(159 downto 152);
      ptr_deref_1265_data_0 <= data_out(151 downto 144);
      ptr_deref_1421_data_0 <= data_out(143 downto 136);
      ptr_deref_1407_data_0 <= data_out(135 downto 128);
      ptr_deref_1442_data_3 <= data_out(127 downto 120);
      ptr_deref_1458_data_1 <= data_out(119 downto 112);
      ptr_deref_1458_data_3 <= data_out(111 downto 104);
      ptr_deref_1442_data_0 <= data_out(103 downto 96);
      ptr_deref_1442_data_2 <= data_out(95 downto 88);
      ptr_deref_1458_data_2 <= data_out(87 downto 80);
      ptr_deref_1407_data_2 <= data_out(79 downto 72);
      ptr_deref_1442_data_1 <= data_out(71 downto 64);
      ptr_deref_1407_data_3 <= data_out(63 downto 56);
      ptr_deref_1407_data_1 <= data_out(55 downto 48);
      ptr_deref_1438_data_3 <= data_out(47 downto 40);
      ptr_deref_1438_data_2 <= data_out(39 downto 32);
      ptr_deref_1438_data_1 <= data_out(31 downto 24);
      ptr_deref_1438_data_0 <= data_out(23 downto 16);
      ptr_deref_1421_data_3 <= data_out(15 downto 8);
      ptr_deref_1421_data_2 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 14,
        num_reqs => 21,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 21,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1565_load_0 ptr_deref_1501_load_0 ptr_deref_1533_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(26 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1565_load_0_req_0,
        ptr_deref_1565_load_0_ack_0,
        ptr_deref_1565_load_0_req_1,
        ptr_deref_1565_load_0_ack_1,
        "ptr_deref_1565_load_0",
        "memory_space_1" ,
        ptr_deref_1565_data_0,
        ptr_deref_1565_word_address_0,
        "ptr_deref_1565_data_0",
        "ptr_deref_1565_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1501_load_0_req_0,
        ptr_deref_1501_load_0_ack_0,
        ptr_deref_1501_load_0_req_1,
        ptr_deref_1501_load_0_ack_1,
        "ptr_deref_1501_load_0",
        "memory_space_1" ,
        ptr_deref_1501_data_0,
        ptr_deref_1501_word_address_0,
        "ptr_deref_1501_data_0",
        "ptr_deref_1501_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1533_load_0_req_0,
        ptr_deref_1533_load_0_ack_0,
        ptr_deref_1533_load_0_req_1,
        ptr_deref_1533_load_0_ack_1,
        "ptr_deref_1533_load_0",
        "memory_space_1" ,
        ptr_deref_1533_data_0,
        ptr_deref_1533_word_address_0,
        "ptr_deref_1533_data_0",
        "ptr_deref_1533_word_address_0" -- 
      );
      reqL(2) <= ptr_deref_1565_load_0_req_0;
      reqL(1) <= ptr_deref_1501_load_0_req_0;
      reqL(0) <= ptr_deref_1533_load_0_req_0;
      ptr_deref_1565_load_0_ack_0 <= ackL(2);
      ptr_deref_1501_load_0_ack_0 <= ackL(1);
      ptr_deref_1533_load_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1565_load_0_req_1;
      reqR(1) <= ptr_deref_1501_load_0_req_1;
      reqR(0) <= ptr_deref_1533_load_0_req_1;
      ptr_deref_1565_load_0_ack_1 <= ackR(2);
      ptr_deref_1501_load_0_ack_1 <= ackR(1);
      ptr_deref_1533_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1565_word_address_0 & ptr_deref_1501_word_address_0 & ptr_deref_1533_word_address_0;
      ptr_deref_1565_data_0 <= data_out(23 downto 16);
      ptr_deref_1501_data_0 <= data_out(15 downto 8);
      ptr_deref_1533_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 9,
        num_reqs => 3,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(8 downto 0),
          mtag => memory_space_1_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : simple_obj_ref_1213_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        simple_obj_ref_1213_load_0_req_0,
        simple_obj_ref_1213_load_0_ack_0,
        simple_obj_ref_1213_load_0_req_1,
        simple_obj_ref_1213_load_0_ack_1,
        "simple_obj_ref_1213_load_0",
        "memory_space_4" ,
        simple_obj_ref_1213_data_0,
        simple_obj_ref_1213_word_address_0,
        "simple_obj_ref_1213_data_0",
        "simple_obj_ref_1213_word_address_0" -- 
      );
      reqL(0) <= simple_obj_ref_1213_load_0_req_0;
      simple_obj_ref_1213_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1213_load_0_req_1;
      simple_obj_ref_1213_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_1213_word_address_0;
      simple_obj_ref_1213_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_1350_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1350_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1350_word_address_0) &  " data ptr_deref_1350_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1350_data_0) severity note; --
        end if;
        if ptr_deref_1336_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1336_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1336_word_address_0) &  " data ptr_deref_1336_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1336_data_0) severity note; --
        end if;
        if ptr_deref_1416_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1416_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1416_word_address_3) &  " data ptr_deref_1416_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1416_data_3) severity note; --
        end if;
        if ptr_deref_1463_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1463_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1463_word_address_0) &  " data ptr_deref_1463_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1463_data_0) severity note; --
        end if;
        if ptr_deref_1416_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1416_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1416_word_address_2) &  " data ptr_deref_1416_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1416_data_2) severity note; --
        end if;
        if ptr_deref_1368_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1368_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1368_word_address_1) &  " data ptr_deref_1368_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1368_data_1) severity note; --
        end if;
        if ptr_deref_1368_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1368_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1368_word_address_2) &  " data ptr_deref_1368_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1368_data_2) severity note; --
        end if;
        if ptr_deref_1368_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1368_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1368_word_address_3) &  " data ptr_deref_1368_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1368_data_3) severity note; --
        end if;
        if ptr_deref_1416_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1416_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1416_word_address_0) &  " data ptr_deref_1416_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1416_data_0) severity note; --
        end if;
        if ptr_deref_1399_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1399_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1399_word_address_0) &  " data ptr_deref_1399_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1399_data_0) severity note; --
        end if;
        if ptr_deref_1416_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1416_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1416_word_address_1) &  " data ptr_deref_1416_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1416_data_1) severity note; --
        end if;
        if ptr_deref_1368_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1368_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1368_word_address_0) &  " data ptr_deref_1368_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1368_data_0) severity note; --
        end if;
        if ptr_deref_1350_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1350_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1350_word_address_1) &  " data ptr_deref_1350_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1350_data_1) severity note; --
        end if;
        if ptr_deref_1350_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1350_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1350_word_address_2) &  " data ptr_deref_1350_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1350_data_2) severity note; --
        end if;
        if ptr_deref_1350_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1350_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1350_word_address_3) &  " data ptr_deref_1350_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1350_data_3) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1350_store_0 ptr_deref_1336_store_0 ptr_deref_1416_store_3 ptr_deref_1463_store_0 ptr_deref_1416_store_2 ptr_deref_1368_store_1 ptr_deref_1368_store_2 ptr_deref_1368_store_3 ptr_deref_1416_store_0 ptr_deref_1399_store_0 ptr_deref_1416_store_1 ptr_deref_1368_store_0 ptr_deref_1350_store_1 ptr_deref_1350_store_2 ptr_deref_1350_store_3 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(209 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= ptr_deref_1350_store_0_req_0;
      reqL(13) <= ptr_deref_1336_store_0_req_0;
      reqL(12) <= ptr_deref_1416_store_3_req_0;
      reqL(11) <= ptr_deref_1463_store_0_req_0;
      reqL(10) <= ptr_deref_1416_store_2_req_0;
      reqL(9) <= ptr_deref_1368_store_1_req_0;
      reqL(8) <= ptr_deref_1368_store_2_req_0;
      reqL(7) <= ptr_deref_1368_store_3_req_0;
      reqL(6) <= ptr_deref_1416_store_0_req_0;
      reqL(5) <= ptr_deref_1399_store_0_req_0;
      reqL(4) <= ptr_deref_1416_store_1_req_0;
      reqL(3) <= ptr_deref_1368_store_0_req_0;
      reqL(2) <= ptr_deref_1350_store_1_req_0;
      reqL(1) <= ptr_deref_1350_store_2_req_0;
      reqL(0) <= ptr_deref_1350_store_3_req_0;
      ptr_deref_1350_store_0_ack_0 <= ackL(14);
      ptr_deref_1336_store_0_ack_0 <= ackL(13);
      ptr_deref_1416_store_3_ack_0 <= ackL(12);
      ptr_deref_1463_store_0_ack_0 <= ackL(11);
      ptr_deref_1416_store_2_ack_0 <= ackL(10);
      ptr_deref_1368_store_1_ack_0 <= ackL(9);
      ptr_deref_1368_store_2_ack_0 <= ackL(8);
      ptr_deref_1368_store_3_ack_0 <= ackL(7);
      ptr_deref_1416_store_0_ack_0 <= ackL(6);
      ptr_deref_1399_store_0_ack_0 <= ackL(5);
      ptr_deref_1416_store_1_ack_0 <= ackL(4);
      ptr_deref_1368_store_0_ack_0 <= ackL(3);
      ptr_deref_1350_store_1_ack_0 <= ackL(2);
      ptr_deref_1350_store_2_ack_0 <= ackL(1);
      ptr_deref_1350_store_3_ack_0 <= ackL(0);
      reqR(14) <= ptr_deref_1350_store_0_req_1;
      reqR(13) <= ptr_deref_1336_store_0_req_1;
      reqR(12) <= ptr_deref_1416_store_3_req_1;
      reqR(11) <= ptr_deref_1463_store_0_req_1;
      reqR(10) <= ptr_deref_1416_store_2_req_1;
      reqR(9) <= ptr_deref_1368_store_1_req_1;
      reqR(8) <= ptr_deref_1368_store_2_req_1;
      reqR(7) <= ptr_deref_1368_store_3_req_1;
      reqR(6) <= ptr_deref_1416_store_0_req_1;
      reqR(5) <= ptr_deref_1399_store_0_req_1;
      reqR(4) <= ptr_deref_1416_store_1_req_1;
      reqR(3) <= ptr_deref_1368_store_0_req_1;
      reqR(2) <= ptr_deref_1350_store_1_req_1;
      reqR(1) <= ptr_deref_1350_store_2_req_1;
      reqR(0) <= ptr_deref_1350_store_3_req_1;
      ptr_deref_1350_store_0_ack_1 <= ackR(14);
      ptr_deref_1336_store_0_ack_1 <= ackR(13);
      ptr_deref_1416_store_3_ack_1 <= ackR(12);
      ptr_deref_1463_store_0_ack_1 <= ackR(11);
      ptr_deref_1416_store_2_ack_1 <= ackR(10);
      ptr_deref_1368_store_1_ack_1 <= ackR(9);
      ptr_deref_1368_store_2_ack_1 <= ackR(8);
      ptr_deref_1368_store_3_ack_1 <= ackR(7);
      ptr_deref_1416_store_0_ack_1 <= ackR(6);
      ptr_deref_1399_store_0_ack_1 <= ackR(5);
      ptr_deref_1416_store_1_ack_1 <= ackR(4);
      ptr_deref_1368_store_0_ack_1 <= ackR(3);
      ptr_deref_1350_store_1_ack_1 <= ackR(2);
      ptr_deref_1350_store_2_ack_1 <= ackR(1);
      ptr_deref_1350_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1350_word_address_0 & ptr_deref_1336_word_address_0 & ptr_deref_1416_word_address_3 & ptr_deref_1463_word_address_0 & ptr_deref_1416_word_address_2 & ptr_deref_1368_word_address_1 & ptr_deref_1368_word_address_2 & ptr_deref_1368_word_address_3 & ptr_deref_1416_word_address_0 & ptr_deref_1399_word_address_0 & ptr_deref_1416_word_address_1 & ptr_deref_1368_word_address_0 & ptr_deref_1350_word_address_1 & ptr_deref_1350_word_address_2 & ptr_deref_1350_word_address_3;
      data_in <= ptr_deref_1350_data_0 & ptr_deref_1336_data_0 & ptr_deref_1416_data_3 & ptr_deref_1463_data_0 & ptr_deref_1416_data_2 & ptr_deref_1368_data_1 & ptr_deref_1368_data_2 & ptr_deref_1368_data_3 & ptr_deref_1416_data_0 & ptr_deref_1399_data_0 & ptr_deref_1416_data_1 & ptr_deref_1368_data_0 & ptr_deref_1350_data_1 & ptr_deref_1350_data_2 & ptr_deref_1350_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 14,
        data_width => 8,
        num_reqs => 15,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1221_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_4 address simple_obj_ref_1221_word_address_0 ="  &  convert_slv_to_hex_string(simple_obj_ref_1221_word_address_0) &  " data simple_obj_ref_1221_data_0 ="  &  convert_slv_to_hex_string(simple_obj_ref_1221_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (1) : simple_obj_ref_1221_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1221_store_0_req_0;
      simple_obj_ref_1221_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1221_store_0_req_1;
      simple_obj_ref_1221_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_1221_word_address_0;
      data_in <= simple_obj_ref_1221_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : simple_obj_ref_1093_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_1093_inst_ack_0 then -- 
            assert false report " ReadPipe rtt_in0 to wire simple_obj_ref_1093_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_1093_inst_req_0;
      simple_obj_ref_1093_inst_ack_0 <= ack(0);
      simple_obj_ref_1093_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => rtt_in0_pipe_read_req(0),
          oack => rtt_in0_pipe_read_ack(0),
          odata => rtt_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1665_inst_ack_0 then -- 
          assert false report " WritePipe to0_in0 from wire type_cast_1667_wire value="  &  convert_slv_to_hex_string(type_cast_1667_wire) severity note; --
        end if;
        if simple_obj_ref_1689_inst_ack_0 then -- 
          assert false report " WritePipe to0_in0 from wire type_cast_1691_wire value="  &  convert_slv_to_hex_string(type_cast_1691_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_1665_inst simple_obj_ref_1689_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_1665_inst_req_0;
      req(0) <= simple_obj_ref_1689_inst_req_0;
      simple_obj_ref_1665_inst_ack_0 <= ack(1);
      simple_obj_ref_1689_inst_ack_0 <= ack(0);
      data_in <= type_cast_1667_wire & type_cast_1691_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to0_in0_pipe_write_req(0),
          oack => to0_in0_pipe_write_ack(0),
          odata => to0_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1671_inst_ack_0 then -- 
          assert false report " WritePipe to1_in0 from wire type_cast_1673_wire value="  &  convert_slv_to_hex_string(type_cast_1673_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_1671_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1671_inst_req_0;
      simple_obj_ref_1671_inst_ack_0 <= ack(0);
      data_in <= type_cast_1673_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to1_in0_pipe_write_req(0),
          oack => to1_in0_pipe_write_ack(0),
          odata => to1_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1677_inst_ack_0 then -- 
          assert false report " WritePipe to2_in0 from wire type_cast_1679_wire value="  &  convert_slv_to_hex_string(type_cast_1679_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (2) : simple_obj_ref_1677_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1677_inst_req_0;
      simple_obj_ref_1677_inst_ack_0 <= ack(0);
      data_in <= type_cast_1679_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to2_in0_pipe_write_req(0),
          oack => to2_in0_pipe_write_ack(0),
          odata => to2_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1683_inst_ack_0 then -- 
          assert false report " WritePipe to3_in0 from wire type_cast_1685_wire value="  &  convert_slv_to_hex_string(type_cast_1685_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (3) : simple_obj_ref_1683_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1683_inst_req_0;
      simple_obj_ref_1683_inst_ack_0 <= ack(0);
      data_in <= type_cast_1685_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to3_in0_pipe_write_req(0),
          oack => to3_in0_pipe_write_ack(0),
          odata => to3_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1470_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1470_call_req_0;
      call_stmt_1470_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1470_call_req_1;
      call_stmt_1470_call_ack_1 <= ackR(0);
      data_in <= tmp_1095;
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 32,
        owidth => 32,
        twidth => 3,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_packet_free_call_reqs(0),
          ackR => ahir_packet_free_call_acks(0),
          dataR => ahir_packet_free_call_data(31 downto 0),
          tagR => ahir_packet_free_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 3, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => ahir_packet_free_return_acks(0), -- cross-over
          ackL => ahir_packet_free_return_reqs(0), -- cross-over
          tagL => ahir_packet_free_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_src is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    src_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    src_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    src_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    chk_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    chk_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    chk_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_src;
architecture Default of ahir_glue_src is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_src_CP_7782_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_1756_root_address_inst_req_1 : boolean;
  signal ptr_deref_1759_addr_3_ack_0 : boolean;
  signal ptr_deref_1759_addr_3_req_1 : boolean;
  signal array_obj_ref_1756_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1759_base_resize_req_0 : boolean;
  signal ptr_deref_1759_addr_2_req_1 : boolean;
  signal array_obj_ref_1756_final_reg_ack_0 : boolean;
  signal ptr_deref_1759_store_3_ack_1 : boolean;
  signal ptr_deref_1759_store_2_req_0 : boolean;
  signal ptr_deref_1759_store_3_ack_0 : boolean;
  signal type_cast_1770_inst_ack_0 : boolean;
  signal ptr_deref_1759_addr_1_ack_1 : boolean;
  signal ptr_deref_1759_addr_0_req_0 : boolean;
  signal ptr_deref_1759_addr_0_ack_0 : boolean;
  signal ptr_deref_1759_addr_3_req_0 : boolean;
  signal binary_1745_inst_req_0 : boolean;
  signal array_obj_ref_1756_final_reg_req_0 : boolean;
  signal binary_1766_inst_ack_1 : boolean;
  signal ptr_deref_1759_addr_0_req_1 : boolean;
  signal ptr_deref_1774_addr_1_ack_1 : boolean;
  signal ptr_deref_1759_store_2_req_1 : boolean;
  signal ptr_deref_1759_base_resize_ack_0 : boolean;
  signal ptr_deref_1759_addr_2_ack_1 : boolean;
  signal ptr_deref_1759_store_1_ack_1 : boolean;
  signal ptr_deref_1759_addr_3_ack_1 : boolean;
  signal ptr_deref_1759_store_0_ack_0 : boolean;
  signal array_obj_ref_1756_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1759_store_3_req_0 : boolean;
  signal ptr_deref_1774_addr_0_ack_1 : boolean;
  signal ptr_deref_1774_load_1_ack_0 : boolean;
  signal ptr_deref_1774_root_address_inst_req_0 : boolean;
  signal ptr_deref_1774_addr_1_ack_0 : boolean;
  signal ptr_deref_1759_addr_2_ack_0 : boolean;
  signal binary_1745_inst_ack_1 : boolean;
  signal ptr_deref_1774_load_0_req_0 : boolean;
  signal ptr_deref_1774_gather_scatter_req_0 : boolean;
  signal ptr_deref_1759_addr_2_req_0 : boolean;
  signal ptr_deref_1759_store_0_req_0 : boolean;
  signal call_stmt_1778_call_req_1 : boolean;
  signal ptr_deref_1759_store_0_req_1 : boolean;
  signal ptr_deref_1774_base_resize_ack_0 : boolean;
  signal type_cast_1749_inst_req_0 : boolean;
  signal array_obj_ref_1756_root_address_inst_req_0 : boolean;
  signal call_stmt_1778_call_ack_1 : boolean;
  signal ptr_deref_1759_store_2_ack_1 : boolean;
  signal type_cast_1749_inst_ack_0 : boolean;
  signal binary_1745_inst_req_1 : boolean;
  signal binary_1745_inst_ack_0 : boolean;
  signal ptr_deref_1774_addr_0_ack_0 : boolean;
  signal ptr_deref_1759_store_0_ack_1 : boolean;
  signal ptr_deref_1759_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1759_addr_1_req_0 : boolean;
  signal ptr_deref_1774_addr_0_req_1 : boolean;
  signal ptr_deref_1774_addr_0_req_0 : boolean;
  signal ptr_deref_1774_addr_1_req_1 : boolean;
  signal ptr_deref_1759_store_1_req_1 : boolean;
  signal ptr_deref_1759_addr_0_ack_1 : boolean;
  signal ptr_deref_1759_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1785_offset_inst_req_0 : boolean;
  signal array_obj_ref_1785_offset_inst_ack_0 : boolean;
  signal call_stmt_1778_call_req_0 : boolean;
  signal ptr_deref_1774_load_1_req_0 : boolean;
  signal ptr_deref_1759_store_3_req_1 : boolean;
  signal ptr_deref_1774_load_0_req_1 : boolean;
  signal array_obj_ref_1785_final_reg_ack_0 : boolean;
  signal ptr_deref_1759_addr_1_ack_0 : boolean;
  signal ptr_deref_1774_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1785_base_resize_req_0 : boolean;
  signal array_obj_ref_1785_base_resize_ack_0 : boolean;
  signal ptr_deref_1774_load_1_req_1 : boolean;
  signal ptr_deref_1759_store_1_req_0 : boolean;
  signal array_obj_ref_1785_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1785_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1774_load_0_ack_1 : boolean;
  signal binary_1766_inst_ack_0 : boolean;
  signal ptr_deref_1774_load_1_ack_1 : boolean;
  signal ptr_deref_1774_base_resize_req_0 : boolean;
  signal ptr_deref_1774_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1759_store_1_ack_0 : boolean;
  signal array_obj_ref_1785_root_address_inst_req_0 : boolean;
  signal binary_1766_inst_req_1 : boolean;
  signal ptr_deref_1774_load_0_ack_0 : boolean;
  signal ptr_deref_1774_addr_1_req_0 : boolean;
  signal type_cast_1770_inst_req_0 : boolean;
  signal ptr_deref_1759_gather_scatter_req_0 : boolean;
  signal type_cast_1781_inst_ack_0 : boolean;
  signal array_obj_ref_1756_base_resize_req_0 : boolean;
  signal ptr_deref_1759_store_2_ack_0 : boolean;
  signal type_cast_1781_inst_req_0 : boolean;
  signal ptr_deref_1759_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1792_base_resize_req_0 : boolean;
  signal array_obj_ref_1792_base_resize_ack_0 : boolean;
  signal array_obj_ref_1785_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1785_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1785_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1785_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1785_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1785_final_reg_req_0 : boolean;
  signal call_stmt_1778_call_ack_0 : boolean;
  signal ptr_deref_1759_addr_1_req_1 : boolean;
  signal binary_1766_inst_req_0 : boolean;
  signal array_obj_ref_1756_base_resize_ack_0 : boolean;
  signal simple_obj_ref_1702_inst_req_0 : boolean;
  signal simple_obj_ref_1702_inst_ack_0 : boolean;
  signal type_cast_1703_inst_req_0 : boolean;
  signal type_cast_1703_inst_ack_0 : boolean;
  signal binary_1709_inst_req_0 : boolean;
  signal binary_1709_inst_ack_0 : boolean;
  signal binary_1709_inst_req_1 : boolean;
  signal binary_1709_inst_ack_1 : boolean;
  signal binary_1715_inst_req_0 : boolean;
  signal binary_1715_inst_ack_0 : boolean;
  signal binary_1715_inst_req_1 : boolean;
  signal binary_1715_inst_ack_1 : boolean;
  signal type_cast_1719_inst_req_0 : boolean;
  signal type_cast_1719_inst_ack_0 : boolean;
  signal type_cast_1723_inst_req_0 : boolean;
  signal type_cast_1723_inst_ack_0 : boolean;
  signal array_obj_ref_1728_base_resize_req_0 : boolean;
  signal array_obj_ref_1728_base_resize_ack_0 : boolean;
  signal array_obj_ref_1728_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1728_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1728_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1728_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1728_final_reg_req_0 : boolean;
  signal array_obj_ref_1728_final_reg_ack_0 : boolean;
  signal array_obj_ref_1735_base_resize_req_0 : boolean;
  signal array_obj_ref_1735_base_resize_ack_0 : boolean;
  signal array_obj_ref_1735_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1735_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1735_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1735_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1735_final_reg_req_0 : boolean;
  signal array_obj_ref_1735_final_reg_ack_0 : boolean;
  signal ptr_deref_1738_base_resize_req_0 : boolean;
  signal ptr_deref_1738_base_resize_ack_0 : boolean;
  signal ptr_deref_1738_root_address_inst_req_0 : boolean;
  signal ptr_deref_1738_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1738_addr_0_req_0 : boolean;
  signal ptr_deref_1738_addr_0_ack_0 : boolean;
  signal ptr_deref_1738_addr_0_req_1 : boolean;
  signal ptr_deref_1738_addr_0_ack_1 : boolean;
  signal ptr_deref_1738_addr_1_req_0 : boolean;
  signal ptr_deref_1738_addr_1_ack_0 : boolean;
  signal ptr_deref_1738_addr_1_req_1 : boolean;
  signal ptr_deref_1738_addr_1_ack_1 : boolean;
  signal ptr_deref_1738_addr_2_req_0 : boolean;
  signal ptr_deref_1738_addr_2_ack_0 : boolean;
  signal ptr_deref_1738_addr_2_req_1 : boolean;
  signal ptr_deref_1738_addr_2_ack_1 : boolean;
  signal ptr_deref_1738_addr_3_req_0 : boolean;
  signal ptr_deref_1738_addr_3_ack_0 : boolean;
  signal ptr_deref_1738_addr_3_req_1 : boolean;
  signal ptr_deref_1738_addr_3_ack_1 : boolean;
  signal ptr_deref_1738_gather_scatter_req_0 : boolean;
  signal ptr_deref_1738_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1738_store_0_req_0 : boolean;
  signal ptr_deref_1738_store_0_ack_0 : boolean;
  signal ptr_deref_1738_store_1_req_0 : boolean;
  signal ptr_deref_1738_store_1_ack_0 : boolean;
  signal ptr_deref_1738_store_2_req_0 : boolean;
  signal ptr_deref_1738_store_2_ack_0 : boolean;
  signal ptr_deref_1738_store_3_req_0 : boolean;
  signal ptr_deref_1738_store_3_ack_0 : boolean;
  signal ptr_deref_1738_store_0_req_1 : boolean;
  signal ptr_deref_1738_store_0_ack_1 : boolean;
  signal ptr_deref_1738_store_1_req_1 : boolean;
  signal ptr_deref_1738_store_1_ack_1 : boolean;
  signal ptr_deref_1738_store_2_req_1 : boolean;
  signal ptr_deref_1738_store_2_ack_1 : boolean;
  signal ptr_deref_1738_store_3_req_1 : boolean;
  signal ptr_deref_1738_store_3_ack_1 : boolean;
  signal array_obj_ref_1792_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1792_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1792_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1792_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1792_final_reg_req_0 : boolean;
  signal array_obj_ref_1792_final_reg_ack_0 : boolean;
  signal ptr_deref_1795_base_resize_req_0 : boolean;
  signal ptr_deref_1795_base_resize_ack_0 : boolean;
  signal ptr_deref_1795_root_address_inst_req_0 : boolean;
  signal ptr_deref_1795_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1795_addr_0_req_0 : boolean;
  signal ptr_deref_1795_addr_0_ack_0 : boolean;
  signal ptr_deref_1795_addr_0_req_1 : boolean;
  signal ptr_deref_1795_addr_0_ack_1 : boolean;
  signal ptr_deref_1795_addr_1_req_0 : boolean;
  signal ptr_deref_1795_addr_1_ack_0 : boolean;
  signal ptr_deref_1795_addr_1_req_1 : boolean;
  signal ptr_deref_1795_addr_1_ack_1 : boolean;
  signal ptr_deref_1795_addr_2_req_0 : boolean;
  signal ptr_deref_1795_addr_2_ack_0 : boolean;
  signal ptr_deref_1795_addr_2_req_1 : boolean;
  signal ptr_deref_1795_addr_2_ack_1 : boolean;
  signal ptr_deref_1795_addr_3_req_0 : boolean;
  signal ptr_deref_1795_addr_3_ack_0 : boolean;
  signal ptr_deref_1795_addr_3_req_1 : boolean;
  signal ptr_deref_1795_addr_3_ack_1 : boolean;
  signal ptr_deref_1795_gather_scatter_req_0 : boolean;
  signal ptr_deref_1795_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1795_store_0_req_0 : boolean;
  signal ptr_deref_1795_store_0_ack_0 : boolean;
  signal ptr_deref_1795_store_1_req_0 : boolean;
  signal ptr_deref_1795_store_1_ack_0 : boolean;
  signal ptr_deref_1795_store_2_req_0 : boolean;
  signal ptr_deref_1795_store_2_ack_0 : boolean;
  signal ptr_deref_1795_store_3_req_0 : boolean;
  signal ptr_deref_1795_store_3_ack_0 : boolean;
  signal ptr_deref_1795_store_0_req_1 : boolean;
  signal ptr_deref_1795_store_0_ack_1 : boolean;
  signal ptr_deref_1795_store_1_req_1 : boolean;
  signal ptr_deref_1795_store_1_ack_1 : boolean;
  signal ptr_deref_1795_store_2_req_1 : boolean;
  signal ptr_deref_1795_store_2_ack_1 : boolean;
  signal ptr_deref_1795_store_3_req_1 : boolean;
  signal ptr_deref_1795_store_3_ack_1 : boolean;
  signal binary_1802_inst_req_0 : boolean;
  signal binary_1802_inst_ack_0 : boolean;
  signal binary_1802_inst_req_1 : boolean;
  signal binary_1802_inst_ack_1 : boolean;
  signal binary_1808_inst_req_0 : boolean;
  signal binary_1808_inst_ack_0 : boolean;
  signal binary_1808_inst_req_1 : boolean;
  signal binary_1808_inst_ack_1 : boolean;
  signal type_cast_1812_inst_req_0 : boolean;
  signal type_cast_1812_inst_ack_0 : boolean;
  signal array_obj_ref_1819_base_resize_req_0 : boolean;
  signal array_obj_ref_1819_base_resize_ack_0 : boolean;
  signal array_obj_ref_1819_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1819_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1819_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1819_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1819_final_reg_req_0 : boolean;
  signal array_obj_ref_1819_final_reg_ack_0 : boolean;
  signal ptr_deref_1822_base_resize_req_0 : boolean;
  signal ptr_deref_1822_base_resize_ack_0 : boolean;
  signal ptr_deref_1822_root_address_inst_req_0 : boolean;
  signal ptr_deref_1822_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1822_addr_0_req_0 : boolean;
  signal ptr_deref_1822_addr_0_ack_0 : boolean;
  signal ptr_deref_1822_addr_0_req_1 : boolean;
  signal ptr_deref_1822_addr_0_ack_1 : boolean;
  signal ptr_deref_1822_addr_1_req_0 : boolean;
  signal ptr_deref_1822_addr_1_ack_0 : boolean;
  signal ptr_deref_1822_addr_1_req_1 : boolean;
  signal ptr_deref_1822_addr_1_ack_1 : boolean;
  signal ptr_deref_1822_addr_2_req_0 : boolean;
  signal ptr_deref_1822_addr_2_ack_0 : boolean;
  signal ptr_deref_1822_addr_2_req_1 : boolean;
  signal ptr_deref_1822_addr_2_ack_1 : boolean;
  signal ptr_deref_1822_addr_3_req_0 : boolean;
  signal ptr_deref_1822_addr_3_ack_0 : boolean;
  signal ptr_deref_1822_addr_3_req_1 : boolean;
  signal ptr_deref_1822_addr_3_ack_1 : boolean;
  signal ptr_deref_1822_gather_scatter_req_0 : boolean;
  signal ptr_deref_1822_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1822_store_0_req_0 : boolean;
  signal ptr_deref_1822_store_0_ack_0 : boolean;
  signal ptr_deref_1822_store_1_req_0 : boolean;
  signal ptr_deref_1822_store_1_ack_0 : boolean;
  signal ptr_deref_1822_store_2_req_0 : boolean;
  signal ptr_deref_1822_store_2_ack_0 : boolean;
  signal ptr_deref_1822_store_3_req_0 : boolean;
  signal ptr_deref_1822_store_3_ack_0 : boolean;
  signal ptr_deref_1822_store_0_req_1 : boolean;
  signal ptr_deref_1822_store_0_ack_1 : boolean;
  signal ptr_deref_1822_store_1_req_1 : boolean;
  signal ptr_deref_1822_store_1_ack_1 : boolean;
  signal ptr_deref_1822_store_2_req_1 : boolean;
  signal ptr_deref_1822_store_2_ack_1 : boolean;
  signal ptr_deref_1822_store_3_req_1 : boolean;
  signal ptr_deref_1822_store_3_ack_1 : boolean;
  signal type_cast_1827_inst_req_0 : boolean;
  signal type_cast_1827_inst_ack_0 : boolean;
  signal simple_obj_ref_1825_inst_req_0 : boolean;
  signal simple_obj_ref_1825_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_src_CP_7782: Block -- control-path 
    signal cp_elements: BooleanArray(284 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(284);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(284), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(160);
    crr_8275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_1778_call_req_0); -- 
    cp_elements(2) <= cp_elements(278);
    cp_elements(3) <= cp_elements(0);
    cpelement_group_4 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(5) & cp_elements(7));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(4),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7818_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => type_cast_1703_inst_req_0); -- 
    cp_elements(5) <= cp_elements(3);
    cp_elements(6) <= cp_elements(3);
    req_7813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => simple_obj_ref_1702_inst_req_0); -- 
    ack_7814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1702_inst_ack_0, ack => cp_elements(7)); -- 
    ack_7819_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1703_inst_ack_0, ack => cp_elements(8)); -- 
    cp_elements(9) <= cp_elements(8);
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(12));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => binary_1709_inst_req_0); -- 
    cp_elements(11) <= cp_elements(9);
    cp_elements(12) <= cp_elements(9);
    ra_7832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1709_inst_ack_0, ack => cp_elements(13)); -- 
    cr_7833_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => binary_1709_inst_req_1); -- 
    cp_elements(14) <= binary_1709_inst_ack_1;
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_1715_inst_req_0); -- 
    cp_elements(16) <= cp_elements(9);
    cp_elements(17) <= cp_elements(14);
    ra_7844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1715_inst_ack_0, ack => cp_elements(18)); -- 
    cr_7845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_1715_inst_req_1); -- 
    cp_elements(19) <= binary_1715_inst_ack_1;
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(21) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_1719_inst_req_0); -- 
    cp_elements(21) <= cp_elements(9);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= type_cast_1719_inst_ack_0;
    cpelement_group_24 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(25) & cp_elements(26));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(24),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => type_cast_1723_inst_req_0); -- 
    cp_elements(25) <= cp_elements(9);
    cp_elements(26) <= cp_elements(19);
    ack_7866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_0, ack => cp_elements(27)); -- 
    base_resize_req_7877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => array_obj_ref_1728_base_resize_req_0); -- 
    cp_elements(28) <= cp_elements(9);
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(28) & cp_elements(32));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7890_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => array_obj_ref_1728_final_reg_req_0); -- 
    base_resize_ack_7878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1728_base_resize_ack_0, ack => cp_elements(30)); -- 
    plus_base_rr_7883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => array_obj_ref_1728_root_address_inst_req_0); -- 
    plus_base_ra_7884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1728_root_address_inst_ack_0, ack => cp_elements(31)); -- 
    plus_base_cr_7885_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_1728_root_address_inst_req_1); -- 
    plus_base_ca_7886_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1728_root_address_inst_ack_1, ack => cp_elements(32)); -- 
    final_reg_ack_7891_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1728_final_reg_ack_0, ack => cp_elements(33)); -- 
    cp_elements(34) <= cp_elements(9);
    cpelement_group_35 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(34) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(35),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => array_obj_ref_1735_final_reg_req_0); -- 
    cp_elements(36) <= cp_elements(23);
    base_resize_req_7902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_1735_base_resize_req_0); -- 
    base_resize_ack_7903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1735_base_resize_ack_0, ack => cp_elements(37)); -- 
    plus_base_rr_7908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_1735_root_address_inst_req_0); -- 
    plus_base_ra_7909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1735_root_address_inst_ack_0, ack => cp_elements(38)); -- 
    plus_base_cr_7910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_1735_root_address_inst_req_1); -- 
    plus_base_ca_7911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1735_root_address_inst_ack_1, ack => cp_elements(39)); -- 
    cp_elements(40) <= array_obj_ref_1735_final_reg_ack_0;
    cpelement_group_41 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(33) & cp_elements(40) & cp_elements(57));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(41),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_7971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_1738_gather_scatter_req_0); -- 
    cp_elements(42) <= cp_elements(40);
    base_resize_req_7930_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_1738_base_resize_req_0); -- 
    base_resize_ack_7931_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_base_resize_ack_0, ack => cp_elements(43)); -- 
    sum_rename_req_7935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_1738_root_address_inst_req_0); -- 
    cp_elements(44) <= ptr_deref_1738_root_address_inst_ack_0;
    cp_elements(45) <= cp_elements(44);
    rr_7943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_1738_addr_0_req_0); -- 
    ra_7944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_0_ack_0, ack => cp_elements(46)); -- 
    cr_7945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_1738_addr_0_req_1); -- 
    ca_7946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_0_ack_1, ack => cp_elements(47)); -- 
    cp_elements(48) <= cp_elements(44);
    rr_7950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_1738_addr_1_req_0); -- 
    ra_7951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_1_ack_0, ack => cp_elements(49)); -- 
    cr_7952_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_1738_addr_1_req_1); -- 
    ca_7953_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_1_ack_1, ack => cp_elements(50)); -- 
    cp_elements(51) <= cp_elements(44);
    rr_7957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => ptr_deref_1738_addr_2_req_0); -- 
    ra_7958_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_2_ack_0, ack => cp_elements(52)); -- 
    cr_7959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => ptr_deref_1738_addr_2_req_1); -- 
    ca_7960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_2_ack_1, ack => cp_elements(53)); -- 
    cp_elements(54) <= cp_elements(44);
    rr_7964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_1738_addr_3_req_0); -- 
    ra_7965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_3_ack_0, ack => cp_elements(55)); -- 
    cr_7966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => ptr_deref_1738_addr_3_req_1); -- 
    ca_7967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_addr_3_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(47) & cp_elements(50) & cp_elements(53) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(58) <= ptr_deref_1738_gather_scatter_ack_0;
    cp_elements(59) <= cp_elements(58);
    rr_7979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => ptr_deref_1738_store_0_req_0); -- 
    ra_7980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_0_ack_0, ack => cp_elements(60)); -- 
    cp_elements(61) <= cp_elements(58);
    rr_7984_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_1738_store_1_req_0); -- 
    ra_7985_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_1_ack_0, ack => cp_elements(62)); -- 
    cp_elements(63) <= cp_elements(58);
    rr_7989_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_1738_store_2_req_0); -- 
    ra_7990_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_2_ack_0, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(58);
    rr_7994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_1738_store_3_req_0); -- 
    ra_7995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_3_ack_0, ack => cp_elements(66)); -- 
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(62) & cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(68) <= cp_elements(67);
    cp_elements(69) <= cp_elements(68);
    cr_8005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_1738_store_0_req_1); -- 
    ca_8006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_0_ack_1, ack => cp_elements(70)); -- 
    cp_elements(71) <= cp_elements(68);
    cr_8010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => ptr_deref_1738_store_1_req_1); -- 
    ca_8011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_1_ack_1, ack => cp_elements(72)); -- 
    cp_elements(73) <= cp_elements(68);
    cr_8015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => ptr_deref_1738_store_2_req_1); -- 
    ca_8016_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_2_ack_1, ack => cp_elements(74)); -- 
    cp_elements(75) <= cp_elements(68);
    cr_8020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => ptr_deref_1738_store_3_req_1); -- 
    ca_8021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1738_store_3_ack_1, ack => cp_elements(76)); -- 
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(72) & cp_elements(74) & cp_elements(76));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_78 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(79) & cp_elements(80));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(78),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => binary_1745_inst_req_0); -- 
    cp_elements(79) <= cp_elements(9);
    cp_elements(80) <= cp_elements(14);
    ra_8031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1745_inst_ack_0, ack => cp_elements(81)); -- 
    cr_8032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => binary_1745_inst_req_1); -- 
    ca_8033_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1745_inst_ack_1, ack => cp_elements(82)); -- 
    cpelement_group_83 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(83),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => type_cast_1749_inst_req_0); -- 
    cp_elements(84) <= cp_elements(9);
    ack_8043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_0, ack => cp_elements(85)); -- 
    cp_elements(86) <= cp_elements(9);
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(86) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8067_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => array_obj_ref_1756_final_reg_req_0); -- 
    cp_elements(88) <= cp_elements(23);
    base_resize_req_8054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => array_obj_ref_1756_base_resize_req_0); -- 
    base_resize_ack_8055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1756_base_resize_ack_0, ack => cp_elements(89)); -- 
    plus_base_rr_8060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => array_obj_ref_1756_root_address_inst_req_0); -- 
    plus_base_ra_8061_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1756_root_address_inst_ack_0, ack => cp_elements(90)); -- 
    plus_base_cr_8062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => array_obj_ref_1756_root_address_inst_req_1); -- 
    plus_base_ca_8063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1756_root_address_inst_ack_1, ack => cp_elements(91)); -- 
    cp_elements(92) <= array_obj_ref_1756_final_reg_ack_0;
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(67) & cp_elements(85) & cp_elements(92) & cp_elements(109));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_1759_gather_scatter_req_0); -- 
    cp_elements(94) <= cp_elements(92);
    base_resize_req_8082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_1759_base_resize_req_0); -- 
    base_resize_ack_8083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_base_resize_ack_0, ack => cp_elements(95)); -- 
    sum_rename_req_8087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => ptr_deref_1759_root_address_inst_req_0); -- 
    cp_elements(96) <= ptr_deref_1759_root_address_inst_ack_0;
    cp_elements(97) <= cp_elements(96);
    rr_8095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => ptr_deref_1759_addr_0_req_0); -- 
    ra_8096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_0_ack_0, ack => cp_elements(98)); -- 
    cr_8097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_1759_addr_0_req_1); -- 
    ca_8098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_0_ack_1, ack => cp_elements(99)); -- 
    cp_elements(100) <= cp_elements(96);
    rr_8102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_1759_addr_1_req_0); -- 
    ra_8103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_1_ack_0, ack => cp_elements(101)); -- 
    cr_8104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_1759_addr_1_req_1); -- 
    ca_8105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_1_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(96);
    rr_8109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_1759_addr_2_req_0); -- 
    ra_8110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_2_ack_0, ack => cp_elements(104)); -- 
    cr_8111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_1759_addr_2_req_1); -- 
    ca_8112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_2_ack_1, ack => cp_elements(105)); -- 
    cp_elements(106) <= cp_elements(96);
    rr_8116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_1759_addr_3_req_0); -- 
    ra_8117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_3_ack_0, ack => cp_elements(107)); -- 
    cr_8118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_1759_addr_3_req_1); -- 
    ca_8119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_addr_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(99) & cp_elements(102) & cp_elements(105) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(110) <= ptr_deref_1759_gather_scatter_ack_0;
    cp_elements(111) <= cp_elements(110);
    rr_8131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_1759_store_0_req_0); -- 
    ra_8132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_0_ack_0, ack => cp_elements(112)); -- 
    cp_elements(113) <= cp_elements(110);
    rr_8136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_1759_store_1_req_0); -- 
    ra_8137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_1_ack_0, ack => cp_elements(114)); -- 
    cp_elements(115) <= cp_elements(110);
    rr_8141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_1759_store_2_req_0); -- 
    ra_8142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_2_ack_0, ack => cp_elements(116)); -- 
    cp_elements(117) <= cp_elements(110);
    rr_8146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_1759_store_3_req_0); -- 
    ra_8147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_3_ack_0, ack => cp_elements(118)); -- 
    cpelement_group_119 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(112) & cp_elements(114) & cp_elements(116) & cp_elements(118));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(120) <= cp_elements(119);
    cp_elements(121) <= cp_elements(120);
    cr_8157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => ptr_deref_1759_store_0_req_1); -- 
    ca_8158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_0_ack_1, ack => cp_elements(122)); -- 
    cp_elements(123) <= cp_elements(120);
    cr_8162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_1759_store_1_req_1); -- 
    ca_8163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_1_ack_1, ack => cp_elements(124)); -- 
    cp_elements(125) <= cp_elements(120);
    cr_8167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_1759_store_2_req_1); -- 
    ca_8168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_2_ack_1, ack => cp_elements(126)); -- 
    cp_elements(127) <= cp_elements(120);
    cr_8172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(127), ack => ptr_deref_1759_store_3_req_1); -- 
    ca_8173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1759_store_3_ack_1, ack => cp_elements(128)); -- 
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(122) & cp_elements(124) & cp_elements(126) & cp_elements(128));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(131) & cp_elements(132));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => binary_1766_inst_req_0); -- 
    cp_elements(131) <= cp_elements(9);
    cp_elements(132) <= cp_elements(14);
    ra_8183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1766_inst_ack_0, ack => cp_elements(133)); -- 
    cr_8184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => binary_1766_inst_req_1); -- 
    ca_8185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1766_inst_ack_1, ack => cp_elements(134)); -- 
    cpelement_group_135 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(135),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8194_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => type_cast_1770_inst_req_0); -- 
    cp_elements(136) <= cp_elements(9);
    cp_elements(137) <= type_cast_1770_inst_ack_0;
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(119) & cp_elements(137) & cp_elements(148));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(139) <= cp_elements(137);
    base_resize_req_8208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => ptr_deref_1774_base_resize_req_0); -- 
    base_resize_ack_8209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_base_resize_ack_0, ack => cp_elements(140)); -- 
    sum_rename_req_8213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_1774_root_address_inst_req_0); -- 
    cp_elements(141) <= ptr_deref_1774_root_address_inst_ack_0;
    cp_elements(142) <= cp_elements(141);
    rr_8221_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_1774_addr_0_req_0); -- 
    ra_8222_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_addr_0_ack_0, ack => cp_elements(143)); -- 
    cr_8223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => ptr_deref_1774_addr_0_req_1); -- 
    ca_8224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_addr_0_ack_1, ack => cp_elements(144)); -- 
    cp_elements(145) <= cp_elements(141);
    rr_8228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => ptr_deref_1774_addr_1_req_0); -- 
    ra_8229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_addr_1_ack_0, ack => cp_elements(146)); -- 
    cr_8230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(146), ack => ptr_deref_1774_addr_1_req_1); -- 
    ca_8231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_addr_1_ack_1, ack => cp_elements(147)); -- 
    cpelement_group_148 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(144) & cp_elements(147));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(148),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(149) <= cp_elements(138);
    rr_8241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_1774_load_0_req_0); -- 
    ra_8242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_load_0_ack_0, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(138);
    rr_8246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_1774_load_1_req_0); -- 
    ra_8247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_load_1_ack_0, ack => cp_elements(152)); -- 
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(150) & cp_elements(152));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(154) <= cp_elements(153);
    cr_8257_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => ptr_deref_1774_load_0_req_1); -- 
    ca_8258_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_load_0_ack_1, ack => cp_elements(155)); -- 
    cp_elements(156) <= cp_elements(153);
    cr_8262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => ptr_deref_1774_load_1_req_1); -- 
    ca_8263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_load_1_ack_1, ack => cp_elements(157)); -- 
    cpelement_group_158 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(155) & cp_elements(157));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_8264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => ptr_deref_1774_gather_scatter_req_0); -- 
    merge_ack_8265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1774_gather_scatter_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(77) & cp_elements(129) & cp_elements(159));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_8276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1778_call_ack_0, ack => cp_elements(161)); -- 
    ccr_8280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => call_stmt_1778_call_req_1); -- 
    cca_8281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1778_call_ack_1, ack => cp_elements(162)); -- 
    cp_elements(163) <= cp_elements(162);
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_1781_inst_req_0); -- 
    cp_elements(165) <= cp_elements(163);
    cp_elements(166) <= cp_elements(163);
    ack_8296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_0, ack => cp_elements(167)); -- 
    index_resize_req_8311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => array_obj_ref_1785_index_0_resize_req_0); -- 
    cp_elements(168) <= cp_elements(163);
    cpelement_group_169 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(168) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(169),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => array_obj_ref_1785_final_reg_req_0); -- 
    cp_elements(170) <= cp_elements(163);
    base_resize_req_8327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => array_obj_ref_1785_base_resize_req_0); -- 
    index_resize_ack_8312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_index_0_resize_ack_0, ack => cp_elements(171)); -- 
    scale_rename_req_8316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => array_obj_ref_1785_index_0_rename_req_0); -- 
    scale_rename_ack_8317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_index_0_rename_ack_0, ack => cp_elements(172)); -- 
    final_index_req_8321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(172), ack => array_obj_ref_1785_offset_inst_req_0); -- 
    final_index_ack_8322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_offset_inst_ack_0, ack => cp_elements(173)); -- 
    base_resize_ack_8328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_base_resize_ack_0, ack => cp_elements(174)); -- 
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(173) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_8333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(175), ack => array_obj_ref_1785_root_address_inst_req_0); -- 
    plus_base_ra_8334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_root_address_inst_ack_0, ack => cp_elements(176)); -- 
    plus_base_cr_8335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => array_obj_ref_1785_root_address_inst_req_1); -- 
    plus_base_ca_8336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_root_address_inst_ack_1, ack => cp_elements(177)); -- 
    final_reg_ack_8341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1785_final_reg_ack_0, ack => cp_elements(178)); -- 
    cp_elements(179) <= cp_elements(163);
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(184));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => array_obj_ref_1792_final_reg_req_0); -- 
    cp_elements(181) <= cp_elements(163);
    base_resize_req_8352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => array_obj_ref_1792_base_resize_req_0); -- 
    base_resize_ack_8353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1792_base_resize_ack_0, ack => cp_elements(182)); -- 
    plus_base_rr_8358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(182), ack => array_obj_ref_1792_root_address_inst_req_0); -- 
    plus_base_ra_8359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1792_root_address_inst_ack_0, ack => cp_elements(183)); -- 
    plus_base_cr_8360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => array_obj_ref_1792_root_address_inst_req_1); -- 
    plus_base_ca_8361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1792_root_address_inst_ack_1, ack => cp_elements(184)); -- 
    cp_elements(185) <= array_obj_ref_1792_final_reg_ack_0;
    cpelement_group_186 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(185) & cp_elements(202));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(186),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => ptr_deref_1795_gather_scatter_req_0); -- 
    cp_elements(187) <= cp_elements(185);
    base_resize_req_8380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => ptr_deref_1795_base_resize_req_0); -- 
    base_resize_ack_8381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_base_resize_ack_0, ack => cp_elements(188)); -- 
    sum_rename_req_8385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => ptr_deref_1795_root_address_inst_req_0); -- 
    cp_elements(189) <= ptr_deref_1795_root_address_inst_ack_0;
    cp_elements(190) <= cp_elements(189);
    rr_8393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_1795_addr_0_req_0); -- 
    ra_8394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_0_ack_0, ack => cp_elements(191)); -- 
    cr_8395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => ptr_deref_1795_addr_0_req_1); -- 
    ca_8396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_0_ack_1, ack => cp_elements(192)); -- 
    cp_elements(193) <= cp_elements(189);
    rr_8400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => ptr_deref_1795_addr_1_req_0); -- 
    ra_8401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_1_ack_0, ack => cp_elements(194)); -- 
    cr_8402_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => ptr_deref_1795_addr_1_req_1); -- 
    ca_8403_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_1_ack_1, ack => cp_elements(195)); -- 
    cp_elements(196) <= cp_elements(189);
    rr_8407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => ptr_deref_1795_addr_2_req_0); -- 
    ra_8408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_2_ack_0, ack => cp_elements(197)); -- 
    cr_8409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => ptr_deref_1795_addr_2_req_1); -- 
    ca_8410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_2_ack_1, ack => cp_elements(198)); -- 
    cp_elements(199) <= cp_elements(189);
    rr_8414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => ptr_deref_1795_addr_3_req_0); -- 
    ra_8415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_3_ack_0, ack => cp_elements(200)); -- 
    cr_8416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => ptr_deref_1795_addr_3_req_1); -- 
    ca_8417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_addr_3_ack_1, ack => cp_elements(201)); -- 
    cpelement_group_202 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(192) & cp_elements(195) & cp_elements(198) & cp_elements(201));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(202),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(203) <= ptr_deref_1795_gather_scatter_ack_0;
    cp_elements(204) <= cp_elements(203);
    rr_8429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_1795_store_0_req_0); -- 
    ra_8430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_0_ack_0, ack => cp_elements(205)); -- 
    cp_elements(206) <= cp_elements(203);
    rr_8434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_1795_store_1_req_0); -- 
    ra_8435_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_1_ack_0, ack => cp_elements(207)); -- 
    cp_elements(208) <= cp_elements(203);
    rr_8439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => ptr_deref_1795_store_2_req_0); -- 
    ra_8440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_2_ack_0, ack => cp_elements(209)); -- 
    cp_elements(210) <= cp_elements(203);
    rr_8444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_1795_store_3_req_0); -- 
    ra_8445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_3_ack_0, ack => cp_elements(211)); -- 
    cpelement_group_212 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(205) & cp_elements(207) & cp_elements(209) & cp_elements(211));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(213) <= cp_elements(212);
    cp_elements(214) <= cp_elements(213);
    cr_8455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => ptr_deref_1795_store_0_req_1); -- 
    ca_8456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_0_ack_1, ack => cp_elements(215)); -- 
    cp_elements(216) <= cp_elements(213);
    cr_8460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(216), ack => ptr_deref_1795_store_1_req_1); -- 
    ca_8461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_1_ack_1, ack => cp_elements(217)); -- 
    cp_elements(218) <= cp_elements(213);
    cr_8465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(218), ack => ptr_deref_1795_store_2_req_1); -- 
    ca_8466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_2_ack_1, ack => cp_elements(219)); -- 
    cp_elements(220) <= cp_elements(213);
    cr_8470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(220), ack => ptr_deref_1795_store_3_req_1); -- 
    ca_8471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1795_store_3_ack_1, ack => cp_elements(221)); -- 
    cpelement_group_222 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(215) & cp_elements(217) & cp_elements(219) & cp_elements(221));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(222),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_223 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(224) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(223),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => binary_1802_inst_req_0); -- 
    cp_elements(224) <= cp_elements(163);
    cp_elements(225) <= cp_elements(163);
    ra_8481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1802_inst_ack_0, ack => cp_elements(226)); -- 
    cr_8482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => binary_1802_inst_req_1); -- 
    ca_8483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1802_inst_ack_1, ack => cp_elements(227)); -- 
    cpelement_group_228 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(227) & cp_elements(229));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(228),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8492_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => binary_1808_inst_req_0); -- 
    cp_elements(229) <= cp_elements(163);
    ra_8493_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1808_inst_ack_0, ack => cp_elements(230)); -- 
    cr_8494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => binary_1808_inst_req_1); -- 
    ca_8495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1808_inst_ack_1, ack => cp_elements(231)); -- 
    cpelement_group_232 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(231) & cp_elements(233));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(232),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(232), ack => type_cast_1812_inst_req_0); -- 
    cp_elements(233) <= cp_elements(163);
    ack_8505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1812_inst_ack_0, ack => cp_elements(234)); -- 
    cp_elements(235) <= cp_elements(163);
    cpelement_group_236 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(235) & cp_elements(240));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(236),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => array_obj_ref_1819_final_reg_req_0); -- 
    cp_elements(237) <= cp_elements(163);
    base_resize_req_8516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => array_obj_ref_1819_base_resize_req_0); -- 
    base_resize_ack_8517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1819_base_resize_ack_0, ack => cp_elements(238)); -- 
    plus_base_rr_8522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => array_obj_ref_1819_root_address_inst_req_0); -- 
    plus_base_ra_8523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1819_root_address_inst_ack_0, ack => cp_elements(239)); -- 
    plus_base_cr_8524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => array_obj_ref_1819_root_address_inst_req_1); -- 
    plus_base_ca_8525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1819_root_address_inst_ack_1, ack => cp_elements(240)); -- 
    cp_elements(241) <= array_obj_ref_1819_final_reg_ack_0;
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(212) & cp_elements(234) & cp_elements(241) & cp_elements(258));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => ptr_deref_1822_gather_scatter_req_0); -- 
    cp_elements(243) <= cp_elements(241);
    base_resize_req_8544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(243), ack => ptr_deref_1822_base_resize_req_0); -- 
    base_resize_ack_8545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_base_resize_ack_0, ack => cp_elements(244)); -- 
    sum_rename_req_8549_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_1822_root_address_inst_req_0); -- 
    cp_elements(245) <= ptr_deref_1822_root_address_inst_ack_0;
    cp_elements(246) <= cp_elements(245);
    rr_8557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_1822_addr_0_req_0); -- 
    ra_8558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_0_ack_0, ack => cp_elements(247)); -- 
    cr_8559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(247), ack => ptr_deref_1822_addr_0_req_1); -- 
    ca_8560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_0_ack_1, ack => cp_elements(248)); -- 
    cp_elements(249) <= cp_elements(245);
    rr_8564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => ptr_deref_1822_addr_1_req_0); -- 
    ra_8565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_1_ack_0, ack => cp_elements(250)); -- 
    cr_8566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_1822_addr_1_req_1); -- 
    ca_8567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_1_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(245);
    rr_8571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_1822_addr_2_req_0); -- 
    ra_8572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_2_ack_0, ack => cp_elements(253)); -- 
    cr_8573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(253), ack => ptr_deref_1822_addr_2_req_1); -- 
    ca_8574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_2_ack_1, ack => cp_elements(254)); -- 
    cp_elements(255) <= cp_elements(245);
    rr_8578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => ptr_deref_1822_addr_3_req_0); -- 
    ra_8579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_3_ack_0, ack => cp_elements(256)); -- 
    cr_8580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => ptr_deref_1822_addr_3_req_1); -- 
    ca_8581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_addr_3_ack_1, ack => cp_elements(257)); -- 
    cpelement_group_258 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(251) & cp_elements(254) & cp_elements(257));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(258),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(259) <= ptr_deref_1822_gather_scatter_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_8593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_1822_store_0_req_0); -- 
    ra_8594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_0_ack_0, ack => cp_elements(261)); -- 
    cp_elements(262) <= cp_elements(259);
    rr_8598_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(262), ack => ptr_deref_1822_store_1_req_0); -- 
    ra_8599_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_1_ack_0, ack => cp_elements(263)); -- 
    cp_elements(264) <= cp_elements(259);
    rr_8603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_1822_store_2_req_0); -- 
    ra_8604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_2_ack_0, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_8608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_1822_store_3_req_0); -- 
    ra_8609_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_3_ack_0, ack => cp_elements(267)); -- 
    cpelement_group_268 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(261) & cp_elements(263) & cp_elements(265) & cp_elements(267));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(268),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(269) <= cp_elements(268);
    cr_8619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_1822_store_0_req_1); -- 
    ca_8620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_0_ack_1, ack => cp_elements(270)); -- 
    cp_elements(271) <= cp_elements(268);
    cr_8624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => ptr_deref_1822_store_1_req_1); -- 
    ca_8625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_1_ack_1, ack => cp_elements(272)); -- 
    cp_elements(273) <= cp_elements(268);
    cr_8629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_1822_store_2_req_1); -- 
    ca_8630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_2_ack_1, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(268);
    cr_8634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_1822_store_3_req_1); -- 
    ca_8635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_3_ack_1, ack => cp_elements(276)); -- 
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(270) & cp_elements(272) & cp_elements(274) & cp_elements(276));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_278 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(222) & cp_elements(277));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(278),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(279) <= cp_elements(2);
    cpelement_group_280 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(281) & cp_elements(282));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(280),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(280), ack => type_cast_1827_inst_req_0); -- 
    cp_elements(281) <= cp_elements(279);
    cp_elements(282) <= cp_elements(279);
    ack_8648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_0, ack => cp_elements(283)); -- 
    pipe_wreq_8653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => simple_obj_ref_1825_inst_req_0); -- 
    pipe_wack_8654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1825_inst_ack_0, ack => cp_elements(284)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1728_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1728_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1728_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1735_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1735_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1735_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1756_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1756_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1756_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1785_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1785_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1785_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1785_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1792_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1792_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1792_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1819_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1819_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1819_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1738_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1738_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1738_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1738_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1738_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1738_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1759_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1759_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1759_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1759_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1759_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1759_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1774_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1774_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1774_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1774_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1774_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1774_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1774_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1774_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1795_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1795_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1795_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1795_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1795_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1795_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1822_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1822_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1822_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1822_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1822_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1822_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1702_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1784_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1784_scaled : std_logic_vector(15 downto 0);
    signal tmp10_1767 : std_logic_vector(31 downto 0);
    signal tmp11_1771 : std_logic_vector(31 downto 0);
    signal tmp12_1775 : std_logic_vector(15 downto 0);
    signal tmp13_1778 : std_logic_vector(15 downto 0);
    signal tmp14_1782 : std_logic_vector(31 downto 0);
    signal tmp15_1786 : std_logic_vector(31 downto 0);
    signal tmp16_1793 : std_logic_vector(31 downto 0);
    signal tmp17_1803 : std_logic_vector(31 downto 0);
    signal tmp18_1809 : std_logic_vector(31 downto 0);
    signal tmp19_1813 : std_logic_vector(31 downto 0);
    signal tmp1_1710 : std_logic_vector(31 downto 0);
    signal tmp20_1820 : std_logic_vector(31 downto 0);
    signal tmp2_1716 : std_logic_vector(31 downto 0);
    signal tmp3_1720 : std_logic_vector(31 downto 0);
    signal tmp4_1724 : std_logic_vector(31 downto 0);
    signal tmp5_1729 : std_logic_vector(31 downto 0);
    signal tmp6_1736 : std_logic_vector(31 downto 0);
    signal tmp7_1746 : std_logic_vector(31 downto 0);
    signal tmp8_1750 : std_logic_vector(31 downto 0);
    signal tmp9_1757 : std_logic_vector(31 downto 0);
    signal tmp_1704 : std_logic_vector(31 downto 0);
    signal type_cast_1708_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1714_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1801_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1807_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1827_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1728_final_offset <= "0000000001101100";
    array_obj_ref_1735_final_offset <= "0000000000001000";
    array_obj_ref_1756_final_offset <= "0000000000001100";
    array_obj_ref_1785_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_1792_final_offset <= "0000000000010000";
    array_obj_ref_1819_final_offset <= "0000000000010100";
    ptr_deref_1738_word_offset_0 <= "0000000000000000";
    ptr_deref_1738_word_offset_1 <= "0000000000000001";
    ptr_deref_1738_word_offset_2 <= "0000000000000010";
    ptr_deref_1738_word_offset_3 <= "0000000000000011";
    ptr_deref_1759_word_offset_0 <= "0000000000000000";
    ptr_deref_1759_word_offset_1 <= "0000000000000001";
    ptr_deref_1759_word_offset_2 <= "0000000000000010";
    ptr_deref_1759_word_offset_3 <= "0000000000000011";
    ptr_deref_1774_word_offset_0 <= "0000000000000000";
    ptr_deref_1774_word_offset_1 <= "0000000000000001";
    ptr_deref_1795_word_offset_0 <= "0000000000000000";
    ptr_deref_1795_word_offset_1 <= "0000000000000001";
    ptr_deref_1795_word_offset_2 <= "0000000000000010";
    ptr_deref_1795_word_offset_3 <= "0000000000000011";
    ptr_deref_1822_word_offset_0 <= "0000000000000000";
    ptr_deref_1822_word_offset_1 <= "0000000000000001";
    ptr_deref_1822_word_offset_2 <= "0000000000000010";
    ptr_deref_1822_word_offset_3 <= "0000000000000011";
    type_cast_1708_wire_constant <= "11111111111111111111100000000000";
    type_cast_1714_wire_constant <= "00000000000000000000000000001000";
    type_cast_1744_wire_constant <= "00000000000000000000000010110100";
    type_cast_1765_wire_constant <= "00000000000000000000000000000110";
    type_cast_1801_wire_constant <= "00000000000000000000011111111111";
    type_cast_1807_wire_constant <= "11111111111111111111111111111000";
    array_obj_ref_1728_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp4_1724, dout => array_obj_ref_1728_resized_base_address, req => array_obj_ref_1728_base_resize_req_0, ack => array_obj_ref_1728_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1728_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1728_root_address, dout => tmp5_1729, req => array_obj_ref_1728_final_reg_req_0, ack => array_obj_ref_1728_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1735_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_1720, dout => array_obj_ref_1735_resized_base_address, req => array_obj_ref_1735_base_resize_req_0, ack => array_obj_ref_1735_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1735_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1735_root_address, dout => tmp6_1736, req => array_obj_ref_1735_final_reg_req_0, ack => array_obj_ref_1735_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1756_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_1720, dout => array_obj_ref_1756_resized_base_address, req => array_obj_ref_1756_base_resize_req_0, ack => array_obj_ref_1756_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1756_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1756_root_address, dout => tmp9_1757, req => array_obj_ref_1756_final_reg_req_0, ack => array_obj_ref_1756_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1785_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_1750, dout => array_obj_ref_1785_resized_base_address, req => array_obj_ref_1785_base_resize_req_0, ack => array_obj_ref_1785_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1785_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1785_root_address, dout => tmp15_1786, req => array_obj_ref_1785_final_reg_req_0, ack => array_obj_ref_1785_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1785_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1782, dout => simple_obj_ref_1784_resized, req => array_obj_ref_1785_index_0_resize_req_0, ack => array_obj_ref_1785_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1785_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_1784_scaled, dout => array_obj_ref_1785_final_offset, req => array_obj_ref_1785_offset_inst_req_0, ack => array_obj_ref_1785_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1792_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_1720, dout => array_obj_ref_1792_resized_base_address, req => array_obj_ref_1792_base_resize_req_0, ack => array_obj_ref_1792_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1792_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1792_root_address, dout => tmp16_1793, req => array_obj_ref_1792_final_reg_req_0, ack => array_obj_ref_1792_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1819_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_1720, dout => array_obj_ref_1819_resized_base_address, req => array_obj_ref_1819_base_resize_req_0, ack => array_obj_ref_1819_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1819_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1819_root_address, dout => tmp20_1820, req => array_obj_ref_1819_final_reg_req_0, ack => array_obj_ref_1819_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1738_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_1736, dout => ptr_deref_1738_resized_base_address, req => ptr_deref_1738_base_resize_req_0, ack => ptr_deref_1738_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1759_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_1757, dout => ptr_deref_1759_resized_base_address, req => ptr_deref_1759_base_resize_req_0, ack => ptr_deref_1759_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1774_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp11_1771, dout => ptr_deref_1774_resized_base_address, req => ptr_deref_1774_base_resize_req_0, ack => ptr_deref_1774_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1795_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1793, dout => ptr_deref_1795_resized_base_address, req => ptr_deref_1795_base_resize_req_0, ack => ptr_deref_1795_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1822_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp20_1820, dout => ptr_deref_1822_resized_base_address, req => ptr_deref_1822_base_resize_req_0, ack => ptr_deref_1822_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1703_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_1702_wire, dout => tmp_1704, req => type_cast_1703_inst_req_0, ack => type_cast_1703_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1719_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_1716, dout => tmp3_1720, req => type_cast_1719_inst_req_0, ack => type_cast_1719_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1723_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_1716, dout => tmp4_1724, req => type_cast_1723_inst_req_0, ack => type_cast_1723_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1749_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_1746, dout => tmp8_1750, req => type_cast_1749_inst_req_0, ack => type_cast_1749_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1770_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_1767, dout => tmp11_1771, req => type_cast_1770_inst_req_0, ack => type_cast_1770_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1781_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_1778, dout => tmp14_1782, req => type_cast_1781_inst_req_0, ack => type_cast_1781_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1812_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp18_1809, dout => tmp19_1813, req => type_cast_1812_inst_req_0, ack => type_cast_1812_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1827_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp2_1716, dout => type_cast_1827_wire, req => type_cast_1827_inst_req_0, ack => type_cast_1827_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1785_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_1785_index_0_rename_ack_0 <= array_obj_ref_1785_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1784_resized;
      simple_obj_ref_1784_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1738_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1738_gather_scatter_ack_0 <= ptr_deref_1738_gather_scatter_req_0;
      aggregated_sig <= tmp5_1729;
      ptr_deref_1738_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1738_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1738_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1738_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1738_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1738_root_address_inst_ack_0 <= ptr_deref_1738_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1738_resized_base_address;
      ptr_deref_1738_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1759_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1759_gather_scatter_ack_0 <= ptr_deref_1759_gather_scatter_req_0;
      aggregated_sig <= tmp8_1750;
      ptr_deref_1759_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1759_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1759_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1759_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1759_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1759_root_address_inst_ack_0 <= ptr_deref_1759_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1759_resized_base_address;
      ptr_deref_1759_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1774_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1774_gather_scatter_ack_0 <= ptr_deref_1774_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1774_data_1 & ptr_deref_1774_data_0;
      tmp12_1775 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1774_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1774_root_address_inst_ack_0 <= ptr_deref_1774_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1774_resized_base_address;
      ptr_deref_1774_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1795_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1795_gather_scatter_ack_0 <= ptr_deref_1795_gather_scatter_req_0;
      aggregated_sig <= tmp15_1786;
      ptr_deref_1795_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1795_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1795_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1795_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1795_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1795_root_address_inst_ack_0 <= ptr_deref_1795_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1795_resized_base_address;
      ptr_deref_1795_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1822_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1822_gather_scatter_ack_0 <= ptr_deref_1822_gather_scatter_req_0;
      aggregated_sig <= tmp19_1813;
      ptr_deref_1822_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1822_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1822_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1822_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1822_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1822_root_address_inst_ack_0 <= ptr_deref_1822_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1822_resized_base_address;
      ptr_deref_1822_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_1728_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1728_resized_base_address;
      array_obj_ref_1728_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001101100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1728_root_address_inst_req_0,
          ackL => array_obj_ref_1728_root_address_inst_ack_0,
          reqR => array_obj_ref_1728_root_address_inst_req_1,
          ackR => array_obj_ref_1728_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1735_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1735_resized_base_address;
      array_obj_ref_1735_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1735_root_address_inst_req_0,
          ackL => array_obj_ref_1735_root_address_inst_ack_0,
          reqR => array_obj_ref_1735_root_address_inst_req_1,
          ackR => array_obj_ref_1735_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1756_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1756_resized_base_address;
      array_obj_ref_1756_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1756_root_address_inst_req_0,
          ackL => array_obj_ref_1756_root_address_inst_ack_0,
          reqR => array_obj_ref_1756_root_address_inst_req_1,
          ackR => array_obj_ref_1756_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1785_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1785_final_offset & array_obj_ref_1785_resized_base_address;
      array_obj_ref_1785_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1785_root_address_inst_req_0,
          ackL => array_obj_ref_1785_root_address_inst_ack_0,
          reqR => array_obj_ref_1785_root_address_inst_req_1,
          ackR => array_obj_ref_1785_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1792_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1792_resized_base_address;
      array_obj_ref_1792_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1792_root_address_inst_req_0,
          ackL => array_obj_ref_1792_root_address_inst_ack_0,
          reqR => array_obj_ref_1792_root_address_inst_req_1,
          ackR => array_obj_ref_1792_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1819_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1819_resized_base_address;
      array_obj_ref_1819_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1819_root_address_inst_req_0,
          ackL => array_obj_ref_1819_root_address_inst_ack_0,
          reqR => array_obj_ref_1819_root_address_inst_req_1,
          ackR => array_obj_ref_1819_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_1709_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1704;
      tmp1_1710 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1709_inst_req_0,
          ackL => binary_1709_inst_ack_0,
          reqR => binary_1709_inst_req_1,
          ackR => binary_1709_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_1715_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_1710;
      tmp2_1716 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1715_inst_req_0,
          ackL => binary_1715_inst_ack_0,
          reqR => binary_1715_inst_req_1,
          ackR => binary_1715_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_1745_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_1710;
      tmp7_1746 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000010110100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1745_inst_req_0,
          ackL => binary_1745_inst_ack_0,
          reqR => binary_1745_inst_req_1,
          ackR => binary_1745_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_1766_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_1710;
      tmp10_1767 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1766_inst_req_0,
          ackL => binary_1766_inst_ack_0,
          reqR => binary_1766_inst_req_1,
          ackR => binary_1766_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_1802_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1704;
      tmp17_1803 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000011111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1802_inst_req_0,
          ackL => binary_1802_inst_ack_0,
          reqR => binary_1802_inst_req_1,
          ackR => binary_1802_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_1808_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp17_1803;
      tmp18_1809 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1808_inst_req_0,
          ackL => binary_1808_inst_ack_0,
          reqR => binary_1808_inst_req_1,
          ackR => binary_1808_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_1738_addr_0 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1738_root_address;
      ptr_deref_1738_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1738_addr_0_req_0,
          ackL => ptr_deref_1738_addr_0_ack_0,
          reqR => ptr_deref_1738_addr_0_req_1,
          ackR => ptr_deref_1738_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_1738_addr_1 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1738_root_address;
      ptr_deref_1738_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1738_addr_1_req_0,
          ackL => ptr_deref_1738_addr_1_ack_0,
          reqR => ptr_deref_1738_addr_1_req_1,
          ackR => ptr_deref_1738_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_1738_addr_2 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1738_root_address;
      ptr_deref_1738_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1738_addr_2_req_0,
          ackL => ptr_deref_1738_addr_2_ack_0,
          reqR => ptr_deref_1738_addr_2_req_1,
          ackR => ptr_deref_1738_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_1738_addr_3 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1738_root_address;
      ptr_deref_1738_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1738_addr_3_req_0,
          ackL => ptr_deref_1738_addr_3_ack_0,
          reqR => ptr_deref_1738_addr_3_req_1,
          ackR => ptr_deref_1738_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_1759_addr_0 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1759_root_address;
      ptr_deref_1759_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1759_addr_0_req_0,
          ackL => ptr_deref_1759_addr_0_ack_0,
          reqR => ptr_deref_1759_addr_0_req_1,
          ackR => ptr_deref_1759_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_1759_addr_1 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1759_root_address;
      ptr_deref_1759_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1759_addr_1_req_0,
          ackL => ptr_deref_1759_addr_1_ack_0,
          reqR => ptr_deref_1759_addr_1_req_1,
          ackR => ptr_deref_1759_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_1759_addr_2 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1759_root_address;
      ptr_deref_1759_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1759_addr_2_req_0,
          ackL => ptr_deref_1759_addr_2_ack_0,
          reqR => ptr_deref_1759_addr_2_req_1,
          ackR => ptr_deref_1759_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_1759_addr_3 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1759_root_address;
      ptr_deref_1759_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1759_addr_3_req_0,
          ackL => ptr_deref_1759_addr_3_ack_0,
          reqR => ptr_deref_1759_addr_3_req_1,
          ackR => ptr_deref_1759_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_1774_addr_0 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1774_root_address;
      ptr_deref_1774_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1774_addr_0_req_0,
          ackL => ptr_deref_1774_addr_0_ack_0,
          reqR => ptr_deref_1774_addr_0_req_1,
          ackR => ptr_deref_1774_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_1774_addr_1 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1774_root_address;
      ptr_deref_1774_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1774_addr_1_req_0,
          ackL => ptr_deref_1774_addr_1_ack_0,
          reqR => ptr_deref_1774_addr_1_req_1,
          ackR => ptr_deref_1774_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_1795_addr_0 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1795_root_address;
      ptr_deref_1795_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1795_addr_0_req_0,
          ackL => ptr_deref_1795_addr_0_ack_0,
          reqR => ptr_deref_1795_addr_0_req_1,
          ackR => ptr_deref_1795_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_1795_addr_1 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1795_root_address;
      ptr_deref_1795_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1795_addr_1_req_0,
          ackL => ptr_deref_1795_addr_1_ack_0,
          reqR => ptr_deref_1795_addr_1_req_1,
          ackR => ptr_deref_1795_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_1795_addr_2 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1795_root_address;
      ptr_deref_1795_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1795_addr_2_req_0,
          ackL => ptr_deref_1795_addr_2_ack_0,
          reqR => ptr_deref_1795_addr_2_req_1,
          ackR => ptr_deref_1795_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_1795_addr_3 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1795_root_address;
      ptr_deref_1795_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1795_addr_3_req_0,
          ackL => ptr_deref_1795_addr_3_ack_0,
          reqR => ptr_deref_1795_addr_3_req_1,
          ackR => ptr_deref_1795_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_1822_addr_0 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1822_root_address;
      ptr_deref_1822_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1822_addr_0_req_0,
          ackL => ptr_deref_1822_addr_0_ack_0,
          reqR => ptr_deref_1822_addr_0_req_1,
          ackR => ptr_deref_1822_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_1822_addr_1 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1822_root_address;
      ptr_deref_1822_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1822_addr_1_req_0,
          ackL => ptr_deref_1822_addr_1_ack_0,
          reqR => ptr_deref_1822_addr_1_req_1,
          ackR => ptr_deref_1822_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_1822_addr_2 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1822_root_address;
      ptr_deref_1822_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1822_addr_2_req_0,
          ackL => ptr_deref_1822_addr_2_ack_0,
          reqR => ptr_deref_1822_addr_2_req_1,
          ackR => ptr_deref_1822_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : ptr_deref_1822_addr_3 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1822_root_address;
      ptr_deref_1822_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1822_addr_3_req_0,
          ackL => ptr_deref_1822_addr_3_ack_0,
          reqR => ptr_deref_1822_addr_3_req_1,
          ackR => ptr_deref_1822_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1774_load_0 ptr_deref_1774_load_1 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1774_load_0_req_0,
        ptr_deref_1774_load_0_ack_0,
        ptr_deref_1774_load_0_req_1,
        ptr_deref_1774_load_0_ack_1,
        "ptr_deref_1774_load_0",
        "memory_space_5" ,
        ptr_deref_1774_data_0,
        ptr_deref_1774_word_address_0,
        "ptr_deref_1774_data_0",
        "ptr_deref_1774_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1774_load_1_req_0,
        ptr_deref_1774_load_1_ack_0,
        ptr_deref_1774_load_1_req_1,
        ptr_deref_1774_load_1_ack_1,
        "ptr_deref_1774_load_1",
        "memory_space_5" ,
        ptr_deref_1774_data_1,
        ptr_deref_1774_word_address_1,
        "ptr_deref_1774_data_1",
        "ptr_deref_1774_word_address_1" -- 
      );
      reqL(1) <= ptr_deref_1774_load_0_req_0;
      reqL(0) <= ptr_deref_1774_load_1_req_0;
      ptr_deref_1774_load_0_ack_0 <= ackL(1);
      ptr_deref_1774_load_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1774_load_0_req_1;
      reqR(0) <= ptr_deref_1774_load_1_req_1;
      ptr_deref_1774_load_0_ack_1 <= ackR(1);
      ptr_deref_1774_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_1774_word_address_0 & ptr_deref_1774_word_address_1;
      ptr_deref_1774_data_0 <= data_out(15 downto 8);
      ptr_deref_1774_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 2,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_1822_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1822_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1822_word_address_1) &  " data ptr_deref_1822_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1822_data_1) severity note; --
        end if;
        if ptr_deref_1759_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1759_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1759_word_address_1) &  " data ptr_deref_1759_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1759_data_1) severity note; --
        end if;
        if ptr_deref_1738_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1738_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1738_word_address_3) &  " data ptr_deref_1738_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1738_data_3) severity note; --
        end if;
        if ptr_deref_1759_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1759_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1759_word_address_2) &  " data ptr_deref_1759_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1759_data_2) severity note; --
        end if;
        if ptr_deref_1795_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1795_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1795_word_address_3) &  " data ptr_deref_1795_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1795_data_3) severity note; --
        end if;
        if ptr_deref_1795_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1795_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1795_word_address_1) &  " data ptr_deref_1795_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1795_data_1) severity note; --
        end if;
        if ptr_deref_1822_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1822_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1822_word_address_0) &  " data ptr_deref_1822_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1822_data_0) severity note; --
        end if;
        if ptr_deref_1738_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1738_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1738_word_address_2) &  " data ptr_deref_1738_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1738_data_2) severity note; --
        end if;
        if ptr_deref_1738_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1738_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1738_word_address_1) &  " data ptr_deref_1738_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1738_data_1) severity note; --
        end if;
        if ptr_deref_1738_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1738_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1738_word_address_0) &  " data ptr_deref_1738_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1738_data_0) severity note; --
        end if;
        if ptr_deref_1822_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1822_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1822_word_address_3) &  " data ptr_deref_1822_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1822_data_3) severity note; --
        end if;
        if ptr_deref_1795_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1795_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1795_word_address_2) &  " data ptr_deref_1795_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1795_data_2) severity note; --
        end if;
        if ptr_deref_1795_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1795_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1795_word_address_0) &  " data ptr_deref_1795_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1795_data_0) severity note; --
        end if;
        if ptr_deref_1759_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1759_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1759_word_address_3) &  " data ptr_deref_1759_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1759_data_3) severity note; --
        end if;
        if ptr_deref_1822_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1822_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1822_word_address_2) &  " data ptr_deref_1822_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1822_data_2) severity note; --
        end if;
        if ptr_deref_1759_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1759_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1759_word_address_0) &  " data ptr_deref_1759_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1759_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1822_store_1 ptr_deref_1759_store_1 ptr_deref_1738_store_3 ptr_deref_1759_store_2 ptr_deref_1795_store_3 ptr_deref_1795_store_1 ptr_deref_1822_store_0 ptr_deref_1738_store_2 ptr_deref_1738_store_1 ptr_deref_1738_store_0 ptr_deref_1822_store_3 ptr_deref_1795_store_2 ptr_deref_1795_store_0 ptr_deref_1759_store_3 ptr_deref_1822_store_2 ptr_deref_1759_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(255 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      -- 
    begin -- 
      reqL(15) <= ptr_deref_1822_store_1_req_0;
      reqL(14) <= ptr_deref_1759_store_1_req_0;
      reqL(13) <= ptr_deref_1738_store_3_req_0;
      reqL(12) <= ptr_deref_1759_store_2_req_0;
      reqL(11) <= ptr_deref_1795_store_3_req_0;
      reqL(10) <= ptr_deref_1795_store_1_req_0;
      reqL(9) <= ptr_deref_1822_store_0_req_0;
      reqL(8) <= ptr_deref_1738_store_2_req_0;
      reqL(7) <= ptr_deref_1738_store_1_req_0;
      reqL(6) <= ptr_deref_1738_store_0_req_0;
      reqL(5) <= ptr_deref_1822_store_3_req_0;
      reqL(4) <= ptr_deref_1795_store_2_req_0;
      reqL(3) <= ptr_deref_1795_store_0_req_0;
      reqL(2) <= ptr_deref_1759_store_3_req_0;
      reqL(1) <= ptr_deref_1822_store_2_req_0;
      reqL(0) <= ptr_deref_1759_store_0_req_0;
      ptr_deref_1822_store_1_ack_0 <= ackL(15);
      ptr_deref_1759_store_1_ack_0 <= ackL(14);
      ptr_deref_1738_store_3_ack_0 <= ackL(13);
      ptr_deref_1759_store_2_ack_0 <= ackL(12);
      ptr_deref_1795_store_3_ack_0 <= ackL(11);
      ptr_deref_1795_store_1_ack_0 <= ackL(10);
      ptr_deref_1822_store_0_ack_0 <= ackL(9);
      ptr_deref_1738_store_2_ack_0 <= ackL(8);
      ptr_deref_1738_store_1_ack_0 <= ackL(7);
      ptr_deref_1738_store_0_ack_0 <= ackL(6);
      ptr_deref_1822_store_3_ack_0 <= ackL(5);
      ptr_deref_1795_store_2_ack_0 <= ackL(4);
      ptr_deref_1795_store_0_ack_0 <= ackL(3);
      ptr_deref_1759_store_3_ack_0 <= ackL(2);
      ptr_deref_1822_store_2_ack_0 <= ackL(1);
      ptr_deref_1759_store_0_ack_0 <= ackL(0);
      reqR(15) <= ptr_deref_1822_store_1_req_1;
      reqR(14) <= ptr_deref_1759_store_1_req_1;
      reqR(13) <= ptr_deref_1738_store_3_req_1;
      reqR(12) <= ptr_deref_1759_store_2_req_1;
      reqR(11) <= ptr_deref_1795_store_3_req_1;
      reqR(10) <= ptr_deref_1795_store_1_req_1;
      reqR(9) <= ptr_deref_1822_store_0_req_1;
      reqR(8) <= ptr_deref_1738_store_2_req_1;
      reqR(7) <= ptr_deref_1738_store_1_req_1;
      reqR(6) <= ptr_deref_1738_store_0_req_1;
      reqR(5) <= ptr_deref_1822_store_3_req_1;
      reqR(4) <= ptr_deref_1795_store_2_req_1;
      reqR(3) <= ptr_deref_1795_store_0_req_1;
      reqR(2) <= ptr_deref_1759_store_3_req_1;
      reqR(1) <= ptr_deref_1822_store_2_req_1;
      reqR(0) <= ptr_deref_1759_store_0_req_1;
      ptr_deref_1822_store_1_ack_1 <= ackR(15);
      ptr_deref_1759_store_1_ack_1 <= ackR(14);
      ptr_deref_1738_store_3_ack_1 <= ackR(13);
      ptr_deref_1759_store_2_ack_1 <= ackR(12);
      ptr_deref_1795_store_3_ack_1 <= ackR(11);
      ptr_deref_1795_store_1_ack_1 <= ackR(10);
      ptr_deref_1822_store_0_ack_1 <= ackR(9);
      ptr_deref_1738_store_2_ack_1 <= ackR(8);
      ptr_deref_1738_store_1_ack_1 <= ackR(7);
      ptr_deref_1738_store_0_ack_1 <= ackR(6);
      ptr_deref_1822_store_3_ack_1 <= ackR(5);
      ptr_deref_1795_store_2_ack_1 <= ackR(4);
      ptr_deref_1795_store_0_ack_1 <= ackR(3);
      ptr_deref_1759_store_3_ack_1 <= ackR(2);
      ptr_deref_1822_store_2_ack_1 <= ackR(1);
      ptr_deref_1759_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1822_word_address_1 & ptr_deref_1759_word_address_1 & ptr_deref_1738_word_address_3 & ptr_deref_1759_word_address_2 & ptr_deref_1795_word_address_3 & ptr_deref_1795_word_address_1 & ptr_deref_1822_word_address_0 & ptr_deref_1738_word_address_2 & ptr_deref_1738_word_address_1 & ptr_deref_1738_word_address_0 & ptr_deref_1822_word_address_3 & ptr_deref_1795_word_address_2 & ptr_deref_1795_word_address_0 & ptr_deref_1759_word_address_3 & ptr_deref_1822_word_address_2 & ptr_deref_1759_word_address_0;
      data_in <= ptr_deref_1822_data_1 & ptr_deref_1759_data_1 & ptr_deref_1738_data_3 & ptr_deref_1759_data_2 & ptr_deref_1795_data_3 & ptr_deref_1795_data_1 & ptr_deref_1822_data_0 & ptr_deref_1738_data_2 & ptr_deref_1738_data_1 & ptr_deref_1738_data_0 & ptr_deref_1822_data_3 & ptr_deref_1795_data_2 & ptr_deref_1795_data_0 & ptr_deref_1759_data_3 & ptr_deref_1822_data_2 & ptr_deref_1759_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 16,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_1702_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_1702_inst_ack_0 then -- 
            assert false report " ReadPipe src_in0 to wire simple_obj_ref_1702_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_1702_inst_req_0;
      simple_obj_ref_1702_inst_ack_0 <= ack(0);
      simple_obj_ref_1702_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => src_in0_pipe_read_req(0),
          oack => src_in0_pipe_read_ack(0),
          odata => src_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1825_inst_ack_0 then -- 
          assert false report " WritePipe chk_in0 from wire type_cast_1827_wire value="  &  convert_slv_to_hex_string(type_cast_1827_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_1825_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1825_inst_req_0;
      simple_obj_ref_1825_inst_ack_0 <= ack(0);
      data_in <= type_cast_1827_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => chk_in0_pipe_write_req(0),
          oack => chk_in0_pipe_write_ack(0),
          odata => chk_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1778_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1778_call_req_0;
      call_stmt_1778_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1778_call_req_1;
      call_stmt_1778_call_ack_1 <= ackR(0);
      data_in <= tmp12_1775;
      tmp13_1778 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 16,
        owidth => 16,
        twidth => 2,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 16, twidth => 2, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to0 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to0_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to0_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to0_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga0_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to0;
architecture Default of ahir_glue_to0 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to0_CP_8663_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_1901_base_resize_req_0 : boolean;
  signal array_obj_ref_1901_base_resize_ack_0 : boolean;
  signal ptr_deref_1905_addr_3_req_1 : boolean;
  signal ptr_deref_1905_addr_3_ack_0 : boolean;
  signal ptr_deref_1905_addr_3_ack_1 : boolean;
  signal ptr_deref_1905_root_address_inst_ack_0 : boolean;
  signal type_cast_1909_inst_ack_0 : boolean;
  signal binary_1914_inst_req_1 : boolean;
  signal binary_1914_inst_ack_1 : boolean;
  signal type_cast_1918_inst_req_0 : boolean;
  signal ptr_deref_1905_load_0_req_0 : boolean;
  signal ptr_deref_1905_load_0_ack_0 : boolean;
  signal type_cast_1918_inst_ack_0 : boolean;
  signal ptr_deref_1905_load_3_req_1 : boolean;
  signal type_cast_1909_inst_req_0 : boolean;
  signal ptr_deref_1905_load_3_ack_1 : boolean;
  signal array_obj_ref_1901_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1901_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1905_load_1_req_0 : boolean;
  signal ptr_deref_1905_load_1_ack_0 : boolean;
  signal ptr_deref_1905_base_resize_req_0 : boolean;
  signal ptr_deref_1905_base_resize_ack_0 : boolean;
  signal ptr_deref_1905_gather_scatter_req_0 : boolean;
  signal ptr_deref_1905_load_0_req_1 : boolean;
  signal ptr_deref_1905_load_2_req_0 : boolean;
  signal ptr_deref_1905_root_address_inst_req_0 : boolean;
  signal type_cast_1894_inst_req_0 : boolean;
  signal ptr_deref_1905_load_0_ack_1 : boolean;
  signal array_obj_ref_1901_root_address_inst_req_1 : boolean;
  signal ptr_deref_1905_load_2_ack_0 : boolean;
  signal type_cast_1894_inst_ack_0 : boolean;
  signal array_obj_ref_1901_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1905_addr_0_req_0 : boolean;
  signal ptr_deref_1905_addr_0_ack_0 : boolean;
  signal ptr_deref_1905_addr_0_req_1 : boolean;
  signal ptr_deref_1905_addr_0_ack_1 : boolean;
  signal ptr_deref_1905_load_3_req_0 : boolean;
  signal ptr_deref_1905_load_1_req_1 : boolean;
  signal ptr_deref_1905_load_1_ack_1 : boolean;
  signal ptr_deref_1905_load_3_ack_0 : boolean;
  signal array_obj_ref_1901_final_reg_req_0 : boolean;
  signal array_obj_ref_1901_final_reg_ack_0 : boolean;
  signal ptr_deref_1905_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1905_addr_1_req_0 : boolean;
  signal ptr_deref_1905_addr_1_ack_0 : boolean;
  signal ptr_deref_1905_addr_1_req_1 : boolean;
  signal ptr_deref_1905_load_2_req_1 : boolean;
  signal ptr_deref_1905_addr_1_ack_1 : boolean;
  signal ptr_deref_1905_addr_2_req_0 : boolean;
  signal ptr_deref_1905_addr_2_ack_0 : boolean;
  signal ptr_deref_1905_addr_2_req_1 : boolean;
  signal ptr_deref_1905_addr_2_ack_1 : boolean;
  signal binary_1914_inst_req_0 : boolean;
  signal binary_1914_inst_ack_0 : boolean;
  signal ptr_deref_1905_load_2_ack_1 : boolean;
  signal ptr_deref_1905_addr_3_req_0 : boolean;
  signal simple_obj_ref_1836_inst_req_0 : boolean;
  signal simple_obj_ref_1836_inst_ack_0 : boolean;
  signal type_cast_1837_inst_req_0 : boolean;
  signal type_cast_1837_inst_ack_0 : boolean;
  signal type_cast_1841_inst_req_0 : boolean;
  signal type_cast_1841_inst_ack_0 : boolean;
  signal binary_1847_inst_req_0 : boolean;
  signal binary_1847_inst_ack_0 : boolean;
  signal binary_1847_inst_req_1 : boolean;
  signal binary_1847_inst_ack_1 : boolean;
  signal type_cast_1851_inst_req_0 : boolean;
  signal type_cast_1851_inst_ack_0 : boolean;
  signal call_stmt_1856_call_req_0 : boolean;
  signal call_stmt_1856_call_ack_0 : boolean;
  signal call_stmt_1856_call_req_1 : boolean;
  signal call_stmt_1856_call_ack_1 : boolean;
  signal ptr_deref_1858_base_resize_req_0 : boolean;
  signal ptr_deref_1858_base_resize_ack_0 : boolean;
  signal ptr_deref_1858_root_address_inst_req_0 : boolean;
  signal ptr_deref_1858_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1858_addr_0_req_0 : boolean;
  signal ptr_deref_1858_addr_0_ack_0 : boolean;
  signal ptr_deref_1858_addr_0_req_1 : boolean;
  signal ptr_deref_1858_addr_0_ack_1 : boolean;
  signal ptr_deref_1858_addr_1_req_0 : boolean;
  signal ptr_deref_1858_addr_1_ack_0 : boolean;
  signal ptr_deref_1858_addr_1_req_1 : boolean;
  signal ptr_deref_1858_addr_1_ack_1 : boolean;
  signal ptr_deref_1858_gather_scatter_req_0 : boolean;
  signal ptr_deref_1858_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1858_store_0_req_0 : boolean;
  signal ptr_deref_1858_store_0_ack_0 : boolean;
  signal ptr_deref_1858_store_1_req_0 : boolean;
  signal ptr_deref_1858_store_1_ack_0 : boolean;
  signal ptr_deref_1858_store_0_req_1 : boolean;
  signal ptr_deref_1858_store_0_ack_1 : boolean;
  signal ptr_deref_1858_store_1_req_1 : boolean;
  signal ptr_deref_1858_store_1_ack_1 : boolean;
  signal binary_1865_inst_req_0 : boolean;
  signal binary_1865_inst_ack_0 : boolean;
  signal binary_1865_inst_req_1 : boolean;
  signal binary_1865_inst_ack_1 : boolean;
  signal type_cast_1869_inst_req_0 : boolean;
  signal type_cast_1869_inst_ack_0 : boolean;
  signal binary_1875_inst_req_0 : boolean;
  signal binary_1875_inst_ack_0 : boolean;
  signal binary_1875_inst_req_1 : boolean;
  signal binary_1875_inst_ack_1 : boolean;
  signal type_cast_1879_inst_req_0 : boolean;
  signal type_cast_1879_inst_ack_0 : boolean;
  signal array_obj_ref_1886_base_resize_req_0 : boolean;
  signal array_obj_ref_1886_base_resize_ack_0 : boolean;
  signal array_obj_ref_1886_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1886_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1886_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1886_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1886_final_reg_req_0 : boolean;
  signal array_obj_ref_1886_final_reg_ack_0 : boolean;
  signal ptr_deref_1890_base_resize_req_0 : boolean;
  signal ptr_deref_1890_base_resize_ack_0 : boolean;
  signal ptr_deref_1890_root_address_inst_req_0 : boolean;
  signal ptr_deref_1890_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1890_addr_0_req_0 : boolean;
  signal ptr_deref_1890_addr_0_ack_0 : boolean;
  signal ptr_deref_1890_addr_0_req_1 : boolean;
  signal ptr_deref_1890_addr_0_ack_1 : boolean;
  signal ptr_deref_1890_addr_1_req_0 : boolean;
  signal ptr_deref_1890_addr_1_ack_0 : boolean;
  signal ptr_deref_1890_addr_1_req_1 : boolean;
  signal ptr_deref_1890_addr_1_ack_1 : boolean;
  signal ptr_deref_1890_addr_2_req_0 : boolean;
  signal ptr_deref_1890_addr_2_ack_0 : boolean;
  signal ptr_deref_1890_addr_2_req_1 : boolean;
  signal ptr_deref_1890_addr_2_ack_1 : boolean;
  signal ptr_deref_1890_addr_3_req_0 : boolean;
  signal ptr_deref_1890_addr_3_ack_0 : boolean;
  signal ptr_deref_1890_addr_3_req_1 : boolean;
  signal ptr_deref_1890_addr_3_ack_1 : boolean;
  signal ptr_deref_1890_load_0_req_0 : boolean;
  signal ptr_deref_1890_load_0_ack_0 : boolean;
  signal ptr_deref_1890_load_1_req_0 : boolean;
  signal ptr_deref_1890_load_1_ack_0 : boolean;
  signal ptr_deref_1890_load_2_req_0 : boolean;
  signal ptr_deref_1890_load_2_ack_0 : boolean;
  signal ptr_deref_1890_load_3_req_0 : boolean;
  signal ptr_deref_1890_load_3_ack_0 : boolean;
  signal ptr_deref_1890_load_0_req_1 : boolean;
  signal ptr_deref_1890_load_0_ack_1 : boolean;
  signal ptr_deref_1890_load_1_req_1 : boolean;
  signal ptr_deref_1890_load_1_ack_1 : boolean;
  signal ptr_deref_1890_load_2_req_1 : boolean;
  signal ptr_deref_1890_load_2_ack_1 : boolean;
  signal ptr_deref_1890_load_3_req_1 : boolean;
  signal ptr_deref_1890_load_3_ack_1 : boolean;
  signal ptr_deref_1890_gather_scatter_req_0 : boolean;
  signal ptr_deref_1890_gather_scatter_ack_0 : boolean;
  signal binary_1924_inst_req_0 : boolean;
  signal binary_1924_inst_ack_0 : boolean;
  signal binary_1924_inst_req_1 : boolean;
  signal binary_1924_inst_ack_1 : boolean;
  signal type_cast_1928_inst_req_0 : boolean;
  signal type_cast_1928_inst_ack_0 : boolean;
  signal binary_1934_inst_req_0 : boolean;
  signal binary_1934_inst_ack_0 : boolean;
  signal binary_1934_inst_req_1 : boolean;
  signal binary_1934_inst_ack_1 : boolean;
  signal binary_1940_inst_req_0 : boolean;
  signal binary_1940_inst_ack_0 : boolean;
  signal binary_1940_inst_req_1 : boolean;
  signal binary_1940_inst_ack_1 : boolean;
  signal type_cast_1944_inst_req_0 : boolean;
  signal type_cast_1944_inst_ack_0 : boolean;
  signal binary_1948_inst_req_0 : boolean;
  signal binary_1948_inst_ack_0 : boolean;
  signal binary_1948_inst_req_1 : boolean;
  signal binary_1948_inst_ack_1 : boolean;
  signal type_cast_1952_inst_req_0 : boolean;
  signal type_cast_1952_inst_ack_0 : boolean;
  signal binary_1957_inst_req_0 : boolean;
  signal binary_1957_inst_ack_0 : boolean;
  signal binary_1957_inst_req_1 : boolean;
  signal binary_1957_inst_ack_1 : boolean;
  signal call_stmt_1961_call_req_0 : boolean;
  signal call_stmt_1961_call_ack_0 : boolean;
  signal call_stmt_1961_call_req_1 : boolean;
  signal call_stmt_1961_call_ack_1 : boolean;
  signal ptr_deref_1963_base_resize_req_0 : boolean;
  signal ptr_deref_1963_base_resize_ack_0 : boolean;
  signal ptr_deref_1963_root_address_inst_req_0 : boolean;
  signal ptr_deref_1963_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1963_addr_0_req_0 : boolean;
  signal ptr_deref_1963_addr_0_ack_0 : boolean;
  signal ptr_deref_1963_addr_0_req_1 : boolean;
  signal ptr_deref_1963_addr_0_ack_1 : boolean;
  signal ptr_deref_1963_addr_1_req_0 : boolean;
  signal ptr_deref_1963_addr_1_ack_0 : boolean;
  signal ptr_deref_1963_addr_1_req_1 : boolean;
  signal ptr_deref_1963_addr_1_ack_1 : boolean;
  signal ptr_deref_1963_gather_scatter_req_0 : boolean;
  signal ptr_deref_1963_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1963_store_0_req_0 : boolean;
  signal ptr_deref_1963_store_0_ack_0 : boolean;
  signal ptr_deref_1963_store_1_req_0 : boolean;
  signal ptr_deref_1963_store_1_ack_0 : boolean;
  signal ptr_deref_1963_store_0_req_1 : boolean;
  signal ptr_deref_1963_store_0_ack_1 : boolean;
  signal ptr_deref_1963_store_1_req_1 : boolean;
  signal ptr_deref_1963_store_1_ack_1 : boolean;
  signal call_stmt_1968_call_req_0 : boolean;
  signal call_stmt_1968_call_ack_0 : boolean;
  signal call_stmt_1968_call_req_1 : boolean;
  signal call_stmt_1968_call_ack_1 : boolean;
  signal ptr_deref_1970_base_resize_req_0 : boolean;
  signal ptr_deref_1970_base_resize_ack_0 : boolean;
  signal ptr_deref_1970_root_address_inst_req_0 : boolean;
  signal ptr_deref_1970_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1970_addr_0_req_0 : boolean;
  signal ptr_deref_1970_addr_0_ack_0 : boolean;
  signal ptr_deref_1970_addr_0_req_1 : boolean;
  signal ptr_deref_1970_addr_0_ack_1 : boolean;
  signal ptr_deref_1970_addr_1_req_0 : boolean;
  signal ptr_deref_1970_addr_1_ack_0 : boolean;
  signal ptr_deref_1970_addr_1_req_1 : boolean;
  signal ptr_deref_1970_addr_1_ack_1 : boolean;
  signal ptr_deref_1970_gather_scatter_req_0 : boolean;
  signal ptr_deref_1970_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1970_store_0_req_0 : boolean;
  signal ptr_deref_1970_store_0_ack_0 : boolean;
  signal ptr_deref_1970_store_1_req_0 : boolean;
  signal ptr_deref_1970_store_1_ack_0 : boolean;
  signal ptr_deref_1970_store_0_req_1 : boolean;
  signal ptr_deref_1970_store_0_ack_1 : boolean;
  signal ptr_deref_1970_store_1_req_1 : boolean;
  signal ptr_deref_1970_store_1_ack_1 : boolean;
  signal ptr_deref_1975_base_resize_req_0 : boolean;
  signal ptr_deref_1975_base_resize_ack_0 : boolean;
  signal ptr_deref_1975_root_address_inst_req_0 : boolean;
  signal ptr_deref_1975_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1975_addr_0_req_0 : boolean;
  signal ptr_deref_1975_addr_0_ack_0 : boolean;
  signal ptr_deref_1975_addr_0_req_1 : boolean;
  signal ptr_deref_1975_addr_0_ack_1 : boolean;
  signal ptr_deref_1975_addr_1_req_0 : boolean;
  signal ptr_deref_1975_addr_1_ack_0 : boolean;
  signal ptr_deref_1975_addr_1_req_1 : boolean;
  signal ptr_deref_1975_addr_1_ack_1 : boolean;
  signal ptr_deref_1975_addr_2_req_0 : boolean;
  signal ptr_deref_1975_addr_2_ack_0 : boolean;
  signal ptr_deref_1975_addr_2_req_1 : boolean;
  signal ptr_deref_1975_addr_2_ack_1 : boolean;
  signal ptr_deref_1975_addr_3_req_0 : boolean;
  signal ptr_deref_1975_addr_3_ack_0 : boolean;
  signal ptr_deref_1975_addr_3_req_1 : boolean;
  signal ptr_deref_1975_addr_3_ack_1 : boolean;
  signal ptr_deref_1975_load_0_req_0 : boolean;
  signal ptr_deref_1975_load_0_ack_0 : boolean;
  signal ptr_deref_1975_load_1_req_0 : boolean;
  signal ptr_deref_1975_load_1_ack_0 : boolean;
  signal ptr_deref_1975_load_2_req_0 : boolean;
  signal ptr_deref_1975_load_2_ack_0 : boolean;
  signal ptr_deref_1975_load_3_req_0 : boolean;
  signal ptr_deref_1975_load_3_ack_0 : boolean;
  signal ptr_deref_1975_load_0_req_1 : boolean;
  signal ptr_deref_1975_load_0_ack_1 : boolean;
  signal ptr_deref_1975_load_1_req_1 : boolean;
  signal ptr_deref_1975_load_1_ack_1 : boolean;
  signal ptr_deref_1975_load_2_req_1 : boolean;
  signal ptr_deref_1975_load_2_ack_1 : boolean;
  signal ptr_deref_1975_load_3_req_1 : boolean;
  signal ptr_deref_1975_load_3_ack_1 : boolean;
  signal ptr_deref_1975_gather_scatter_req_0 : boolean;
  signal ptr_deref_1975_gather_scatter_ack_0 : boolean;
  signal type_cast_1979_inst_req_0 : boolean;
  signal type_cast_1979_inst_ack_0 : boolean;
  signal simple_obj_ref_1981_inst_req_0 : boolean;
  signal simple_obj_ref_1981_inst_ack_0 : boolean;
  signal type_cast_1987_inst_req_0 : boolean;
  signal type_cast_1987_inst_ack_0 : boolean;
  signal simple_obj_ref_1985_inst_req_0 : boolean;
  signal simple_obj_ref_1985_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to0_CP_8663: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_8754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_1856_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_9279_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_1961_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_9577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_1981_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8709_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_1837_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_8704_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_1836_inst_req_0); -- 
    ack_8705_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1836_inst_ack_0, ack => cp_elements(8)); -- 
    ack_8710_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_1841_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_8723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1841_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_1847_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_8733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1847_inst_ack_0, ack => cp_elements(18)); -- 
    cr_8734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_1847_inst_req_1); -- 
    ca_8735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1847_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_1851_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_8745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1851_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_8755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1856_call_ack_0, ack => cp_elements(24)); -- 
    ccr_8759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_1856_call_req_1); -- 
    cca_8760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1856_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_1858_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_8779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_1858_base_resize_req_0); -- 
    base_resize_ack_8780_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_8784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_1858_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_1858_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_8792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_1858_addr_0_req_0); -- 
    ra_8793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_8794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_1858_addr_0_req_1); -- 
    ca_8795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_8799_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_1858_addr_1_req_0); -- 
    ra_8800_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_8801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_1858_addr_1_req_1); -- 
    ca_8802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_1858_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_8814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_1858_store_0_req_0); -- 
    ra_8815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_8819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_1858_store_1_req_0); -- 
    ra_8820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_8830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_1858_store_0_req_1); -- 
    ca_8831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_8835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_1858_store_1_req_1); -- 
    ca_8836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1858_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_1865_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_8846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1865_inst_ack_0, ack => cp_elements(55)); -- 
    cr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_1865_inst_req_1); -- 
    ca_8848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1865_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_1869_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_8858_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1869_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_1875_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_8868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1875_inst_ack_0, ack => cp_elements(63)); -- 
    cr_8869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_1875_inst_req_1); -- 
    ca_8870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1875_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_1879_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_8880_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1879_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_1886_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_8891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_1886_base_resize_req_0); -- 
    base_resize_ack_8892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1886_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_8897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_1886_root_address_inst_req_0); -- 
    plus_base_ra_8898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1886_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_8899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_1886_root_address_inst_req_1); -- 
    plus_base_ca_8900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1886_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_1886_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_8918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_1890_base_resize_req_0); -- 
    base_resize_ack_8919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_8923_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_1890_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_1890_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_8931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_1890_addr_0_req_0); -- 
    ra_8932_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_8933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_1890_addr_0_req_1); -- 
    ca_8934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_8938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_1890_addr_1_req_0); -- 
    ra_8939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_8940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_1890_addr_1_req_1); -- 
    ca_8941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_8945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_1890_addr_2_req_0); -- 
    ra_8946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_8947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_1890_addr_2_req_1); -- 
    ca_8948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_8952_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_1890_addr_3_req_0); -- 
    ra_8953_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_8954_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_1890_addr_3_req_1); -- 
    ca_8955_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_8965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_1890_load_0_req_0); -- 
    ra_8966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_8970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_1890_load_1_req_0); -- 
    ra_8971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_8975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_1890_load_2_req_0); -- 
    ra_8976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_8980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_1890_load_3_req_0); -- 
    ra_8981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_8991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_1890_load_0_req_1); -- 
    ca_8992_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_8996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_1890_load_1_req_1); -- 
    ca_8997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_9001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_1890_load_2_req_1); -- 
    ca_9002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_9006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_1890_load_3_req_1); -- 
    ca_9007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_1890_gather_scatter_req_0); -- 
    merge_ack_9009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1890_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_1894_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_9019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_9043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_1901_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_9030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_1901_base_resize_req_0); -- 
    base_resize_ack_9031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1901_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_9036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_1901_root_address_inst_req_0); -- 
    plus_base_ra_9037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1901_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_9038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_1901_root_address_inst_req_1); -- 
    plus_base_ca_9039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1901_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_1901_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_9057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_1905_base_resize_req_0); -- 
    base_resize_ack_9058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_9062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_1905_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_1905_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_9070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_1905_addr_0_req_0); -- 
    ra_9071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_9072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_1905_addr_0_req_1); -- 
    ca_9073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_9077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_1905_addr_1_req_0); -- 
    ra_9078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_9079_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_1905_addr_1_req_1); -- 
    ca_9080_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_9084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_1905_addr_2_req_0); -- 
    ra_9085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_9086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_1905_addr_2_req_1); -- 
    ca_9087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_9091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_1905_addr_3_req_0); -- 
    ra_9092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_9093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_1905_addr_3_req_1); -- 
    ca_9094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_9104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_1905_load_0_req_0); -- 
    ra_9105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_9109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_1905_load_1_req_0); -- 
    ra_9110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_9114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_1905_load_2_req_0); -- 
    ra_9115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_9119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_1905_load_3_req_0); -- 
    ra_9120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_9130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_1905_load_0_req_1); -- 
    ca_9131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_9135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_1905_load_1_req_1); -- 
    ca_9136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_9140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_1905_load_2_req_1); -- 
    ca_9141_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_9145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_1905_load_3_req_1); -- 
    ca_9146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_1905_gather_scatter_req_0); -- 
    merge_ack_9148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_1909_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_9158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1909_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_1914_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_9169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1914_inst_ack_0, ack => cp_elements(162)); -- 
    cr_9170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_1914_inst_req_1); -- 
    cp_elements(163) <= binary_1914_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_1918_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_9181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1918_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_1924_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_9191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1924_inst_ack_0, ack => cp_elements(171)); -- 
    cr_9192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_1924_inst_req_1); -- 
    ca_9193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1924_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9202_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_1928_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_9203_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1928_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_1934_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_9213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1934_inst_ack_0, ack => cp_elements(178)); -- 
    cr_9214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_1934_inst_req_1); -- 
    ca_9215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1934_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_1940_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_9225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1940_inst_ack_0, ack => cp_elements(183)); -- 
    cr_9226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_1940_inst_req_1); -- 
    ca_9227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1940_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_1948_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_1944_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_9239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_0, ack => cp_elements(189)); -- 
    ra_9244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1948_inst_ack_0, ack => cp_elements(190)); -- 
    cr_9245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_1948_inst_req_1); -- 
    ca_9246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1948_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9255_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_1952_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_9256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1952_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_1957_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_9267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1957_inst_ack_0, ack => cp_elements(197)); -- 
    cr_9268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_1957_inst_req_1); -- 
    ca_9269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1957_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_9280_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1961_call_ack_0, ack => cp_elements(200)); -- 
    ccr_9284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_1961_call_req_1); -- 
    cca_9285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1961_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_9331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_1963_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_9304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_1963_base_resize_req_0); -- 
    base_resize_ack_9305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_9309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_1963_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_1963_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_9317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_1963_addr_0_req_0); -- 
    ra_9318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_9319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_1963_addr_0_req_1); -- 
    ca_9320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_9324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_1963_addr_1_req_0); -- 
    ra_9325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_9326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_1963_addr_1_req_1); -- 
    ca_9327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_1963_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_9339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_1963_store_0_req_0); -- 
    ra_9340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_9344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_1963_store_1_req_0); -- 
    ra_9345_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_9355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_1963_store_0_req_1); -- 
    ca_9356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_9360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_1963_store_1_req_1); -- 
    ca_9361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_9371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_1968_call_req_0); -- 
    cra_9372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1968_call_ack_0, ack => cp_elements(227)); -- 
    ccr_9376_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_1968_call_req_1); -- 
    cca_9377_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1968_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_9423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_1970_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_9396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_1970_base_resize_req_0); -- 
    base_resize_ack_9397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_9401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_1970_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_1970_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_9409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_1970_addr_0_req_0); -- 
    ra_9410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_9411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_1970_addr_0_req_1); -- 
    ca_9412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_9416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_1970_addr_1_req_0); -- 
    ra_9417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_9418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_1970_addr_1_req_1); -- 
    ca_9419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_1970_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_9431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_1970_store_0_req_0); -- 
    ra_9432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_9436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_1970_store_1_req_0); -- 
    ra_9437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_9447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_1970_store_0_req_1); -- 
    ca_9448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_9452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_1970_store_1_req_1); -- 
    ca_9453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1970_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_9466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_1975_base_resize_req_0); -- 
    base_resize_ack_9467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_9471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_1975_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_1975_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_9479_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_1975_addr_0_req_0); -- 
    ra_9480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_9481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_1975_addr_0_req_1); -- 
    ca_9482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_9486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_1975_addr_1_req_0); -- 
    ra_9487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_9488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_1975_addr_1_req_1); -- 
    ca_9489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_9493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_1975_addr_2_req_0); -- 
    ra_9494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_9495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_1975_addr_2_req_1); -- 
    ca_9496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_9500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_1975_addr_3_req_0); -- 
    ra_9501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_9502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_1975_addr_3_req_1); -- 
    ca_9503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_9513_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_1975_load_0_req_0); -- 
    ra_9514_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_9518_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_1975_load_1_req_0); -- 
    ra_9519_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_9523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_1975_load_2_req_0); -- 
    ra_9524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_9528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_1975_load_3_req_0); -- 
    ra_9529_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_9539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_1975_load_0_req_1); -- 
    ca_9540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_9544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_1975_load_1_req_1); -- 
    ca_9545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_9549_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_1975_load_2_req_1); -- 
    ca_9550_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_9554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_1975_load_3_req_1); -- 
    ca_9555_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_1975_gather_scatter_req_0); -- 
    merge_ack_9557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1975_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_1979_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_9567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_9578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1981_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_1987_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_9591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_9596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_1985_inst_req_0); -- 
    pipe_wack_9597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1985_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1886_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1886_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1886_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1901_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1901_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1901_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_1949 : std_logic_vector(0 downto 0);
    signal ptr_deref_1858_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1858_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1858_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1858_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1858_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_1858_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1858_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1858_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1858_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1890_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1890_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1890_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1890_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1890_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1905_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1905_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1905_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1905_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1905_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1963_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1963_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1963_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1970_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1970_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1970_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1975_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1975_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1975_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1975_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1975_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1836_wire : std_logic_vector(31 downto 0);
    signal tmp10_1891 : std_logic_vector(31 downto 0);
    signal tmp11_1895 : std_logic_vector(31 downto 0);
    signal tmp12_1902 : std_logic_vector(31 downto 0);
    signal tmp13_1906 : std_logic_vector(31 downto 0);
    signal tmp14_1910 : std_logic_vector(31 downto 0);
    signal tmp15_1915 : std_logic_vector(31 downto 0);
    signal tmp16_1919 : std_logic_vector(15 downto 0);
    signal tmp17_1925 : std_logic_vector(31 downto 0);
    signal tmp18_1935 : std_logic_vector(15 downto 0);
    signal tmp19_1941 : std_logic_vector(31 downto 0);
    signal tmp1_1842 : std_logic_vector(31 downto 0);
    signal tmp20_1953 : std_logic_vector(15 downto 0);
    signal tmp21_1958 : std_logic_vector(15 downto 0);
    signal tmp22_1961 : std_logic_vector(15 downto 0);
    signal tmp23_1968 : std_logic_vector(15 downto 0);
    signal tmp24_1976 : std_logic_vector(31 downto 0);
    signal tmp25_1980 : std_logic_vector(31 downto 0);
    signal tmp2_1848 : std_logic_vector(31 downto 0);
    signal tmp3_1852 : std_logic_vector(31 downto 0);
    signal tmp4_1856 : std_logic_vector(15 downto 0);
    signal tmp5_1866 : std_logic_vector(31 downto 0);
    signal tmp6_1870 : std_logic_vector(31 downto 0);
    signal tmp7_1876 : std_logic_vector(31 downto 0);
    signal tmp8_1880 : std_logic_vector(31 downto 0);
    signal tmp9_1887 : std_logic_vector(31 downto 0);
    signal tmp_1838 : std_logic_vector(31 downto 0);
    signal type_cast_1846_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1854_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1864_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1923_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1933_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1939_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1944_wire : std_logic_vector(31 downto 0);
    signal type_cast_1947_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1983_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1987_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_1929 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1886_final_offset <= "0000000000010000";
    array_obj_ref_1901_final_offset <= "0000000000001100";
    ptr_deref_1858_word_offset_0 <= "0000000000000000";
    ptr_deref_1858_word_offset_1 <= "0000000000000001";
    ptr_deref_1890_word_offset_0 <= "0000000000000000";
    ptr_deref_1890_word_offset_1 <= "0000000000000001";
    ptr_deref_1890_word_offset_2 <= "0000000000000010";
    ptr_deref_1890_word_offset_3 <= "0000000000000011";
    ptr_deref_1905_word_offset_0 <= "0000000000000000";
    ptr_deref_1905_word_offset_1 <= "0000000000000001";
    ptr_deref_1905_word_offset_2 <= "0000000000000010";
    ptr_deref_1905_word_offset_3 <= "0000000000000011";
    ptr_deref_1963_word_offset_0 <= "0000000000000000";
    ptr_deref_1963_word_offset_1 <= "0000000000000001";
    ptr_deref_1970_word_offset_0 <= "0000000000000000";
    ptr_deref_1970_word_offset_1 <= "0000000000000001";
    ptr_deref_1975_word_offset_0 <= "0000000000000000";
    ptr_deref_1975_word_offset_1 <= "0000000000000001";
    ptr_deref_1975_word_offset_2 <= "0000000000000010";
    ptr_deref_1975_word_offset_3 <= "0000000000000011";
    type_cast_1846_wire_constant <= "11111111111111111111100000000000";
    type_cast_1854_wire_constant <= "0000000000000001";
    type_cast_1864_wire_constant <= "00000000000000000000000000000110";
    type_cast_1874_wire_constant <= "00000000000000000000000000000010";
    type_cast_1923_wire_constant <= "00000000000000000000000000000011";
    type_cast_1933_wire_constant <= "0001111111111111";
    type_cast_1939_wire_constant <= "00000000000000000000000000000111";
    type_cast_1947_wire_constant <= "00000000000000000000000000000000";
    type_cast_1983_wire_constant <= "00000000000000000000000000000001";
    array_obj_ref_1886_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_1842, dout => array_obj_ref_1886_resized_base_address, req => array_obj_ref_1886_base_resize_req_0, ack => array_obj_ref_1886_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1886_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1886_root_address, dout => tmp9_1887, req => array_obj_ref_1886_final_reg_req_0, ack => array_obj_ref_1886_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1901_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_1842, dout => array_obj_ref_1901_resized_base_address, req => array_obj_ref_1901_base_resize_req_0, ack => array_obj_ref_1901_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1901_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1901_root_address, dout => tmp12_1902, req => array_obj_ref_1901_final_reg_req_0, ack => array_obj_ref_1901_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1858_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_1852, dout => ptr_deref_1858_resized_base_address, req => ptr_deref_1858_base_resize_req_0, ack => ptr_deref_1858_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1890_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_1887, dout => ptr_deref_1890_resized_base_address, req => ptr_deref_1890_base_resize_req_0, ack => ptr_deref_1890_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1905_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_1902, dout => ptr_deref_1905_resized_base_address, req => ptr_deref_1905_base_resize_req_0, ack => ptr_deref_1905_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1963_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_1870, dout => ptr_deref_1963_resized_base_address, req => ptr_deref_1963_base_resize_req_0, ack => ptr_deref_1963_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1970_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_1880, dout => ptr_deref_1970_resized_base_address, req => ptr_deref_1970_base_resize_req_0, ack => ptr_deref_1970_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1975_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_1902, dout => ptr_deref_1975_resized_base_address, req => ptr_deref_1975_base_resize_req_0, ack => ptr_deref_1975_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1837_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_1836_wire, dout => tmp_1838, req => type_cast_1837_inst_req_0, ack => type_cast_1837_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1841_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_1838, dout => tmp1_1842, req => type_cast_1841_inst_req_0, ack => type_cast_1841_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1851_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_1848, dout => tmp3_1852, req => type_cast_1851_inst_req_0, ack => type_cast_1851_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1869_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_1866, dout => tmp6_1870, req => type_cast_1869_inst_req_0, ack => type_cast_1869_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1879_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_1876, dout => tmp8_1880, req => type_cast_1879_inst_req_0, ack => type_cast_1879_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1894_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_1891, dout => tmp11_1895, req => type_cast_1894_inst_req_0, ack => type_cast_1894_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1909_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_1906, dout => tmp14_1910, req => type_cast_1909_inst_req_0, ack => type_cast_1909_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1918_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_1915, dout => tmp16_1919, req => type_cast_1918_inst_req_0, ack => type_cast_1918_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1928_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_1925, dout => xx_xtrx_xi_1929, req => type_cast_1928_inst_req_0, ack => type_cast_1928_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1944_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_1941, dout => type_cast_1944_wire, req => type_cast_1944_inst_req_0, ack => type_cast_1944_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1952_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_1949, dout => tmp20_1953, req => type_cast_1952_inst_req_0, ack => type_cast_1952_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1979_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_1976, dout => tmp25_1980, req => type_cast_1979_inst_req_0, ack => type_cast_1979_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1987_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_1980, dout => type_cast_1987_wire, req => type_cast_1987_inst_req_0, ack => type_cast_1987_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1858_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1858_gather_scatter_ack_0 <= ptr_deref_1858_gather_scatter_req_0;
      aggregated_sig <= tmp4_1856;
      ptr_deref_1858_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1858_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1858_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1858_root_address_inst_ack_0 <= ptr_deref_1858_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1858_resized_base_address;
      ptr_deref_1858_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1890_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1890_gather_scatter_ack_0 <= ptr_deref_1890_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1890_data_3 & ptr_deref_1890_data_2 & ptr_deref_1890_data_1 & ptr_deref_1890_data_0;
      tmp10_1891 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1890_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1890_root_address_inst_ack_0 <= ptr_deref_1890_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1890_resized_base_address;
      ptr_deref_1890_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1905_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1905_gather_scatter_ack_0 <= ptr_deref_1905_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1905_data_3 & ptr_deref_1905_data_2 & ptr_deref_1905_data_1 & ptr_deref_1905_data_0;
      tmp13_1906 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1905_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1905_root_address_inst_ack_0 <= ptr_deref_1905_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1905_resized_base_address;
      ptr_deref_1905_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1963_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1963_gather_scatter_ack_0 <= ptr_deref_1963_gather_scatter_req_0;
      aggregated_sig <= tmp22_1961;
      ptr_deref_1963_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1963_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1963_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1963_root_address_inst_ack_0 <= ptr_deref_1963_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1963_resized_base_address;
      ptr_deref_1963_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1970_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1970_gather_scatter_ack_0 <= ptr_deref_1970_gather_scatter_req_0;
      aggregated_sig <= tmp23_1968;
      ptr_deref_1970_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1970_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1970_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1970_root_address_inst_ack_0 <= ptr_deref_1970_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1970_resized_base_address;
      ptr_deref_1970_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1975_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1975_gather_scatter_ack_0 <= ptr_deref_1975_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1975_data_3 & ptr_deref_1975_data_2 & ptr_deref_1975_data_1 & ptr_deref_1975_data_0;
      tmp24_1976 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1975_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1975_root_address_inst_ack_0 <= ptr_deref_1975_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1975_resized_base_address;
      ptr_deref_1975_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_1886_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1886_resized_base_address;
      array_obj_ref_1886_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1886_root_address_inst_req_0,
          ackL => array_obj_ref_1886_root_address_inst_ack_0,
          reqR => array_obj_ref_1886_root_address_inst_req_1,
          ackR => array_obj_ref_1886_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1901_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1901_resized_base_address;
      array_obj_ref_1901_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1901_root_address_inst_req_0,
          ackL => array_obj_ref_1901_root_address_inst_ack_0,
          reqR => array_obj_ref_1901_root_address_inst_req_1,
          ackR => array_obj_ref_1901_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1847_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1838;
      tmp2_1848 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1847_inst_req_0,
          ackL => binary_1847_inst_ack_0,
          reqR => binary_1847_inst_req_1,
          ackR => binary_1847_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1865_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_1848;
      tmp5_1866 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1865_inst_req_0,
          ackL => binary_1865_inst_ack_0,
          reqR => binary_1865_inst_req_1,
          ackR => binary_1865_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_1875_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_1848;
      tmp7_1876 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1875_inst_req_0,
          ackL => binary_1875_inst_ack_0,
          reqR => binary_1875_inst_req_1,
          ackR => binary_1875_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_1914_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_1895 & tmp14_1910;
      tmp15_1915 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1914_inst_req_0,
          ackL => binary_1914_inst_ack_0,
          reqR => binary_1914_inst_req_1,
          ackR => binary_1914_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_1924_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_1915;
      tmp17_1925 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1924_inst_req_0,
          ackL => binary_1924_inst_ack_0,
          reqR => binary_1924_inst_req_1,
          ackR => binary_1924_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_1934_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_1929;
      tmp18_1935 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1934_inst_req_0,
          ackL => binary_1934_inst_ack_0,
          reqR => binary_1934_inst_req_1,
          ackR => binary_1934_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_1940_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_1915;
      tmp19_1941 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1940_inst_req_0,
          ackL => binary_1940_inst_ack_0,
          reqR => binary_1940_inst_req_1,
          ackR => binary_1940_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_1948_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1944_wire;
      notx_xx_xi_1949 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1948_inst_req_0,
          ackL => binary_1948_inst_ack_0,
          reqR => binary_1948_inst_req_1,
          ackR => binary_1948_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_1957_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_1935 & tmp20_1953;
      tmp21_1958 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1957_inst_req_0,
          ackL => binary_1957_inst_ack_0,
          reqR => binary_1957_inst_req_1,
          ackR => binary_1957_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_1858_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1858_root_address;
      ptr_deref_1858_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1858_addr_0_req_0,
          ackL => ptr_deref_1858_addr_0_ack_0,
          reqR => ptr_deref_1858_addr_0_req_1,
          ackR => ptr_deref_1858_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_1858_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1858_root_address;
      ptr_deref_1858_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1858_addr_1_req_0,
          ackL => ptr_deref_1858_addr_1_ack_0,
          reqR => ptr_deref_1858_addr_1_req_1,
          ackR => ptr_deref_1858_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_1890_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1890_root_address;
      ptr_deref_1890_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1890_addr_0_req_0,
          ackL => ptr_deref_1890_addr_0_ack_0,
          reqR => ptr_deref_1890_addr_0_req_1,
          ackR => ptr_deref_1890_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_1890_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1890_root_address;
      ptr_deref_1890_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1890_addr_1_req_0,
          ackL => ptr_deref_1890_addr_1_ack_0,
          reqR => ptr_deref_1890_addr_1_req_1,
          ackR => ptr_deref_1890_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_1890_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1890_root_address;
      ptr_deref_1890_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1890_addr_2_req_0,
          ackL => ptr_deref_1890_addr_2_ack_0,
          reqR => ptr_deref_1890_addr_2_req_1,
          ackR => ptr_deref_1890_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_1890_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1890_root_address;
      ptr_deref_1890_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1890_addr_3_req_0,
          ackL => ptr_deref_1890_addr_3_ack_0,
          reqR => ptr_deref_1890_addr_3_req_1,
          ackR => ptr_deref_1890_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_1905_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1905_root_address;
      ptr_deref_1905_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1905_addr_0_req_0,
          ackL => ptr_deref_1905_addr_0_ack_0,
          reqR => ptr_deref_1905_addr_0_req_1,
          ackR => ptr_deref_1905_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_1905_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1905_root_address;
      ptr_deref_1905_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1905_addr_1_req_0,
          ackL => ptr_deref_1905_addr_1_ack_0,
          reqR => ptr_deref_1905_addr_1_req_1,
          ackR => ptr_deref_1905_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_1905_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1905_root_address;
      ptr_deref_1905_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1905_addr_2_req_0,
          ackL => ptr_deref_1905_addr_2_ack_0,
          reqR => ptr_deref_1905_addr_2_req_1,
          ackR => ptr_deref_1905_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_1905_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1905_root_address;
      ptr_deref_1905_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1905_addr_3_req_0,
          ackL => ptr_deref_1905_addr_3_ack_0,
          reqR => ptr_deref_1905_addr_3_req_1,
          ackR => ptr_deref_1905_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_1963_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1963_root_address;
      ptr_deref_1963_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1963_addr_0_req_0,
          ackL => ptr_deref_1963_addr_0_ack_0,
          reqR => ptr_deref_1963_addr_0_req_1,
          ackR => ptr_deref_1963_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_1963_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1963_root_address;
      ptr_deref_1963_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1963_addr_1_req_0,
          ackL => ptr_deref_1963_addr_1_ack_0,
          reqR => ptr_deref_1963_addr_1_req_1,
          ackR => ptr_deref_1963_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_1970_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1970_root_address;
      ptr_deref_1970_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1970_addr_0_req_0,
          ackL => ptr_deref_1970_addr_0_ack_0,
          reqR => ptr_deref_1970_addr_0_req_1,
          ackR => ptr_deref_1970_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_1970_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1970_root_address;
      ptr_deref_1970_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1970_addr_1_req_0,
          ackL => ptr_deref_1970_addr_1_ack_0,
          reqR => ptr_deref_1970_addr_1_req_1,
          ackR => ptr_deref_1970_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_1975_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1975_root_address;
      ptr_deref_1975_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1975_addr_0_req_0,
          ackL => ptr_deref_1975_addr_0_ack_0,
          reqR => ptr_deref_1975_addr_0_req_1,
          ackR => ptr_deref_1975_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_1975_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1975_root_address;
      ptr_deref_1975_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1975_addr_1_req_0,
          ackL => ptr_deref_1975_addr_1_ack_0,
          reqR => ptr_deref_1975_addr_1_req_1,
          ackR => ptr_deref_1975_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_1975_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1975_root_address;
      ptr_deref_1975_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1975_addr_2_req_0,
          ackL => ptr_deref_1975_addr_2_ack_0,
          reqR => ptr_deref_1975_addr_2_req_1,
          ackR => ptr_deref_1975_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_1975_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1975_root_address;
      ptr_deref_1975_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1975_addr_3_req_0,
          ackL => ptr_deref_1975_addr_3_ack_0,
          reqR => ptr_deref_1975_addr_3_req_1,
          ackR => ptr_deref_1975_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_1905_load_0 ptr_deref_1975_load_0 ptr_deref_1905_load_3 ptr_deref_1905_load_1 ptr_deref_1905_load_2 ptr_deref_1975_load_3 ptr_deref_1890_load_0 ptr_deref_1890_load_1 ptr_deref_1890_load_2 ptr_deref_1890_load_3 ptr_deref_1975_load_2 ptr_deref_1975_load_1 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1905_load_0_req_0,
        ptr_deref_1905_load_0_ack_0,
        ptr_deref_1905_load_0_req_1,
        ptr_deref_1905_load_0_ack_1,
        "ptr_deref_1905_load_0",
        "memory_space_5" ,
        ptr_deref_1905_data_0,
        ptr_deref_1905_word_address_0,
        "ptr_deref_1905_data_0",
        "ptr_deref_1905_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1975_load_0_req_0,
        ptr_deref_1975_load_0_ack_0,
        ptr_deref_1975_load_0_req_1,
        ptr_deref_1975_load_0_ack_1,
        "ptr_deref_1975_load_0",
        "memory_space_5" ,
        ptr_deref_1975_data_0,
        ptr_deref_1975_word_address_0,
        "ptr_deref_1975_data_0",
        "ptr_deref_1975_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1905_load_3_req_0,
        ptr_deref_1905_load_3_ack_0,
        ptr_deref_1905_load_3_req_1,
        ptr_deref_1905_load_3_ack_1,
        "ptr_deref_1905_load_3",
        "memory_space_5" ,
        ptr_deref_1905_data_3,
        ptr_deref_1905_word_address_3,
        "ptr_deref_1905_data_3",
        "ptr_deref_1905_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1905_load_1_req_0,
        ptr_deref_1905_load_1_ack_0,
        ptr_deref_1905_load_1_req_1,
        ptr_deref_1905_load_1_ack_1,
        "ptr_deref_1905_load_1",
        "memory_space_5" ,
        ptr_deref_1905_data_1,
        ptr_deref_1905_word_address_1,
        "ptr_deref_1905_data_1",
        "ptr_deref_1905_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1905_load_2_req_0,
        ptr_deref_1905_load_2_ack_0,
        ptr_deref_1905_load_2_req_1,
        ptr_deref_1905_load_2_ack_1,
        "ptr_deref_1905_load_2",
        "memory_space_5" ,
        ptr_deref_1905_data_2,
        ptr_deref_1905_word_address_2,
        "ptr_deref_1905_data_2",
        "ptr_deref_1905_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1975_load_3_req_0,
        ptr_deref_1975_load_3_ack_0,
        ptr_deref_1975_load_3_req_1,
        ptr_deref_1975_load_3_ack_1,
        "ptr_deref_1975_load_3",
        "memory_space_5" ,
        ptr_deref_1975_data_3,
        ptr_deref_1975_word_address_3,
        "ptr_deref_1975_data_3",
        "ptr_deref_1975_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1890_load_0_req_0,
        ptr_deref_1890_load_0_ack_0,
        ptr_deref_1890_load_0_req_1,
        ptr_deref_1890_load_0_ack_1,
        "ptr_deref_1890_load_0",
        "memory_space_5" ,
        ptr_deref_1890_data_0,
        ptr_deref_1890_word_address_0,
        "ptr_deref_1890_data_0",
        "ptr_deref_1890_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1890_load_1_req_0,
        ptr_deref_1890_load_1_ack_0,
        ptr_deref_1890_load_1_req_1,
        ptr_deref_1890_load_1_ack_1,
        "ptr_deref_1890_load_1",
        "memory_space_5" ,
        ptr_deref_1890_data_1,
        ptr_deref_1890_word_address_1,
        "ptr_deref_1890_data_1",
        "ptr_deref_1890_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1890_load_2_req_0,
        ptr_deref_1890_load_2_ack_0,
        ptr_deref_1890_load_2_req_1,
        ptr_deref_1890_load_2_ack_1,
        "ptr_deref_1890_load_2",
        "memory_space_5" ,
        ptr_deref_1890_data_2,
        ptr_deref_1890_word_address_2,
        "ptr_deref_1890_data_2",
        "ptr_deref_1890_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1890_load_3_req_0,
        ptr_deref_1890_load_3_ack_0,
        ptr_deref_1890_load_3_req_1,
        ptr_deref_1890_load_3_ack_1,
        "ptr_deref_1890_load_3",
        "memory_space_5" ,
        ptr_deref_1890_data_3,
        ptr_deref_1890_word_address_3,
        "ptr_deref_1890_data_3",
        "ptr_deref_1890_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1975_load_2_req_0,
        ptr_deref_1975_load_2_ack_0,
        ptr_deref_1975_load_2_req_1,
        ptr_deref_1975_load_2_ack_1,
        "ptr_deref_1975_load_2",
        "memory_space_5" ,
        ptr_deref_1975_data_2,
        ptr_deref_1975_word_address_2,
        "ptr_deref_1975_data_2",
        "ptr_deref_1975_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1975_load_1_req_0,
        ptr_deref_1975_load_1_ack_0,
        ptr_deref_1975_load_1_req_1,
        ptr_deref_1975_load_1_ack_1,
        "ptr_deref_1975_load_1",
        "memory_space_5" ,
        ptr_deref_1975_data_1,
        ptr_deref_1975_word_address_1,
        "ptr_deref_1975_data_1",
        "ptr_deref_1975_word_address_1" -- 
      );
      reqL(11) <= ptr_deref_1905_load_0_req_0;
      reqL(10) <= ptr_deref_1975_load_0_req_0;
      reqL(9) <= ptr_deref_1905_load_3_req_0;
      reqL(8) <= ptr_deref_1905_load_1_req_0;
      reqL(7) <= ptr_deref_1905_load_2_req_0;
      reqL(6) <= ptr_deref_1975_load_3_req_0;
      reqL(5) <= ptr_deref_1890_load_0_req_0;
      reqL(4) <= ptr_deref_1890_load_1_req_0;
      reqL(3) <= ptr_deref_1890_load_2_req_0;
      reqL(2) <= ptr_deref_1890_load_3_req_0;
      reqL(1) <= ptr_deref_1975_load_2_req_0;
      reqL(0) <= ptr_deref_1975_load_1_req_0;
      ptr_deref_1905_load_0_ack_0 <= ackL(11);
      ptr_deref_1975_load_0_ack_0 <= ackL(10);
      ptr_deref_1905_load_3_ack_0 <= ackL(9);
      ptr_deref_1905_load_1_ack_0 <= ackL(8);
      ptr_deref_1905_load_2_ack_0 <= ackL(7);
      ptr_deref_1975_load_3_ack_0 <= ackL(6);
      ptr_deref_1890_load_0_ack_0 <= ackL(5);
      ptr_deref_1890_load_1_ack_0 <= ackL(4);
      ptr_deref_1890_load_2_ack_0 <= ackL(3);
      ptr_deref_1890_load_3_ack_0 <= ackL(2);
      ptr_deref_1975_load_2_ack_0 <= ackL(1);
      ptr_deref_1975_load_1_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_1905_load_0_req_1;
      reqR(10) <= ptr_deref_1975_load_0_req_1;
      reqR(9) <= ptr_deref_1905_load_3_req_1;
      reqR(8) <= ptr_deref_1905_load_1_req_1;
      reqR(7) <= ptr_deref_1905_load_2_req_1;
      reqR(6) <= ptr_deref_1975_load_3_req_1;
      reqR(5) <= ptr_deref_1890_load_0_req_1;
      reqR(4) <= ptr_deref_1890_load_1_req_1;
      reqR(3) <= ptr_deref_1890_load_2_req_1;
      reqR(2) <= ptr_deref_1890_load_3_req_1;
      reqR(1) <= ptr_deref_1975_load_2_req_1;
      reqR(0) <= ptr_deref_1975_load_1_req_1;
      ptr_deref_1905_load_0_ack_1 <= ackR(11);
      ptr_deref_1975_load_0_ack_1 <= ackR(10);
      ptr_deref_1905_load_3_ack_1 <= ackR(9);
      ptr_deref_1905_load_1_ack_1 <= ackR(8);
      ptr_deref_1905_load_2_ack_1 <= ackR(7);
      ptr_deref_1975_load_3_ack_1 <= ackR(6);
      ptr_deref_1890_load_0_ack_1 <= ackR(5);
      ptr_deref_1890_load_1_ack_1 <= ackR(4);
      ptr_deref_1890_load_2_ack_1 <= ackR(3);
      ptr_deref_1890_load_3_ack_1 <= ackR(2);
      ptr_deref_1975_load_2_ack_1 <= ackR(1);
      ptr_deref_1975_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_1905_word_address_0 & ptr_deref_1975_word_address_0 & ptr_deref_1905_word_address_3 & ptr_deref_1905_word_address_1 & ptr_deref_1905_word_address_2 & ptr_deref_1975_word_address_3 & ptr_deref_1890_word_address_0 & ptr_deref_1890_word_address_1 & ptr_deref_1890_word_address_2 & ptr_deref_1890_word_address_3 & ptr_deref_1975_word_address_2 & ptr_deref_1975_word_address_1;
      ptr_deref_1905_data_0 <= data_out(95 downto 88);
      ptr_deref_1975_data_0 <= data_out(87 downto 80);
      ptr_deref_1905_data_3 <= data_out(79 downto 72);
      ptr_deref_1905_data_1 <= data_out(71 downto 64);
      ptr_deref_1905_data_2 <= data_out(63 downto 56);
      ptr_deref_1975_data_3 <= data_out(55 downto 48);
      ptr_deref_1890_data_0 <= data_out(47 downto 40);
      ptr_deref_1890_data_1 <= data_out(39 downto 32);
      ptr_deref_1890_data_2 <= data_out(31 downto 24);
      ptr_deref_1890_data_3 <= data_out(23 downto 16);
      ptr_deref_1975_data_2 <= data_out(15 downto 8);
      ptr_deref_1975_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_1963_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1963_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1963_word_address_1) &  " data ptr_deref_1963_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1963_data_1) severity note; --
        end if;
        if ptr_deref_1858_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1858_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1858_word_address_0) &  " data ptr_deref_1858_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1858_data_0) severity note; --
        end if;
        if ptr_deref_1963_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1963_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1963_word_address_0) &  " data ptr_deref_1963_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1963_data_0) severity note; --
        end if;
        if ptr_deref_1970_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1970_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1970_word_address_1) &  " data ptr_deref_1970_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1970_data_1) severity note; --
        end if;
        if ptr_deref_1970_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1970_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1970_word_address_0) &  " data ptr_deref_1970_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1970_data_0) severity note; --
        end if;
        if ptr_deref_1858_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1858_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1858_word_address_1) &  " data ptr_deref_1858_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1858_data_1) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1963_store_1 ptr_deref_1858_store_0 ptr_deref_1963_store_0 ptr_deref_1970_store_1 ptr_deref_1970_store_0 ptr_deref_1858_store_1 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_1963_store_1_req_0;
      reqL(4) <= ptr_deref_1858_store_0_req_0;
      reqL(3) <= ptr_deref_1963_store_0_req_0;
      reqL(2) <= ptr_deref_1970_store_1_req_0;
      reqL(1) <= ptr_deref_1970_store_0_req_0;
      reqL(0) <= ptr_deref_1858_store_1_req_0;
      ptr_deref_1963_store_1_ack_0 <= ackL(5);
      ptr_deref_1858_store_0_ack_0 <= ackL(4);
      ptr_deref_1963_store_0_ack_0 <= ackL(3);
      ptr_deref_1970_store_1_ack_0 <= ackL(2);
      ptr_deref_1970_store_0_ack_0 <= ackL(1);
      ptr_deref_1858_store_1_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_1963_store_1_req_1;
      reqR(4) <= ptr_deref_1858_store_0_req_1;
      reqR(3) <= ptr_deref_1963_store_0_req_1;
      reqR(2) <= ptr_deref_1970_store_1_req_1;
      reqR(1) <= ptr_deref_1970_store_0_req_1;
      reqR(0) <= ptr_deref_1858_store_1_req_1;
      ptr_deref_1963_store_1_ack_1 <= ackR(5);
      ptr_deref_1858_store_0_ack_1 <= ackR(4);
      ptr_deref_1963_store_0_ack_1 <= ackR(3);
      ptr_deref_1970_store_1_ack_1 <= ackR(2);
      ptr_deref_1970_store_0_ack_1 <= ackR(1);
      ptr_deref_1858_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1963_word_address_1 & ptr_deref_1858_word_address_0 & ptr_deref_1963_word_address_0 & ptr_deref_1970_word_address_1 & ptr_deref_1970_word_address_0 & ptr_deref_1858_word_address_1;
      data_in <= ptr_deref_1963_data_1 & ptr_deref_1858_data_0 & ptr_deref_1963_data_0 & ptr_deref_1970_data_1 & ptr_deref_1970_data_0 & ptr_deref_1858_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_1836_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_1836_inst_ack_0 then -- 
            assert false report " ReadPipe to0_in0 to wire simple_obj_ref_1836_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_1836_inst_req_0;
      simple_obj_ref_1836_inst_ack_0 <= ack(0);
      simple_obj_ref_1836_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to0_in0_pipe_read_req(0),
          oack => to0_in0_pipe_read_ack(0),
          odata => to0_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1981_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_1983_wire_constant value="  &  convert_slv_to_hex_string(type_cast_1983_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_1981_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1981_inst_req_0;
      simple_obj_ref_1981_inst_ack_0 <= ack(0);
      data_in <= type_cast_1983_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1985_inst_ack_0 then -- 
          assert false report " WritePipe tofpga0_out0 from wire type_cast_1987_wire value="  &  convert_slv_to_hex_string(type_cast_1987_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_1985_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1985_inst_req_0;
      simple_obj_ref_1985_inst_ack_0 <= ack(0);
      data_in <= type_cast_1987_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga0_out0_pipe_write_req(0),
          oack => tofpga0_out0_pipe_write_ack(0),
          odata => tofpga0_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1968_call call_stmt_1961_call call_stmt_1856_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_1968_call_req_0;
      reqL(1) <= call_stmt_1961_call_req_0;
      reqL(0) <= call_stmt_1856_call_req_0;
      call_stmt_1968_call_ack_0 <= ackL(2);
      call_stmt_1961_call_ack_0 <= ackL(1);
      call_stmt_1856_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_1968_call_req_1;
      reqR(1) <= call_stmt_1961_call_req_1;
      reqR(0) <= call_stmt_1856_call_req_1;
      call_stmt_1968_call_ack_1 <= ackR(2);
      call_stmt_1961_call_ack_1 <= ackR(1);
      call_stmt_1856_call_ack_1 <= ackR(0);
      data_in <= tmp21_1958 & tmp16_1919 & type_cast_1854_wire_constant;
      tmp23_1968 <= data_out(47 downto 32);
      tmp22_1961 <= data_out(31 downto 16);
      tmp4_1856 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to1_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to1_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to1_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga1_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to1;
architecture Default of ahir_glue_to1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to1_CP_9606_start: Boolean;
  -- links between control-path and data-path
  signal binary_2007_inst_ack_0 : boolean;
  signal array_obj_ref_2046_final_reg_ack_0 : boolean;
  signal type_cast_2054_inst_ack_0 : boolean;
  signal type_cast_2039_inst_req_0 : boolean;
  signal ptr_deref_2018_gather_scatter_ack_0 : boolean;
  signal call_stmt_2016_call_ack_0 : boolean;
  signal type_cast_2029_inst_ack_0 : boolean;
  signal binary_2007_inst_ack_1 : boolean;
  signal array_obj_ref_2061_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2050_addr_3_req_0 : boolean;
  signal type_cast_2029_inst_req_0 : boolean;
  signal ptr_deref_2018_base_resize_req_0 : boolean;
  signal ptr_deref_2050_load_2_req_0 : boolean;
  signal array_obj_ref_2046_final_reg_req_0 : boolean;
  signal ptr_deref_2018_addr_1_ack_1 : boolean;
  signal ptr_deref_2065_addr_0_ack_0 : boolean;
  signal ptr_deref_2065_base_resize_ack_0 : boolean;
  signal ptr_deref_2018_gather_scatter_req_0 : boolean;
  signal ptr_deref_2065_addr_1_ack_1 : boolean;
  signal ptr_deref_2065_load_1_ack_1 : boolean;
  signal call_stmt_2016_call_req_0 : boolean;
  signal ptr_deref_2065_load_1_req_0 : boolean;
  signal array_obj_ref_2046_root_address_inst_req_0 : boolean;
  signal ptr_deref_2018_addr_1_req_1 : boolean;
  signal ptr_deref_2018_store_1_req_0 : boolean;
  signal ptr_deref_2018_addr_1_ack_0 : boolean;
  signal binary_2025_inst_req_1 : boolean;
  signal simple_obj_ref_1996_inst_req_0 : boolean;
  signal binary_2025_inst_ack_1 : boolean;
  signal binary_2025_inst_req_0 : boolean;
  signal ptr_deref_2065_addr_3_req_1 : boolean;
  signal ptr_deref_2018_root_address_inst_ack_0 : boolean;
  signal type_cast_2054_inst_req_0 : boolean;
  signal ptr_deref_2018_addr_0_ack_1 : boolean;
  signal ptr_deref_2050_load_2_ack_0 : boolean;
  signal binary_2025_inst_ack_0 : boolean;
  signal ptr_deref_2065_load_2_req_1 : boolean;
  signal ptr_deref_2018_store_1_req_1 : boolean;
  signal type_cast_2011_inst_ack_0 : boolean;
  signal ptr_deref_2050_load_1_req_0 : boolean;
  signal ptr_deref_2018_store_0_ack_1 : boolean;
  signal type_cast_1997_inst_ack_0 : boolean;
  signal ptr_deref_2065_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2018_root_address_inst_req_0 : boolean;
  signal ptr_deref_2065_load_3_ack_0 : boolean;
  signal ptr_deref_2050_addr_0_req_1 : boolean;
  signal type_cast_2001_inst_ack_0 : boolean;
  signal ptr_deref_2065_load_0_req_0 : boolean;
  signal array_obj_ref_2061_final_reg_req_0 : boolean;
  signal ptr_deref_2065_addr_1_req_0 : boolean;
  signal ptr_deref_2050_addr_2_req_0 : boolean;
  signal binary_2084_inst_req_0 : boolean;
  signal ptr_deref_2065_gather_scatter_req_0 : boolean;
  signal ptr_deref_2065_load_2_ack_0 : boolean;
  signal ptr_deref_2050_addr_3_ack_0 : boolean;
  signal ptr_deref_2065_addr_1_req_1 : boolean;
  signal array_obj_ref_2046_base_resize_req_0 : boolean;
  signal ptr_deref_2018_store_0_req_1 : boolean;
  signal array_obj_ref_2046_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2018_base_resize_ack_0 : boolean;
  signal ptr_deref_2018_addr_0_req_1 : boolean;
  signal type_cast_1997_inst_req_0 : boolean;
  signal ptr_deref_2065_load_0_ack_0 : boolean;
  signal ptr_deref_2018_addr_1_req_0 : boolean;
  signal binary_2074_inst_req_1 : boolean;
  signal ptr_deref_2050_addr_1_req_0 : boolean;
  signal binary_2007_inst_req_1 : boolean;
  signal ptr_deref_2018_store_0_req_0 : boolean;
  signal ptr_deref_2065_addr_2_req_0 : boolean;
  signal ptr_deref_2065_load_2_ack_1 : boolean;
  signal type_cast_2039_inst_ack_0 : boolean;
  signal ptr_deref_2018_store_0_ack_0 : boolean;
  signal type_cast_2011_inst_req_0 : boolean;
  signal ptr_deref_2050_load_1_ack_0 : boolean;
  signal ptr_deref_2065_load_3_req_0 : boolean;
  signal array_obj_ref_2046_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2050_addr_3_ack_1 : boolean;
  signal binary_2108_inst_ack_1 : boolean;
  signal ptr_deref_2065_load_1_req_1 : boolean;
  signal binary_2100_inst_req_1 : boolean;
  signal ptr_deref_2018_addr_0_ack_0 : boolean;
  signal binary_2084_inst_ack_0 : boolean;
  signal ptr_deref_2065_base_resize_req_0 : boolean;
  signal binary_2074_inst_ack_1 : boolean;
  signal ptr_deref_2065_addr_3_ack_0 : boolean;
  signal array_obj_ref_2046_root_address_inst_req_1 : boolean;
  signal binary_2100_inst_ack_0 : boolean;
  signal binary_2074_inst_ack_0 : boolean;
  signal ptr_deref_2050_load_0_req_0 : boolean;
  signal type_cast_2088_inst_req_0 : boolean;
  signal ptr_deref_2065_load_0_req_1 : boolean;
  signal ptr_deref_2065_load_3_ack_1 : boolean;
  signal type_cast_2078_inst_ack_0 : boolean;
  signal ptr_deref_2065_load_0_ack_1 : boolean;
  signal ptr_deref_2018_addr_0_req_0 : boolean;
  signal ptr_deref_2018_store_1_ack_1 : boolean;
  signal binary_2094_inst_req_1 : boolean;
  signal ptr_deref_2065_addr_0_req_0 : boolean;
  signal ptr_deref_2050_addr_0_ack_1 : boolean;
  signal ptr_deref_2050_load_0_ack_0 : boolean;
  signal binary_2117_inst_req_0 : boolean;
  signal array_obj_ref_2046_base_resize_ack_0 : boolean;
  signal ptr_deref_2065_load_3_req_1 : boolean;
  signal ptr_deref_2050_addr_0_ack_0 : boolean;
  signal ptr_deref_2065_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2050_addr_3_req_1 : boolean;
  signal binary_2108_inst_req_1 : boolean;
  signal binary_2007_inst_req_0 : boolean;
  signal simple_obj_ref_1996_inst_ack_0 : boolean;
  signal binary_2117_inst_ack_0 : boolean;
  signal binary_2117_inst_req_1 : boolean;
  signal binary_2117_inst_ack_1 : boolean;
  signal type_cast_2104_inst_req_0 : boolean;
  signal binary_2108_inst_req_0 : boolean;
  signal binary_2108_inst_ack_0 : boolean;
  signal type_cast_2112_inst_req_0 : boolean;
  signal type_cast_2104_inst_ack_0 : boolean;
  signal ptr_deref_2050_addr_0_req_0 : boolean;
  signal ptr_deref_2050_addr_2_ack_0 : boolean;
  signal ptr_deref_2050_load_3_req_0 : boolean;
  signal ptr_deref_2050_load_3_ack_0 : boolean;
  signal ptr_deref_2065_load_1_ack_0 : boolean;
  signal array_obj_ref_2061_final_reg_ack_0 : boolean;
  signal binary_2035_inst_req_0 : boolean;
  signal array_obj_ref_2061_base_resize_req_0 : boolean;
  signal array_obj_ref_2061_base_resize_ack_0 : boolean;
  signal ptr_deref_2065_addr_2_ack_0 : boolean;
  signal type_cast_2069_inst_req_0 : boolean;
  signal ptr_deref_2050_addr_1_ack_0 : boolean;
  signal binary_2035_inst_req_1 : boolean;
  signal type_cast_2069_inst_ack_0 : boolean;
  signal binary_2035_inst_ack_0 : boolean;
  signal ptr_deref_2065_addr_3_ack_1 : boolean;
  signal ptr_deref_2050_base_resize_req_0 : boolean;
  signal ptr_deref_2018_store_1_ack_0 : boolean;
  signal binary_2035_inst_ack_1 : boolean;
  signal ptr_deref_2050_addr_2_req_1 : boolean;
  signal call_stmt_2016_call_req_1 : boolean;
  signal ptr_deref_2050_base_resize_ack_0 : boolean;
  signal ptr_deref_2065_load_2_req_0 : boolean;
  signal ptr_deref_2065_addr_1_ack_0 : boolean;
  signal ptr_deref_2050_load_0_req_1 : boolean;
  signal ptr_deref_2050_load_0_ack_1 : boolean;
  signal call_stmt_2016_call_ack_1 : boolean;
  signal ptr_deref_2050_addr_1_req_1 : boolean;
  signal ptr_deref_2050_addr_2_ack_1 : boolean;
  signal array_obj_ref_2061_root_address_inst_req_0 : boolean;
  signal ptr_deref_2050_load_1_req_1 : boolean;
  signal ptr_deref_2050_load_1_ack_1 : boolean;
  signal type_cast_2001_inst_req_0 : boolean;
  signal ptr_deref_2050_root_address_inst_req_0 : boolean;
  signal ptr_deref_2050_root_address_inst_ack_0 : boolean;
  signal binary_2094_inst_req_0 : boolean;
  signal binary_2084_inst_req_1 : boolean;
  signal ptr_deref_2050_load_2_req_1 : boolean;
  signal array_obj_ref_2061_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2050_load_2_ack_1 : boolean;
  signal binary_2074_inst_req_0 : boolean;
  signal type_cast_2088_inst_ack_0 : boolean;
  signal type_cast_2078_inst_req_0 : boolean;
  signal ptr_deref_2050_addr_1_ack_1 : boolean;
  signal binary_2100_inst_req_0 : boolean;
  signal ptr_deref_2065_addr_0_req_1 : boolean;
  signal ptr_deref_2050_load_3_req_1 : boolean;
  signal binary_2084_inst_ack_1 : boolean;
  signal ptr_deref_2050_load_3_ack_1 : boolean;
  signal ptr_deref_2050_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2061_root_address_inst_req_1 : boolean;
  signal binary_2094_inst_ack_0 : boolean;
  signal binary_2094_inst_ack_1 : boolean;
  signal ptr_deref_2065_addr_0_ack_1 : boolean;
  signal binary_2100_inst_ack_1 : boolean;
  signal ptr_deref_2050_gather_scatter_ack_0 : boolean;
  signal type_cast_2112_inst_ack_0 : boolean;
  signal ptr_deref_2123_base_resize_req_0 : boolean;
  signal ptr_deref_2123_base_resize_ack_0 : boolean;
  signal ptr_deref_2123_gather_scatter_req_0 : boolean;
  signal ptr_deref_2123_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2123_store_0_req_0 : boolean;
  signal ptr_deref_2123_addr_0_req_1 : boolean;
  signal ptr_deref_2123_addr_0_ack_1 : boolean;
  signal ptr_deref_2123_addr_1_req_0 : boolean;
  signal ptr_deref_2123_addr_1_ack_0 : boolean;
  signal call_stmt_2121_call_req_1 : boolean;
  signal call_stmt_2121_call_ack_1 : boolean;
  signal call_stmt_2128_call_req_0 : boolean;
  signal call_stmt_2128_call_ack_0 : boolean;
  signal ptr_deref_2123_store_0_ack_0 : boolean;
  signal ptr_deref_2123_store_1_req_0 : boolean;
  signal ptr_deref_2123_store_1_ack_0 : boolean;
  signal ptr_deref_2123_addr_0_req_0 : boolean;
  signal ptr_deref_2123_addr_0_ack_0 : boolean;
  signal ptr_deref_2123_root_address_inst_req_0 : boolean;
  signal ptr_deref_2123_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2123_addr_1_req_1 : boolean;
  signal ptr_deref_2123_addr_1_ack_1 : boolean;
  signal call_stmt_2128_call_req_1 : boolean;
  signal call_stmt_2128_call_ack_1 : boolean;
  signal ptr_deref_2123_store_1_req_1 : boolean;
  signal ptr_deref_2123_store_1_ack_1 : boolean;
  signal ptr_deref_2123_store_0_req_1 : boolean;
  signal ptr_deref_2123_store_0_ack_1 : boolean;
  signal call_stmt_2121_call_req_0 : boolean;
  signal call_stmt_2121_call_ack_0 : boolean;
  signal ptr_deref_2065_root_address_inst_req_0 : boolean;
  signal ptr_deref_2065_addr_3_req_0 : boolean;
  signal ptr_deref_2065_addr_2_ack_1 : boolean;
  signal ptr_deref_2065_addr_2_req_1 : boolean;
  signal ptr_deref_2130_base_resize_req_0 : boolean;
  signal ptr_deref_2130_base_resize_ack_0 : boolean;
  signal ptr_deref_2130_root_address_inst_req_0 : boolean;
  signal ptr_deref_2130_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2130_addr_0_req_0 : boolean;
  signal ptr_deref_2130_addr_0_ack_0 : boolean;
  signal ptr_deref_2130_addr_0_req_1 : boolean;
  signal ptr_deref_2130_addr_0_ack_1 : boolean;
  signal ptr_deref_2130_addr_1_req_0 : boolean;
  signal ptr_deref_2130_addr_1_ack_0 : boolean;
  signal ptr_deref_2130_addr_1_req_1 : boolean;
  signal ptr_deref_2130_addr_1_ack_1 : boolean;
  signal ptr_deref_2130_gather_scatter_req_0 : boolean;
  signal ptr_deref_2130_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2130_store_0_req_0 : boolean;
  signal ptr_deref_2130_store_0_ack_0 : boolean;
  signal ptr_deref_2130_store_1_req_0 : boolean;
  signal ptr_deref_2130_store_1_ack_0 : boolean;
  signal ptr_deref_2130_store_0_req_1 : boolean;
  signal ptr_deref_2130_store_0_ack_1 : boolean;
  signal ptr_deref_2130_store_1_req_1 : boolean;
  signal ptr_deref_2130_store_1_ack_1 : boolean;
  signal ptr_deref_2135_base_resize_req_0 : boolean;
  signal ptr_deref_2135_base_resize_ack_0 : boolean;
  signal ptr_deref_2135_root_address_inst_req_0 : boolean;
  signal ptr_deref_2135_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2135_addr_0_req_0 : boolean;
  signal ptr_deref_2135_addr_0_ack_0 : boolean;
  signal ptr_deref_2135_addr_0_req_1 : boolean;
  signal ptr_deref_2135_addr_0_ack_1 : boolean;
  signal ptr_deref_2135_addr_1_req_0 : boolean;
  signal ptr_deref_2135_addr_1_ack_0 : boolean;
  signal ptr_deref_2135_addr_1_req_1 : boolean;
  signal ptr_deref_2135_addr_1_ack_1 : boolean;
  signal ptr_deref_2135_addr_2_req_0 : boolean;
  signal ptr_deref_2135_addr_2_ack_0 : boolean;
  signal ptr_deref_2135_addr_2_req_1 : boolean;
  signal ptr_deref_2135_addr_2_ack_1 : boolean;
  signal ptr_deref_2135_addr_3_req_0 : boolean;
  signal ptr_deref_2135_addr_3_ack_0 : boolean;
  signal ptr_deref_2135_addr_3_req_1 : boolean;
  signal ptr_deref_2135_addr_3_ack_1 : boolean;
  signal ptr_deref_2135_load_0_req_0 : boolean;
  signal ptr_deref_2135_load_0_ack_0 : boolean;
  signal ptr_deref_2135_load_1_req_0 : boolean;
  signal ptr_deref_2135_load_1_ack_0 : boolean;
  signal ptr_deref_2135_load_2_req_0 : boolean;
  signal ptr_deref_2135_load_2_ack_0 : boolean;
  signal ptr_deref_2135_load_3_req_0 : boolean;
  signal ptr_deref_2135_load_3_ack_0 : boolean;
  signal ptr_deref_2135_load_0_req_1 : boolean;
  signal ptr_deref_2135_load_0_ack_1 : boolean;
  signal ptr_deref_2135_load_1_req_1 : boolean;
  signal ptr_deref_2135_load_1_ack_1 : boolean;
  signal ptr_deref_2135_load_2_req_1 : boolean;
  signal ptr_deref_2135_load_2_ack_1 : boolean;
  signal ptr_deref_2135_load_3_req_1 : boolean;
  signal ptr_deref_2135_load_3_ack_1 : boolean;
  signal ptr_deref_2135_gather_scatter_req_0 : boolean;
  signal ptr_deref_2135_gather_scatter_ack_0 : boolean;
  signal type_cast_2139_inst_req_0 : boolean;
  signal type_cast_2139_inst_ack_0 : boolean;
  signal simple_obj_ref_2141_inst_req_0 : boolean;
  signal simple_obj_ref_2141_inst_ack_0 : boolean;
  signal type_cast_2147_inst_req_0 : boolean;
  signal type_cast_2147_inst_ack_0 : boolean;
  signal simple_obj_ref_2145_inst_req_0 : boolean;
  signal simple_obj_ref_2145_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to1_CP_9606: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_9697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2016_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_10222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2121_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_10520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2141_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9652_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_1997_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_9647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_1996_inst_req_0); -- 
    ack_9648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1996_inst_ack_0, ack => cp_elements(8)); -- 
    ack_9653_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1997_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2001_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_9666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9675_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2007_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_9676_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2007_inst_ack_0, ack => cp_elements(18)); -- 
    cr_9677_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2007_inst_req_1); -- 
    ca_9678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2007_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2011_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_9688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2011_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_9698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2016_call_ack_0, ack => cp_elements(24)); -- 
    ccr_9702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2016_call_req_1); -- 
    cca_9703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2016_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_9749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2018_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_9722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2018_base_resize_req_0); -- 
    base_resize_ack_9723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_9727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2018_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2018_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_9735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2018_addr_0_req_0); -- 
    ra_9736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_9737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2018_addr_0_req_1); -- 
    ca_9738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_9742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2018_addr_1_req_0); -- 
    ra_9743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_9744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2018_addr_1_req_1); -- 
    ca_9745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2018_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_9757_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2018_store_0_req_0); -- 
    ra_9758_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_9762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2018_store_1_req_0); -- 
    ra_9763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_9773_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2018_store_0_req_1); -- 
    ca_9774_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_9778_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2018_store_1_req_1); -- 
    ca_9779_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2025_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_9789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2025_inst_ack_0, ack => cp_elements(55)); -- 
    cr_9790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2025_inst_req_1); -- 
    ca_9791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2025_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2029_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_9801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2029_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2035_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_9811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2035_inst_ack_0, ack => cp_elements(63)); -- 
    cr_9812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2035_inst_req_1); -- 
    ca_9813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2035_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2039_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_9823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2039_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_9847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2046_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_9834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2046_base_resize_req_0); -- 
    base_resize_ack_9835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2046_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_9840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2046_root_address_inst_req_0); -- 
    plus_base_ra_9841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2046_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_9842_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2046_root_address_inst_req_1); -- 
    plus_base_ca_9843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2046_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2046_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_9861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2050_base_resize_req_0); -- 
    base_resize_ack_9862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_9866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2050_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2050_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_9874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2050_addr_0_req_0); -- 
    ra_9875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_9876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2050_addr_0_req_1); -- 
    ca_9877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_9881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2050_addr_1_req_0); -- 
    ra_9882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_9883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2050_addr_1_req_1); -- 
    ca_9884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_9888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2050_addr_2_req_0); -- 
    ra_9889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_9890_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2050_addr_2_req_1); -- 
    ca_9891_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_9895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2050_addr_3_req_0); -- 
    ra_9896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_9897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2050_addr_3_req_1); -- 
    ca_9898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_9908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2050_load_0_req_0); -- 
    ra_9909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_9913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2050_load_1_req_0); -- 
    ra_9914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_9918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2050_load_2_req_0); -- 
    ra_9919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_9923_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2050_load_3_req_0); -- 
    ra_9924_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_9934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2050_load_0_req_1); -- 
    ca_9935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_9939_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2050_load_1_req_1); -- 
    ca_9940_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_9944_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2050_load_2_req_1); -- 
    ca_9945_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_9949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2050_load_3_req_1); -- 
    ca_9950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2050_gather_scatter_req_0); -- 
    merge_ack_9952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2050_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_9961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2054_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_9962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2054_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_9986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2061_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_9973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2061_base_resize_req_0); -- 
    base_resize_ack_9974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2061_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_9979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2061_root_address_inst_req_0); -- 
    plus_base_ra_9980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2061_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_9981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2061_root_address_inst_req_1); -- 
    plus_base_ca_9982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2061_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2061_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_10000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2065_base_resize_req_0); -- 
    base_resize_ack_10001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_10005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2065_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2065_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_10013_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2065_addr_0_req_0); -- 
    ra_10014_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_10015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2065_addr_0_req_1); -- 
    ca_10016_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_10020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2065_addr_1_req_0); -- 
    ra_10021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_10022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2065_addr_1_req_1); -- 
    ca_10023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_10027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2065_addr_2_req_0); -- 
    ra_10028_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_10029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2065_addr_2_req_1); -- 
    ca_10030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_10034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2065_addr_3_req_0); -- 
    ra_10035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_10036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2065_addr_3_req_1); -- 
    ca_10037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_10047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2065_load_0_req_0); -- 
    ra_10048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_10052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2065_load_1_req_0); -- 
    ra_10053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_10057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2065_load_2_req_0); -- 
    ra_10058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_10062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2065_load_3_req_0); -- 
    ra_10063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_10073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2065_load_0_req_1); -- 
    ca_10074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_10078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2065_load_1_req_1); -- 
    ca_10079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_10083_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2065_load_2_req_1); -- 
    ca_10084_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_10088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2065_load_3_req_1); -- 
    ca_10089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_10090_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2065_gather_scatter_req_0); -- 
    merge_ack_10091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2065_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2069_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_10101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2069_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_2074_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_10112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2074_inst_ack_0, ack => cp_elements(162)); -- 
    cr_10113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_2074_inst_req_1); -- 
    cp_elements(163) <= binary_2074_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_2078_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_10124_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2078_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10133_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_2084_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_10134_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2084_inst_ack_0, ack => cp_elements(171)); -- 
    cr_10135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_2084_inst_req_1); -- 
    ca_10136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2084_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_2088_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_10146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2088_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2094_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_10156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2094_inst_ack_0, ack => cp_elements(178)); -- 
    cr_10157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_2094_inst_req_1); -- 
    ca_10158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2094_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_2100_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_10168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2100_inst_ack_0, ack => cp_elements(183)); -- 
    cr_10169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2100_inst_req_1); -- 
    ca_10170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2100_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_2108_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_2104_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_10182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_0, ack => cp_elements(189)); -- 
    ra_10187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2108_inst_ack_0, ack => cp_elements(190)); -- 
    cr_10188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_2108_inst_req_1); -- 
    ca_10189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2108_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_2112_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_10199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2112_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_2117_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_10210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2117_inst_ack_0, ack => cp_elements(197)); -- 
    cr_10211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_2117_inst_req_1); -- 
    ca_10212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2117_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_10223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2121_call_ack_0, ack => cp_elements(200)); -- 
    ccr_10227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_2121_call_req_1); -- 
    cca_10228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2121_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_10274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_2123_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_10247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_2123_base_resize_req_0); -- 
    base_resize_ack_10248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_10252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2123_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_2123_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_10260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2123_addr_0_req_0); -- 
    ra_10261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_10262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_2123_addr_0_req_1); -- 
    ca_10263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_10267_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_2123_addr_1_req_0); -- 
    ra_10268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_10269_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2123_addr_1_req_1); -- 
    ca_10270_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_2123_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_10282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2123_store_0_req_0); -- 
    ra_10283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_10287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2123_store_1_req_0); -- 
    ra_10288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_10298_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_2123_store_0_req_1); -- 
    ca_10299_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_10303_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_2123_store_1_req_1); -- 
    ca_10304_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_10314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_2128_call_req_0); -- 
    cra_10315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2128_call_ack_0, ack => cp_elements(227)); -- 
    ccr_10319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_2128_call_req_1); -- 
    cca_10320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2128_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_10366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_2130_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_10339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_2130_base_resize_req_0); -- 
    base_resize_ack_10340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_10344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_2130_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_2130_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_10352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_2130_addr_0_req_0); -- 
    ra_10353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_10354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_2130_addr_0_req_1); -- 
    ca_10355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_10359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_2130_addr_1_req_0); -- 
    ra_10360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_10361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_2130_addr_1_req_1); -- 
    ca_10362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_2130_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_10374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_2130_store_0_req_0); -- 
    ra_10375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_10379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2130_store_1_req_0); -- 
    ra_10380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_10390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_2130_store_0_req_1); -- 
    ca_10391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_10395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2130_store_1_req_1); -- 
    ca_10396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2130_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_10409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_2135_base_resize_req_0); -- 
    base_resize_ack_10410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_10414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_2135_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_2135_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_10422_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_2135_addr_0_req_0); -- 
    ra_10423_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_10424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2135_addr_0_req_1); -- 
    ca_10425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_10429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2135_addr_1_req_0); -- 
    ra_10430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_10431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_2135_addr_1_req_1); -- 
    ca_10432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_10436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_2135_addr_2_req_0); -- 
    ra_10437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_10438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_2135_addr_2_req_1); -- 
    ca_10439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_10443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_2135_addr_3_req_0); -- 
    ra_10444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_10445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2135_addr_3_req_1); -- 
    ca_10446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_10456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2135_load_0_req_0); -- 
    ra_10457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_10461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_2135_load_1_req_0); -- 
    ra_10462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_10466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2135_load_2_req_0); -- 
    ra_10467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_10471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2135_load_3_req_0); -- 
    ra_10472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_10482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2135_load_0_req_1); -- 
    ca_10483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_10487_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_2135_load_1_req_1); -- 
    ca_10488_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_10492_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2135_load_2_req_1); -- 
    ca_10493_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_10497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2135_load_3_req_1); -- 
    ca_10498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_10499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_2135_gather_scatter_req_0); -- 
    merge_ack_10500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_2139_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_10510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2139_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_10521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2141_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_2147_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_10534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_10539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_2145_inst_req_0); -- 
    pipe_wack_10540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2145_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2046_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2046_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2046_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2061_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2061_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2061_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_2109 : std_logic_vector(0 downto 0);
    signal ptr_deref_2018_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2018_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2018_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2018_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2018_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2018_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2018_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2018_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2018_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2050_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2050_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2050_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2050_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2050_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2065_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2065_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2065_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2065_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2065_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2123_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2123_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2130_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2130_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2130_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2135_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2135_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2135_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2135_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1996_wire : std_logic_vector(31 downto 0);
    signal tmp10_2051 : std_logic_vector(31 downto 0);
    signal tmp11_2055 : std_logic_vector(31 downto 0);
    signal tmp12_2062 : std_logic_vector(31 downto 0);
    signal tmp13_2066 : std_logic_vector(31 downto 0);
    signal tmp14_2070 : std_logic_vector(31 downto 0);
    signal tmp15_2075 : std_logic_vector(31 downto 0);
    signal tmp16_2079 : std_logic_vector(15 downto 0);
    signal tmp17_2085 : std_logic_vector(31 downto 0);
    signal tmp18_2095 : std_logic_vector(15 downto 0);
    signal tmp19_2101 : std_logic_vector(31 downto 0);
    signal tmp1_2002 : std_logic_vector(31 downto 0);
    signal tmp20_2113 : std_logic_vector(15 downto 0);
    signal tmp21_2118 : std_logic_vector(15 downto 0);
    signal tmp22_2121 : std_logic_vector(15 downto 0);
    signal tmp23_2128 : std_logic_vector(15 downto 0);
    signal tmp24_2136 : std_logic_vector(31 downto 0);
    signal tmp25_2140 : std_logic_vector(31 downto 0);
    signal tmp2_2008 : std_logic_vector(31 downto 0);
    signal tmp3_2012 : std_logic_vector(31 downto 0);
    signal tmp4_2016 : std_logic_vector(15 downto 0);
    signal tmp5_2026 : std_logic_vector(31 downto 0);
    signal tmp6_2030 : std_logic_vector(31 downto 0);
    signal tmp7_2036 : std_logic_vector(31 downto 0);
    signal tmp8_2040 : std_logic_vector(31 downto 0);
    signal tmp9_2047 : std_logic_vector(31 downto 0);
    signal tmp_1998 : std_logic_vector(31 downto 0);
    signal type_cast_2006_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2014_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2024_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2034_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2083_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2093_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2099_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2104_wire : std_logic_vector(31 downto 0);
    signal type_cast_2107_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2143_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2147_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_2089 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2046_final_offset <= "0000000000010000";
    array_obj_ref_2061_final_offset <= "0000000000001100";
    ptr_deref_2018_word_offset_0 <= "0000000000000000";
    ptr_deref_2018_word_offset_1 <= "0000000000000001";
    ptr_deref_2050_word_offset_0 <= "0000000000000000";
    ptr_deref_2050_word_offset_1 <= "0000000000000001";
    ptr_deref_2050_word_offset_2 <= "0000000000000010";
    ptr_deref_2050_word_offset_3 <= "0000000000000011";
    ptr_deref_2065_word_offset_0 <= "0000000000000000";
    ptr_deref_2065_word_offset_1 <= "0000000000000001";
    ptr_deref_2065_word_offset_2 <= "0000000000000010";
    ptr_deref_2065_word_offset_3 <= "0000000000000011";
    ptr_deref_2123_word_offset_0 <= "0000000000000000";
    ptr_deref_2123_word_offset_1 <= "0000000000000001";
    ptr_deref_2130_word_offset_0 <= "0000000000000000";
    ptr_deref_2130_word_offset_1 <= "0000000000000001";
    ptr_deref_2135_word_offset_0 <= "0000000000000000";
    ptr_deref_2135_word_offset_1 <= "0000000000000001";
    ptr_deref_2135_word_offset_2 <= "0000000000000010";
    ptr_deref_2135_word_offset_3 <= "0000000000000011";
    type_cast_2006_wire_constant <= "11111111111111111111100000000000";
    type_cast_2014_wire_constant <= "0000000000000010";
    type_cast_2024_wire_constant <= "00000000000000000000000000000110";
    type_cast_2034_wire_constant <= "00000000000000000000000000000010";
    type_cast_2083_wire_constant <= "00000000000000000000000000000011";
    type_cast_2093_wire_constant <= "0001111111111111";
    type_cast_2099_wire_constant <= "00000000000000000000000000000111";
    type_cast_2107_wire_constant <= "00000000000000000000000000000000";
    type_cast_2143_wire_constant <= "00000000000000000000000000000010";
    array_obj_ref_2046_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2002, dout => array_obj_ref_2046_resized_base_address, req => array_obj_ref_2046_base_resize_req_0, ack => array_obj_ref_2046_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2046_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2046_root_address, dout => tmp9_2047, req => array_obj_ref_2046_final_reg_req_0, ack => array_obj_ref_2046_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2061_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2002, dout => array_obj_ref_2061_resized_base_address, req => array_obj_ref_2061_base_resize_req_0, ack => array_obj_ref_2061_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2061_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2061_root_address, dout => tmp12_2062, req => array_obj_ref_2061_final_reg_req_0, ack => array_obj_ref_2061_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2018_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2012, dout => ptr_deref_2018_resized_base_address, req => ptr_deref_2018_base_resize_req_0, ack => ptr_deref_2018_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2050_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2047, dout => ptr_deref_2050_resized_base_address, req => ptr_deref_2050_base_resize_req_0, ack => ptr_deref_2050_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2065_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2062, dout => ptr_deref_2065_resized_base_address, req => ptr_deref_2065_base_resize_req_0, ack => ptr_deref_2065_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2123_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2030, dout => ptr_deref_2123_resized_base_address, req => ptr_deref_2123_base_resize_req_0, ack => ptr_deref_2123_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2130_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2040, dout => ptr_deref_2130_resized_base_address, req => ptr_deref_2130_base_resize_req_0, ack => ptr_deref_2130_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2135_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2062, dout => ptr_deref_2135_resized_base_address, req => ptr_deref_2135_base_resize_req_0, ack => ptr_deref_2135_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1997_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_1996_wire, dout => tmp_1998, req => type_cast_1997_inst_req_0, ack => type_cast_1997_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2001_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_1998, dout => tmp1_2002, req => type_cast_2001_inst_req_0, ack => type_cast_2001_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2011_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2008, dout => tmp3_2012, req => type_cast_2011_inst_req_0, ack => type_cast_2011_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2029_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2026, dout => tmp6_2030, req => type_cast_2029_inst_req_0, ack => type_cast_2029_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2039_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2036, dout => tmp8_2040, req => type_cast_2039_inst_req_0, ack => type_cast_2039_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2054_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2051, dout => tmp11_2055, req => type_cast_2054_inst_req_0, ack => type_cast_2054_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2069_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2066, dout => tmp14_2070, req => type_cast_2069_inst_req_0, ack => type_cast_2069_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2078_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_2075, dout => tmp16_2079, req => type_cast_2078_inst_req_0, ack => type_cast_2078_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2088_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_2085, dout => xx_xtrx_xi_2089, req => type_cast_2088_inst_req_0, ack => type_cast_2088_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2104_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_2101, dout => type_cast_2104_wire, req => type_cast_2104_inst_req_0, ack => type_cast_2104_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2112_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_2109, dout => tmp20_2113, req => type_cast_2112_inst_req_0, ack => type_cast_2112_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2139_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_2136, dout => tmp25_2140, req => type_cast_2139_inst_req_0, ack => type_cast_2139_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2147_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_2140, dout => type_cast_2147_wire, req => type_cast_2147_inst_req_0, ack => type_cast_2147_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2018_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2018_gather_scatter_ack_0 <= ptr_deref_2018_gather_scatter_req_0;
      aggregated_sig <= tmp4_2016;
      ptr_deref_2018_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2018_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2018_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2018_root_address_inst_ack_0 <= ptr_deref_2018_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2018_resized_base_address;
      ptr_deref_2018_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2050_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2050_gather_scatter_ack_0 <= ptr_deref_2050_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2050_data_3 & ptr_deref_2050_data_2 & ptr_deref_2050_data_1 & ptr_deref_2050_data_0;
      tmp10_2051 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2050_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2050_root_address_inst_ack_0 <= ptr_deref_2050_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2050_resized_base_address;
      ptr_deref_2050_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2065_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2065_gather_scatter_ack_0 <= ptr_deref_2065_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2065_data_3 & ptr_deref_2065_data_2 & ptr_deref_2065_data_1 & ptr_deref_2065_data_0;
      tmp13_2066 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2065_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2065_root_address_inst_ack_0 <= ptr_deref_2065_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2065_resized_base_address;
      ptr_deref_2065_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2123_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2123_gather_scatter_ack_0 <= ptr_deref_2123_gather_scatter_req_0;
      aggregated_sig <= tmp22_2121;
      ptr_deref_2123_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2123_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2123_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2123_root_address_inst_ack_0 <= ptr_deref_2123_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2123_resized_base_address;
      ptr_deref_2123_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2130_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2130_gather_scatter_ack_0 <= ptr_deref_2130_gather_scatter_req_0;
      aggregated_sig <= tmp23_2128;
      ptr_deref_2130_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2130_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2130_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2130_root_address_inst_ack_0 <= ptr_deref_2130_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2130_resized_base_address;
      ptr_deref_2130_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2135_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2135_gather_scatter_ack_0 <= ptr_deref_2135_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2135_data_3 & ptr_deref_2135_data_2 & ptr_deref_2135_data_1 & ptr_deref_2135_data_0;
      tmp24_2136 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2135_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2135_root_address_inst_ack_0 <= ptr_deref_2135_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2135_resized_base_address;
      ptr_deref_2135_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2046_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2046_resized_base_address;
      array_obj_ref_2046_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2046_root_address_inst_req_0,
          ackL => array_obj_ref_2046_root_address_inst_ack_0,
          reqR => array_obj_ref_2046_root_address_inst_req_1,
          ackR => array_obj_ref_2046_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2061_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2061_resized_base_address;
      array_obj_ref_2061_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2061_root_address_inst_req_0,
          ackL => array_obj_ref_2061_root_address_inst_ack_0,
          reqR => array_obj_ref_2061_root_address_inst_req_1,
          ackR => array_obj_ref_2061_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2007_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1998;
      tmp2_2008 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2007_inst_req_0,
          ackL => binary_2007_inst_ack_0,
          reqR => binary_2007_inst_req_1,
          ackR => binary_2007_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2025_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2008;
      tmp5_2026 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2025_inst_req_0,
          ackL => binary_2025_inst_ack_0,
          reqR => binary_2025_inst_req_1,
          ackR => binary_2025_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2035_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2008;
      tmp7_2036 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2035_inst_req_0,
          ackL => binary_2035_inst_ack_0,
          reqR => binary_2035_inst_req_1,
          ackR => binary_2035_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2074_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2055 & tmp14_2070;
      tmp15_2075 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2074_inst_req_0,
          ackL => binary_2074_inst_ack_0,
          reqR => binary_2074_inst_req_1,
          ackR => binary_2074_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2084_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2075;
      tmp17_2085 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2084_inst_req_0,
          ackL => binary_2084_inst_ack_0,
          reqR => binary_2084_inst_req_1,
          ackR => binary_2084_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2094_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_2089;
      tmp18_2095 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2094_inst_req_0,
          ackL => binary_2094_inst_ack_0,
          reqR => binary_2094_inst_req_1,
          ackR => binary_2094_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2100_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2075;
      tmp19_2101 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2100_inst_req_0,
          ackL => binary_2100_inst_ack_0,
          reqR => binary_2100_inst_req_1,
          ackR => binary_2100_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2108_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2104_wire;
      notx_xx_xi_2109 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2108_inst_req_0,
          ackL => binary_2108_inst_ack_0,
          reqR => binary_2108_inst_req_1,
          ackR => binary_2108_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2117_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_2095 & tmp20_2113;
      tmp21_2118 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2117_inst_req_0,
          ackL => binary_2117_inst_ack_0,
          reqR => binary_2117_inst_req_1,
          ackR => binary_2117_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2018_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2018_root_address;
      ptr_deref_2018_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2018_addr_0_req_0,
          ackL => ptr_deref_2018_addr_0_ack_0,
          reqR => ptr_deref_2018_addr_0_req_1,
          ackR => ptr_deref_2018_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2018_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2018_root_address;
      ptr_deref_2018_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2018_addr_1_req_0,
          ackL => ptr_deref_2018_addr_1_ack_0,
          reqR => ptr_deref_2018_addr_1_req_1,
          ackR => ptr_deref_2018_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2050_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2050_root_address;
      ptr_deref_2050_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2050_addr_0_req_0,
          ackL => ptr_deref_2050_addr_0_ack_0,
          reqR => ptr_deref_2050_addr_0_req_1,
          ackR => ptr_deref_2050_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2050_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2050_root_address;
      ptr_deref_2050_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2050_addr_1_req_0,
          ackL => ptr_deref_2050_addr_1_ack_0,
          reqR => ptr_deref_2050_addr_1_req_1,
          ackR => ptr_deref_2050_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2050_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2050_root_address;
      ptr_deref_2050_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2050_addr_2_req_0,
          ackL => ptr_deref_2050_addr_2_ack_0,
          reqR => ptr_deref_2050_addr_2_req_1,
          ackR => ptr_deref_2050_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2050_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2050_root_address;
      ptr_deref_2050_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2050_addr_3_req_0,
          ackL => ptr_deref_2050_addr_3_ack_0,
          reqR => ptr_deref_2050_addr_3_req_1,
          ackR => ptr_deref_2050_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2065_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2065_root_address;
      ptr_deref_2065_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2065_addr_0_req_0,
          ackL => ptr_deref_2065_addr_0_ack_0,
          reqR => ptr_deref_2065_addr_0_req_1,
          ackR => ptr_deref_2065_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2065_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2065_root_address;
      ptr_deref_2065_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2065_addr_1_req_0,
          ackL => ptr_deref_2065_addr_1_ack_0,
          reqR => ptr_deref_2065_addr_1_req_1,
          ackR => ptr_deref_2065_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2065_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2065_root_address;
      ptr_deref_2065_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2065_addr_2_req_0,
          ackL => ptr_deref_2065_addr_2_ack_0,
          reqR => ptr_deref_2065_addr_2_req_1,
          ackR => ptr_deref_2065_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2065_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2065_root_address;
      ptr_deref_2065_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2065_addr_3_req_0,
          ackL => ptr_deref_2065_addr_3_ack_0,
          reqR => ptr_deref_2065_addr_3_req_1,
          ackR => ptr_deref_2065_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2123_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2123_root_address;
      ptr_deref_2123_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2123_addr_0_req_0,
          ackL => ptr_deref_2123_addr_0_ack_0,
          reqR => ptr_deref_2123_addr_0_req_1,
          ackR => ptr_deref_2123_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2123_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2123_root_address;
      ptr_deref_2123_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2123_addr_1_req_0,
          ackL => ptr_deref_2123_addr_1_ack_0,
          reqR => ptr_deref_2123_addr_1_req_1,
          ackR => ptr_deref_2123_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2130_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2130_root_address;
      ptr_deref_2130_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2130_addr_0_req_0,
          ackL => ptr_deref_2130_addr_0_ack_0,
          reqR => ptr_deref_2130_addr_0_req_1,
          ackR => ptr_deref_2130_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2130_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2130_root_address;
      ptr_deref_2130_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2130_addr_1_req_0,
          ackL => ptr_deref_2130_addr_1_ack_0,
          reqR => ptr_deref_2130_addr_1_req_1,
          ackR => ptr_deref_2130_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2135_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2135_root_address;
      ptr_deref_2135_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2135_addr_0_req_0,
          ackL => ptr_deref_2135_addr_0_ack_0,
          reqR => ptr_deref_2135_addr_0_req_1,
          ackR => ptr_deref_2135_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2135_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2135_root_address;
      ptr_deref_2135_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2135_addr_1_req_0,
          ackL => ptr_deref_2135_addr_1_ack_0,
          reqR => ptr_deref_2135_addr_1_req_1,
          ackR => ptr_deref_2135_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2135_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2135_root_address;
      ptr_deref_2135_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2135_addr_2_req_0,
          ackL => ptr_deref_2135_addr_2_ack_0,
          reqR => ptr_deref_2135_addr_2_req_1,
          ackR => ptr_deref_2135_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2135_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2135_root_address;
      ptr_deref_2135_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2135_addr_3_req_0,
          ackL => ptr_deref_2135_addr_3_ack_0,
          reqR => ptr_deref_2135_addr_3_req_1,
          ackR => ptr_deref_2135_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2135_load_1 ptr_deref_2065_load_3 ptr_deref_2050_load_0 ptr_deref_2135_load_0 ptr_deref_2050_load_2 ptr_deref_2050_load_1 ptr_deref_2135_load_3 ptr_deref_2065_load_2 ptr_deref_2050_load_3 ptr_deref_2065_load_0 ptr_deref_2135_load_2 ptr_deref_2065_load_1 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2135_load_1_req_0,
        ptr_deref_2135_load_1_ack_0,
        ptr_deref_2135_load_1_req_1,
        ptr_deref_2135_load_1_ack_1,
        "ptr_deref_2135_load_1",
        "memory_space_5" ,
        ptr_deref_2135_data_1,
        ptr_deref_2135_word_address_1,
        "ptr_deref_2135_data_1",
        "ptr_deref_2135_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2065_load_3_req_0,
        ptr_deref_2065_load_3_ack_0,
        ptr_deref_2065_load_3_req_1,
        ptr_deref_2065_load_3_ack_1,
        "ptr_deref_2065_load_3",
        "memory_space_5" ,
        ptr_deref_2065_data_3,
        ptr_deref_2065_word_address_3,
        "ptr_deref_2065_data_3",
        "ptr_deref_2065_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2050_load_0_req_0,
        ptr_deref_2050_load_0_ack_0,
        ptr_deref_2050_load_0_req_1,
        ptr_deref_2050_load_0_ack_1,
        "ptr_deref_2050_load_0",
        "memory_space_5" ,
        ptr_deref_2050_data_0,
        ptr_deref_2050_word_address_0,
        "ptr_deref_2050_data_0",
        "ptr_deref_2050_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2135_load_0_req_0,
        ptr_deref_2135_load_0_ack_0,
        ptr_deref_2135_load_0_req_1,
        ptr_deref_2135_load_0_ack_1,
        "ptr_deref_2135_load_0",
        "memory_space_5" ,
        ptr_deref_2135_data_0,
        ptr_deref_2135_word_address_0,
        "ptr_deref_2135_data_0",
        "ptr_deref_2135_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2050_load_2_req_0,
        ptr_deref_2050_load_2_ack_0,
        ptr_deref_2050_load_2_req_1,
        ptr_deref_2050_load_2_ack_1,
        "ptr_deref_2050_load_2",
        "memory_space_5" ,
        ptr_deref_2050_data_2,
        ptr_deref_2050_word_address_2,
        "ptr_deref_2050_data_2",
        "ptr_deref_2050_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2050_load_1_req_0,
        ptr_deref_2050_load_1_ack_0,
        ptr_deref_2050_load_1_req_1,
        ptr_deref_2050_load_1_ack_1,
        "ptr_deref_2050_load_1",
        "memory_space_5" ,
        ptr_deref_2050_data_1,
        ptr_deref_2050_word_address_1,
        "ptr_deref_2050_data_1",
        "ptr_deref_2050_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2135_load_3_req_0,
        ptr_deref_2135_load_3_ack_0,
        ptr_deref_2135_load_3_req_1,
        ptr_deref_2135_load_3_ack_1,
        "ptr_deref_2135_load_3",
        "memory_space_5" ,
        ptr_deref_2135_data_3,
        ptr_deref_2135_word_address_3,
        "ptr_deref_2135_data_3",
        "ptr_deref_2135_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2065_load_2_req_0,
        ptr_deref_2065_load_2_ack_0,
        ptr_deref_2065_load_2_req_1,
        ptr_deref_2065_load_2_ack_1,
        "ptr_deref_2065_load_2",
        "memory_space_5" ,
        ptr_deref_2065_data_2,
        ptr_deref_2065_word_address_2,
        "ptr_deref_2065_data_2",
        "ptr_deref_2065_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2050_load_3_req_0,
        ptr_deref_2050_load_3_ack_0,
        ptr_deref_2050_load_3_req_1,
        ptr_deref_2050_load_3_ack_1,
        "ptr_deref_2050_load_3",
        "memory_space_5" ,
        ptr_deref_2050_data_3,
        ptr_deref_2050_word_address_3,
        "ptr_deref_2050_data_3",
        "ptr_deref_2050_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2065_load_0_req_0,
        ptr_deref_2065_load_0_ack_0,
        ptr_deref_2065_load_0_req_1,
        ptr_deref_2065_load_0_ack_1,
        "ptr_deref_2065_load_0",
        "memory_space_5" ,
        ptr_deref_2065_data_0,
        ptr_deref_2065_word_address_0,
        "ptr_deref_2065_data_0",
        "ptr_deref_2065_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2135_load_2_req_0,
        ptr_deref_2135_load_2_ack_0,
        ptr_deref_2135_load_2_req_1,
        ptr_deref_2135_load_2_ack_1,
        "ptr_deref_2135_load_2",
        "memory_space_5" ,
        ptr_deref_2135_data_2,
        ptr_deref_2135_word_address_2,
        "ptr_deref_2135_data_2",
        "ptr_deref_2135_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2065_load_1_req_0,
        ptr_deref_2065_load_1_ack_0,
        ptr_deref_2065_load_1_req_1,
        ptr_deref_2065_load_1_ack_1,
        "ptr_deref_2065_load_1",
        "memory_space_5" ,
        ptr_deref_2065_data_1,
        ptr_deref_2065_word_address_1,
        "ptr_deref_2065_data_1",
        "ptr_deref_2065_word_address_1" -- 
      );
      reqL(11) <= ptr_deref_2135_load_1_req_0;
      reqL(10) <= ptr_deref_2065_load_3_req_0;
      reqL(9) <= ptr_deref_2050_load_0_req_0;
      reqL(8) <= ptr_deref_2135_load_0_req_0;
      reqL(7) <= ptr_deref_2050_load_2_req_0;
      reqL(6) <= ptr_deref_2050_load_1_req_0;
      reqL(5) <= ptr_deref_2135_load_3_req_0;
      reqL(4) <= ptr_deref_2065_load_2_req_0;
      reqL(3) <= ptr_deref_2050_load_3_req_0;
      reqL(2) <= ptr_deref_2065_load_0_req_0;
      reqL(1) <= ptr_deref_2135_load_2_req_0;
      reqL(0) <= ptr_deref_2065_load_1_req_0;
      ptr_deref_2135_load_1_ack_0 <= ackL(11);
      ptr_deref_2065_load_3_ack_0 <= ackL(10);
      ptr_deref_2050_load_0_ack_0 <= ackL(9);
      ptr_deref_2135_load_0_ack_0 <= ackL(8);
      ptr_deref_2050_load_2_ack_0 <= ackL(7);
      ptr_deref_2050_load_1_ack_0 <= ackL(6);
      ptr_deref_2135_load_3_ack_0 <= ackL(5);
      ptr_deref_2065_load_2_ack_0 <= ackL(4);
      ptr_deref_2050_load_3_ack_0 <= ackL(3);
      ptr_deref_2065_load_0_ack_0 <= ackL(2);
      ptr_deref_2135_load_2_ack_0 <= ackL(1);
      ptr_deref_2065_load_1_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2135_load_1_req_1;
      reqR(10) <= ptr_deref_2065_load_3_req_1;
      reqR(9) <= ptr_deref_2050_load_0_req_1;
      reqR(8) <= ptr_deref_2135_load_0_req_1;
      reqR(7) <= ptr_deref_2050_load_2_req_1;
      reqR(6) <= ptr_deref_2050_load_1_req_1;
      reqR(5) <= ptr_deref_2135_load_3_req_1;
      reqR(4) <= ptr_deref_2065_load_2_req_1;
      reqR(3) <= ptr_deref_2050_load_3_req_1;
      reqR(2) <= ptr_deref_2065_load_0_req_1;
      reqR(1) <= ptr_deref_2135_load_2_req_1;
      reqR(0) <= ptr_deref_2065_load_1_req_1;
      ptr_deref_2135_load_1_ack_1 <= ackR(11);
      ptr_deref_2065_load_3_ack_1 <= ackR(10);
      ptr_deref_2050_load_0_ack_1 <= ackR(9);
      ptr_deref_2135_load_0_ack_1 <= ackR(8);
      ptr_deref_2050_load_2_ack_1 <= ackR(7);
      ptr_deref_2050_load_1_ack_1 <= ackR(6);
      ptr_deref_2135_load_3_ack_1 <= ackR(5);
      ptr_deref_2065_load_2_ack_1 <= ackR(4);
      ptr_deref_2050_load_3_ack_1 <= ackR(3);
      ptr_deref_2065_load_0_ack_1 <= ackR(2);
      ptr_deref_2135_load_2_ack_1 <= ackR(1);
      ptr_deref_2065_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_2135_word_address_1 & ptr_deref_2065_word_address_3 & ptr_deref_2050_word_address_0 & ptr_deref_2135_word_address_0 & ptr_deref_2050_word_address_2 & ptr_deref_2050_word_address_1 & ptr_deref_2135_word_address_3 & ptr_deref_2065_word_address_2 & ptr_deref_2050_word_address_3 & ptr_deref_2065_word_address_0 & ptr_deref_2135_word_address_2 & ptr_deref_2065_word_address_1;
      ptr_deref_2135_data_1 <= data_out(95 downto 88);
      ptr_deref_2065_data_3 <= data_out(87 downto 80);
      ptr_deref_2050_data_0 <= data_out(79 downto 72);
      ptr_deref_2135_data_0 <= data_out(71 downto 64);
      ptr_deref_2050_data_2 <= data_out(63 downto 56);
      ptr_deref_2050_data_1 <= data_out(55 downto 48);
      ptr_deref_2135_data_3 <= data_out(47 downto 40);
      ptr_deref_2065_data_2 <= data_out(39 downto 32);
      ptr_deref_2050_data_3 <= data_out(31 downto 24);
      ptr_deref_2065_data_0 <= data_out(23 downto 16);
      ptr_deref_2135_data_2 <= data_out(15 downto 8);
      ptr_deref_2065_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2018_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2018_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2018_word_address_0) &  " data ptr_deref_2018_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2018_data_0) severity note; --
        end if;
        if ptr_deref_2018_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2018_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2018_word_address_1) &  " data ptr_deref_2018_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2018_data_1) severity note; --
        end if;
        if ptr_deref_2130_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2130_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2130_word_address_1) &  " data ptr_deref_2130_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2130_data_1) severity note; --
        end if;
        if ptr_deref_2130_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2130_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2130_word_address_0) &  " data ptr_deref_2130_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2130_data_0) severity note; --
        end if;
        if ptr_deref_2123_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2123_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2123_word_address_1) &  " data ptr_deref_2123_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2123_data_1) severity note; --
        end if;
        if ptr_deref_2123_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2123_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2123_word_address_0) &  " data ptr_deref_2123_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2123_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2018_store_0 ptr_deref_2018_store_1 ptr_deref_2130_store_1 ptr_deref_2130_store_0 ptr_deref_2123_store_1 ptr_deref_2123_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2018_store_0_req_0;
      reqL(4) <= ptr_deref_2018_store_1_req_0;
      reqL(3) <= ptr_deref_2130_store_1_req_0;
      reqL(2) <= ptr_deref_2130_store_0_req_0;
      reqL(1) <= ptr_deref_2123_store_1_req_0;
      reqL(0) <= ptr_deref_2123_store_0_req_0;
      ptr_deref_2018_store_0_ack_0 <= ackL(5);
      ptr_deref_2018_store_1_ack_0 <= ackL(4);
      ptr_deref_2130_store_1_ack_0 <= ackL(3);
      ptr_deref_2130_store_0_ack_0 <= ackL(2);
      ptr_deref_2123_store_1_ack_0 <= ackL(1);
      ptr_deref_2123_store_0_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2018_store_0_req_1;
      reqR(4) <= ptr_deref_2018_store_1_req_1;
      reqR(3) <= ptr_deref_2130_store_1_req_1;
      reqR(2) <= ptr_deref_2130_store_0_req_1;
      reqR(1) <= ptr_deref_2123_store_1_req_1;
      reqR(0) <= ptr_deref_2123_store_0_req_1;
      ptr_deref_2018_store_0_ack_1 <= ackR(5);
      ptr_deref_2018_store_1_ack_1 <= ackR(4);
      ptr_deref_2130_store_1_ack_1 <= ackR(3);
      ptr_deref_2130_store_0_ack_1 <= ackR(2);
      ptr_deref_2123_store_1_ack_1 <= ackR(1);
      ptr_deref_2123_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2018_word_address_0 & ptr_deref_2018_word_address_1 & ptr_deref_2130_word_address_1 & ptr_deref_2130_word_address_0 & ptr_deref_2123_word_address_1 & ptr_deref_2123_word_address_0;
      data_in <= ptr_deref_2018_data_0 & ptr_deref_2018_data_1 & ptr_deref_2130_data_1 & ptr_deref_2130_data_0 & ptr_deref_2123_data_1 & ptr_deref_2123_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_1996_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_1996_inst_ack_0 then -- 
            assert false report " ReadPipe to1_in0 to wire simple_obj_ref_1996_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_1996_inst_req_0;
      simple_obj_ref_1996_inst_ack_0 <= ack(0);
      simple_obj_ref_1996_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to1_in0_pipe_read_req(0),
          oack => to1_in0_pipe_read_ack(0),
          odata => to1_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2141_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_2143_wire_constant value="  &  convert_slv_to_hex_string(type_cast_2143_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2141_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2141_inst_req_0;
      simple_obj_ref_2141_inst_ack_0 <= ack(0);
      data_in <= type_cast_2143_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2145_inst_ack_0 then -- 
          assert false report " WritePipe tofpga1_out0 from wire type_cast_2147_wire value="  &  convert_slv_to_hex_string(type_cast_2147_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2145_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2145_inst_req_0;
      simple_obj_ref_2145_inst_ack_0 <= ack(0);
      data_in <= type_cast_2147_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga1_out0_pipe_write_req(0),
          oack => tofpga1_out0_pipe_write_ack(0),
          odata => tofpga1_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2128_call call_stmt_2121_call call_stmt_2016_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2128_call_req_0;
      reqL(1) <= call_stmt_2121_call_req_0;
      reqL(0) <= call_stmt_2016_call_req_0;
      call_stmt_2128_call_ack_0 <= ackL(2);
      call_stmt_2121_call_ack_0 <= ackL(1);
      call_stmt_2016_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2128_call_req_1;
      reqR(1) <= call_stmt_2121_call_req_1;
      reqR(0) <= call_stmt_2016_call_req_1;
      call_stmt_2128_call_ack_1 <= ackR(2);
      call_stmt_2121_call_ack_1 <= ackR(1);
      call_stmt_2016_call_ack_1 <= ackR(0);
      data_in <= tmp21_2118 & tmp16_2079 & type_cast_2014_wire_constant;
      tmp23_2128 <= data_out(47 downto 32);
      tmp22_2121 <= data_out(31 downto 16);
      tmp4_2016 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to2_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to2_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to2_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga2_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to2;
architecture Default of ahir_glue_to2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to2_CP_10549_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_2290_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2221_base_resize_ack_0 : boolean;
  signal type_cast_2214_inst_req_0 : boolean;
  signal ptr_deref_2295_addr_0_req_0 : boolean;
  signal ptr_deref_2283_store_1_ack_1 : boolean;
  signal ptr_deref_2295_addr_0_req_1 : boolean;
  signal binary_2234_inst_req_1 : boolean;
  signal binary_2234_inst_ack_0 : boolean;
  signal call_stmt_2288_call_req_1 : boolean;
  signal type_cast_2214_inst_ack_0 : boolean;
  signal ptr_deref_2225_addr_0_ack_0 : boolean;
  signal ptr_deref_2290_gather_scatter_ack_0 : boolean;
  signal binary_2268_inst_ack_1 : boolean;
  signal ptr_deref_2290_root_address_inst_ack_0 : boolean;
  signal type_cast_2264_inst_ack_0 : boolean;
  signal array_obj_ref_2221_base_resize_req_0 : boolean;
  signal ptr_deref_2290_gather_scatter_req_0 : boolean;
  signal type_cast_2238_inst_req_0 : boolean;
  signal binary_2234_inst_req_0 : boolean;
  signal binary_2244_inst_req_1 : boolean;
  signal ptr_deref_2225_base_resize_req_0 : boolean;
  signal ptr_deref_2225_addr_1_req_0 : boolean;
  signal ptr_deref_2295_load_1_req_0 : boolean;
  signal ptr_deref_2290_addr_0_req_0 : boolean;
  signal ptr_deref_2290_addr_1_ack_1 : boolean;
  signal ptr_deref_2295_load_1_ack_0 : boolean;
  signal ptr_deref_2295_addr_3_ack_1 : boolean;
  signal binary_2244_inst_ack_1 : boolean;
  signal ptr_deref_2295_load_3_req_0 : boolean;
  signal ptr_deref_2295_addr_3_req_0 : boolean;
  signal ptr_deref_2290_addr_1_req_1 : boolean;
  signal ptr_deref_2225_addr_0_req_1 : boolean;
  signal ptr_deref_2225_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2283_addr_1_req_1 : boolean;
  signal type_cast_2264_inst_req_0 : boolean;
  signal ptr_deref_2225_root_address_inst_ack_0 : boolean;
  signal binary_2260_inst_ack_0 : boolean;
  signal binary_2268_inst_req_0 : boolean;
  signal ptr_deref_2290_store_0_req_0 : boolean;
  signal ptr_deref_2290_base_resize_req_0 : boolean;
  signal binary_2234_inst_ack_1 : boolean;
  signal ptr_deref_2290_store_1_ack_0 : boolean;
  signal ptr_deref_2290_store_0_ack_0 : boolean;
  signal ptr_deref_2225_load_0_ack_0 : boolean;
  signal ptr_deref_2225_addr_3_req_0 : boolean;
  signal ptr_deref_2225_addr_2_ack_1 : boolean;
  signal ptr_deref_2225_addr_3_ack_1 : boolean;
  signal ptr_deref_2283_addr_1_req_0 : boolean;
  signal ptr_deref_2295_addr_2_ack_0 : boolean;
  signal ptr_deref_2225_load_0_req_0 : boolean;
  signal ptr_deref_2283_addr_0_req_1 : boolean;
  signal binary_2260_inst_req_1 : boolean;
  signal binary_2268_inst_ack_0 : boolean;
  signal binary_2244_inst_req_0 : boolean;
  signal ptr_deref_2283_addr_1_ack_0 : boolean;
  signal ptr_deref_2225_load_0_ack_1 : boolean;
  signal ptr_deref_2283_store_1_ack_0 : boolean;
  signal ptr_deref_2295_addr_1_req_0 : boolean;
  signal binary_2268_inst_req_1 : boolean;
  signal binary_2244_inst_ack_0 : boolean;
  signal ptr_deref_2225_base_resize_ack_0 : boolean;
  signal ptr_deref_2225_load_1_req_1 : boolean;
  signal ptr_deref_2225_load_1_req_0 : boolean;
  signal call_stmt_2281_call_req_1 : boolean;
  signal ptr_deref_2283_addr_1_ack_1 : boolean;
  signal ptr_deref_2283_gather_scatter_req_0 : boolean;
  signal ptr_deref_2295_base_resize_req_0 : boolean;
  signal ptr_deref_2290_addr_0_ack_0 : boolean;
  signal type_cast_2248_inst_req_0 : boolean;
  signal ptr_deref_2225_load_1_ack_1 : boolean;
  signal ptr_deref_2290_store_1_req_0 : boolean;
  signal ptr_deref_2295_load_2_ack_1 : boolean;
  signal ptr_deref_2295_load_1_ack_1 : boolean;
  signal ptr_deref_2290_addr_1_req_0 : boolean;
  signal ptr_deref_2283_store_1_req_1 : boolean;
  signal type_cast_2272_inst_req_0 : boolean;
  signal ptr_deref_2283_addr_0_ack_0 : boolean;
  signal ptr_deref_2295_load_0_req_0 : boolean;
  signal ptr_deref_2225_load_2_req_0 : boolean;
  signal type_cast_2248_inst_ack_0 : boolean;
  signal ptr_deref_2225_load_1_ack_0 : boolean;
  signal ptr_deref_2290_store_0_req_1 : boolean;
  signal ptr_deref_2295_load_0_req_1 : boolean;
  signal type_cast_2238_inst_ack_0 : boolean;
  signal ptr_deref_2295_addr_0_ack_0 : boolean;
  signal ptr_deref_2225_addr_0_ack_1 : boolean;
  signal ptr_deref_2283_store_1_req_0 : boolean;
  signal ptr_deref_2295_addr_2_req_0 : boolean;
  signal ptr_deref_2225_addr_3_req_1 : boolean;
  signal ptr_deref_2225_addr_3_ack_0 : boolean;
  signal ptr_deref_2225_load_2_ack_0 : boolean;
  signal ptr_deref_2295_addr_0_ack_1 : boolean;
  signal type_cast_2229_inst_req_0 : boolean;
  signal type_cast_2272_inst_ack_0 : boolean;
  signal ptr_deref_2283_base_resize_req_0 : boolean;
  signal ptr_deref_2290_store_0_ack_1 : boolean;
  signal ptr_deref_2283_base_resize_ack_0 : boolean;
  signal ptr_deref_2295_base_resize_ack_0 : boolean;
  signal binary_2260_inst_ack_1 : boolean;
  signal array_obj_ref_2221_root_address_inst_ack_1 : boolean;
  signal call_stmt_2281_call_ack_1 : boolean;
  signal ptr_deref_2295_addr_1_ack_1 : boolean;
  signal ptr_deref_2295_load_3_req_1 : boolean;
  signal ptr_deref_2295_load_3_ack_1 : boolean;
  signal ptr_deref_2295_addr_3_ack_0 : boolean;
  signal ptr_deref_2225_load_2_req_1 : boolean;
  signal ptr_deref_2283_gather_scatter_ack_0 : boolean;
  signal binary_2254_inst_req_0 : boolean;
  signal binary_2254_inst_ack_0 : boolean;
  signal binary_2277_inst_ack_1 : boolean;
  signal ptr_deref_2290_addr_0_req_1 : boolean;
  signal ptr_deref_2283_root_address_inst_req_0 : boolean;
  signal ptr_deref_2290_addr_0_ack_1 : boolean;
  signal binary_2254_inst_req_1 : boolean;
  signal ptr_deref_2283_root_address_inst_ack_0 : boolean;
  signal binary_2254_inst_ack_1 : boolean;
  signal ptr_deref_2290_store_1_req_1 : boolean;
  signal call_stmt_2288_call_ack_1 : boolean;
  signal ptr_deref_2283_store_0_req_1 : boolean;
  signal ptr_deref_2290_base_resize_ack_0 : boolean;
  signal call_stmt_2281_call_req_0 : boolean;
  signal array_obj_ref_2221_final_reg_ack_0 : boolean;
  signal ptr_deref_2283_store_0_ack_0 : boolean;
  signal ptr_deref_2295_load_1_req_1 : boolean;
  signal ptr_deref_2295_addr_1_req_1 : boolean;
  signal ptr_deref_2295_gather_scatter_req_0 : boolean;
  signal ptr_deref_2225_load_3_req_0 : boolean;
  signal ptr_deref_2283_store_0_ack_1 : boolean;
  signal type_cast_2229_inst_ack_0 : boolean;
  signal ptr_deref_2295_addr_1_ack_0 : boolean;
  signal ptr_deref_2290_addr_1_ack_0 : boolean;
  signal ptr_deref_2295_load_2_req_1 : boolean;
  signal binary_2277_inst_req_1 : boolean;
  signal ptr_deref_2295_load_3_ack_0 : boolean;
  signal ptr_deref_2225_root_address_inst_req_0 : boolean;
  signal ptr_deref_2225_load_2_ack_1 : boolean;
  signal ptr_deref_2295_load_2_req_0 : boolean;
  signal ptr_deref_2225_load_3_ack_0 : boolean;
  signal ptr_deref_2225_addr_0_req_0 : boolean;
  signal ptr_deref_2283_addr_0_req_0 : boolean;
  signal ptr_deref_2283_store_0_req_0 : boolean;
  signal ptr_deref_2295_root_address_inst_req_0 : boolean;
  signal ptr_deref_2295_load_0_ack_0 : boolean;
  signal binary_2260_inst_req_0 : boolean;
  signal ptr_deref_2295_addr_3_req_1 : boolean;
  signal ptr_deref_2295_addr_2_req_1 : boolean;
  signal ptr_deref_2295_load_0_ack_1 : boolean;
  signal type_cast_2299_inst_req_0 : boolean;
  signal ptr_deref_2225_addr_1_ack_0 : boolean;
  signal type_cast_2299_inst_ack_0 : boolean;
  signal ptr_deref_2295_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2225_addr_1_req_1 : boolean;
  signal call_stmt_2288_call_req_0 : boolean;
  signal ptr_deref_2225_addr_1_ack_1 : boolean;
  signal call_stmt_2288_call_ack_0 : boolean;
  signal ptr_deref_2225_load_0_req_1 : boolean;
  signal ptr_deref_2295_load_2_ack_0 : boolean;
  signal ptr_deref_2290_store_1_ack_1 : boolean;
  signal ptr_deref_2225_load_3_req_1 : boolean;
  signal ptr_deref_2283_addr_0_ack_1 : boolean;
  signal ptr_deref_2225_addr_2_req_0 : boolean;
  signal ptr_deref_2225_load_3_ack_1 : boolean;
  signal ptr_deref_2225_addr_2_ack_0 : boolean;
  signal ptr_deref_2225_addr_2_req_1 : boolean;
  signal ptr_deref_2225_gather_scatter_req_0 : boolean;
  signal call_stmt_2281_call_ack_0 : boolean;
  signal array_obj_ref_2221_final_reg_req_0 : boolean;
  signal binary_2277_inst_ack_0 : boolean;
  signal binary_2277_inst_req_0 : boolean;
  signal array_obj_ref_2221_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2221_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2221_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2295_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2295_addr_2_ack_1 : boolean;
  signal simple_obj_ref_2156_inst_req_0 : boolean;
  signal simple_obj_ref_2156_inst_ack_0 : boolean;
  signal type_cast_2157_inst_req_0 : boolean;
  signal type_cast_2157_inst_ack_0 : boolean;
  signal type_cast_2161_inst_req_0 : boolean;
  signal type_cast_2161_inst_ack_0 : boolean;
  signal binary_2167_inst_req_0 : boolean;
  signal binary_2167_inst_ack_0 : boolean;
  signal binary_2167_inst_req_1 : boolean;
  signal binary_2167_inst_ack_1 : boolean;
  signal type_cast_2171_inst_req_0 : boolean;
  signal type_cast_2171_inst_ack_0 : boolean;
  signal call_stmt_2176_call_req_0 : boolean;
  signal call_stmt_2176_call_ack_0 : boolean;
  signal call_stmt_2176_call_req_1 : boolean;
  signal call_stmt_2176_call_ack_1 : boolean;
  signal ptr_deref_2178_base_resize_req_0 : boolean;
  signal ptr_deref_2178_base_resize_ack_0 : boolean;
  signal ptr_deref_2178_root_address_inst_req_0 : boolean;
  signal ptr_deref_2178_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2178_addr_0_req_0 : boolean;
  signal ptr_deref_2178_addr_0_ack_0 : boolean;
  signal ptr_deref_2178_addr_0_req_1 : boolean;
  signal ptr_deref_2178_addr_0_ack_1 : boolean;
  signal ptr_deref_2178_addr_1_req_0 : boolean;
  signal ptr_deref_2178_addr_1_ack_0 : boolean;
  signal ptr_deref_2178_addr_1_req_1 : boolean;
  signal ptr_deref_2178_addr_1_ack_1 : boolean;
  signal ptr_deref_2178_gather_scatter_req_0 : boolean;
  signal ptr_deref_2178_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2178_store_0_req_0 : boolean;
  signal ptr_deref_2178_store_0_ack_0 : boolean;
  signal ptr_deref_2178_store_1_req_0 : boolean;
  signal ptr_deref_2178_store_1_ack_0 : boolean;
  signal ptr_deref_2178_store_0_req_1 : boolean;
  signal ptr_deref_2178_store_0_ack_1 : boolean;
  signal ptr_deref_2178_store_1_req_1 : boolean;
  signal ptr_deref_2178_store_1_ack_1 : boolean;
  signal binary_2185_inst_req_0 : boolean;
  signal binary_2185_inst_ack_0 : boolean;
  signal binary_2185_inst_req_1 : boolean;
  signal binary_2185_inst_ack_1 : boolean;
  signal type_cast_2189_inst_req_0 : boolean;
  signal type_cast_2189_inst_ack_0 : boolean;
  signal binary_2195_inst_req_0 : boolean;
  signal binary_2195_inst_ack_0 : boolean;
  signal binary_2195_inst_req_1 : boolean;
  signal binary_2195_inst_ack_1 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal array_obj_ref_2206_base_resize_req_0 : boolean;
  signal array_obj_ref_2206_base_resize_ack_0 : boolean;
  signal array_obj_ref_2206_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2206_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2206_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2206_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2206_final_reg_req_0 : boolean;
  signal array_obj_ref_2206_final_reg_ack_0 : boolean;
  signal ptr_deref_2210_base_resize_req_0 : boolean;
  signal ptr_deref_2210_base_resize_ack_0 : boolean;
  signal ptr_deref_2210_root_address_inst_req_0 : boolean;
  signal ptr_deref_2210_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2210_addr_0_req_0 : boolean;
  signal ptr_deref_2210_addr_0_ack_0 : boolean;
  signal ptr_deref_2210_addr_0_req_1 : boolean;
  signal ptr_deref_2210_addr_0_ack_1 : boolean;
  signal ptr_deref_2210_addr_1_req_0 : boolean;
  signal ptr_deref_2210_addr_1_ack_0 : boolean;
  signal ptr_deref_2210_addr_1_req_1 : boolean;
  signal ptr_deref_2210_addr_1_ack_1 : boolean;
  signal ptr_deref_2210_addr_2_req_0 : boolean;
  signal ptr_deref_2210_addr_2_ack_0 : boolean;
  signal ptr_deref_2210_addr_2_req_1 : boolean;
  signal ptr_deref_2210_addr_2_ack_1 : boolean;
  signal ptr_deref_2210_addr_3_req_0 : boolean;
  signal ptr_deref_2210_addr_3_ack_0 : boolean;
  signal ptr_deref_2210_addr_3_req_1 : boolean;
  signal ptr_deref_2210_addr_3_ack_1 : boolean;
  signal ptr_deref_2210_load_0_req_0 : boolean;
  signal ptr_deref_2210_load_0_ack_0 : boolean;
  signal ptr_deref_2210_load_1_req_0 : boolean;
  signal ptr_deref_2210_load_1_ack_0 : boolean;
  signal ptr_deref_2210_load_2_req_0 : boolean;
  signal ptr_deref_2210_load_2_ack_0 : boolean;
  signal ptr_deref_2210_load_3_req_0 : boolean;
  signal ptr_deref_2210_load_3_ack_0 : boolean;
  signal ptr_deref_2210_load_0_req_1 : boolean;
  signal ptr_deref_2210_load_0_ack_1 : boolean;
  signal ptr_deref_2210_load_1_req_1 : boolean;
  signal ptr_deref_2210_load_1_ack_1 : boolean;
  signal ptr_deref_2210_load_2_req_1 : boolean;
  signal ptr_deref_2210_load_2_ack_1 : boolean;
  signal ptr_deref_2210_load_3_req_1 : boolean;
  signal ptr_deref_2210_load_3_ack_1 : boolean;
  signal ptr_deref_2210_gather_scatter_req_0 : boolean;
  signal ptr_deref_2210_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_2301_inst_req_0 : boolean;
  signal simple_obj_ref_2301_inst_ack_0 : boolean;
  signal type_cast_2307_inst_req_0 : boolean;
  signal type_cast_2307_inst_ack_0 : boolean;
  signal simple_obj_ref_2305_inst_req_0 : boolean;
  signal simple_obj_ref_2305_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to2_CP_10549: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_10640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2176_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_11165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2281_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_11463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2301_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_2157_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_10590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_2156_inst_req_0); -- 
    ack_10591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2156_inst_ack_0, ack => cp_elements(8)); -- 
    ack_10596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2161_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_10609_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2161_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2167_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_10619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2167_inst_ack_0, ack => cp_elements(18)); -- 
    cr_10620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2167_inst_req_1); -- 
    ca_10621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2167_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2171_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_10631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2171_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_10641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2176_call_ack_0, ack => cp_elements(24)); -- 
    ccr_10645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2176_call_req_1); -- 
    cca_10646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2176_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_10692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2178_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_10665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2178_base_resize_req_0); -- 
    base_resize_ack_10666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_10670_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2178_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2178_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_10678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2178_addr_0_req_0); -- 
    ra_10679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_10680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2178_addr_0_req_1); -- 
    ca_10681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_10685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2178_addr_1_req_0); -- 
    ra_10686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_10687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2178_addr_1_req_1); -- 
    ca_10688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2178_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_10700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2178_store_0_req_0); -- 
    ra_10701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_10705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2178_store_1_req_0); -- 
    ra_10706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_10716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2178_store_0_req_1); -- 
    ca_10717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_10721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2178_store_1_req_1); -- 
    ca_10722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2178_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10731_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2185_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_10732_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2185_inst_ack_0, ack => cp_elements(55)); -- 
    cr_10733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2185_inst_req_1); -- 
    ca_10734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2185_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2189_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_10744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2195_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_10754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2195_inst_ack_0, ack => cp_elements(63)); -- 
    cr_10755_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2195_inst_req_1); -- 
    ca_10756_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2195_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10765_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2199_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_10766_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_10790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2206_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_10777_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2206_base_resize_req_0); -- 
    base_resize_ack_10778_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2206_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_10783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2206_root_address_inst_req_0); -- 
    plus_base_ra_10784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2206_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_10785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2206_root_address_inst_req_1); -- 
    plus_base_ca_10786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2206_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2206_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_10804_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2210_base_resize_req_0); -- 
    base_resize_ack_10805_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_10809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2210_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2210_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_10817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2210_addr_0_req_0); -- 
    ra_10818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_10819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2210_addr_0_req_1); -- 
    ca_10820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_10824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2210_addr_1_req_0); -- 
    ra_10825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_10826_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2210_addr_1_req_1); -- 
    ca_10827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_10831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2210_addr_2_req_0); -- 
    ra_10832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_10833_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2210_addr_2_req_1); -- 
    ca_10834_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_10838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2210_addr_3_req_0); -- 
    ra_10839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_10840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2210_addr_3_req_1); -- 
    ca_10841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_10851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2210_load_0_req_0); -- 
    ra_10852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_10856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2210_load_1_req_0); -- 
    ra_10857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_10861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2210_load_2_req_0); -- 
    ra_10862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_10866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2210_load_3_req_0); -- 
    ra_10867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_10877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2210_load_0_req_1); -- 
    ca_10878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_10882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2210_load_1_req_1); -- 
    ca_10883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_10887_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2210_load_2_req_1); -- 
    ca_10888_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_10892_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2210_load_3_req_1); -- 
    ca_10893_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_10894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2210_gather_scatter_req_0); -- 
    merge_ack_10895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2210_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2214_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_10905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_10929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2221_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_10916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2221_base_resize_req_0); -- 
    base_resize_ack_10917_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2221_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_10922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2221_root_address_inst_req_0); -- 
    plus_base_ra_10923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2221_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_10924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2221_root_address_inst_req_1); -- 
    plus_base_ca_10925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2221_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2221_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_10943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2225_base_resize_req_0); -- 
    base_resize_ack_10944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_10948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2225_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2225_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_10956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2225_addr_0_req_0); -- 
    ra_10957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_10958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2225_addr_0_req_1); -- 
    ca_10959_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_10963_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2225_addr_1_req_0); -- 
    ra_10964_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_10965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2225_addr_1_req_1); -- 
    ca_10966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_10970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2225_addr_2_req_0); -- 
    ra_10971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_10972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2225_addr_2_req_1); -- 
    ca_10973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_10977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2225_addr_3_req_0); -- 
    ra_10978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_10979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2225_addr_3_req_1); -- 
    ca_10980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_10990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2225_load_0_req_0); -- 
    ra_10991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_10995_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2225_load_1_req_0); -- 
    ra_10996_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_11000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2225_load_2_req_0); -- 
    ra_11001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_11005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2225_load_3_req_0); -- 
    ra_11006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_11016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2225_load_0_req_1); -- 
    ca_11017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_11021_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2225_load_1_req_1); -- 
    ca_11022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_11026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2225_load_2_req_1); -- 
    ca_11027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_11031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2225_load_3_req_1); -- 
    ca_11032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_11033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2225_gather_scatter_req_0); -- 
    merge_ack_11034_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2225_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2229_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_11044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2229_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_2234_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_11055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2234_inst_ack_0, ack => cp_elements(162)); -- 
    cr_11056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_2234_inst_req_1); -- 
    cp_elements(163) <= binary_2234_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_2238_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_11067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_2244_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_11077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2244_inst_ack_0, ack => cp_elements(171)); -- 
    cr_11078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_2244_inst_req_1); -- 
    ca_11079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2244_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_2248_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_11089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2254_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_11099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2254_inst_ack_0, ack => cp_elements(178)); -- 
    cr_11100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_2254_inst_req_1); -- 
    ca_11101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2254_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_2260_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_11111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2260_inst_ack_0, ack => cp_elements(183)); -- 
    cr_11112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2260_inst_req_1); -- 
    ca_11113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2260_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_2268_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_2264_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_11125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2264_inst_ack_0, ack => cp_elements(189)); -- 
    ra_11130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2268_inst_ack_0, ack => cp_elements(190)); -- 
    cr_11131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_2268_inst_req_1); -- 
    ca_11132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2268_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_2272_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_11142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_2277_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_11153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2277_inst_ack_0, ack => cp_elements(197)); -- 
    cr_11154_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_2277_inst_req_1); -- 
    ca_11155_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2277_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_11166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2281_call_ack_0, ack => cp_elements(200)); -- 
    ccr_11170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_2281_call_req_1); -- 
    cca_11171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2281_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11217_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_2283_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_11190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_2283_base_resize_req_0); -- 
    base_resize_ack_11191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_11195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2283_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_2283_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_11203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2283_addr_0_req_0); -- 
    ra_11204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_11205_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_2283_addr_0_req_1); -- 
    ca_11206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_11210_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_2283_addr_1_req_0); -- 
    ra_11211_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_11212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2283_addr_1_req_1); -- 
    ca_11213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_2283_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_11225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2283_store_0_req_0); -- 
    ra_11226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_11230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2283_store_1_req_0); -- 
    ra_11231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_11241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_2283_store_0_req_1); -- 
    ca_11242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_11246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_2283_store_1_req_1); -- 
    ca_11247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_11257_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_2288_call_req_0); -- 
    cra_11258_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2288_call_ack_0, ack => cp_elements(227)); -- 
    ccr_11262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_2288_call_req_1); -- 
    cca_11263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2288_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_2290_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_11282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_2290_base_resize_req_0); -- 
    base_resize_ack_11283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_11287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_2290_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_2290_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_11295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_2290_addr_0_req_0); -- 
    ra_11296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_11297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_2290_addr_0_req_1); -- 
    ca_11298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_11302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_2290_addr_1_req_0); -- 
    ra_11303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_11304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_2290_addr_1_req_1); -- 
    ca_11305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_2290_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_11317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_2290_store_0_req_0); -- 
    ra_11318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_11322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2290_store_1_req_0); -- 
    ra_11323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_11333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_2290_store_0_req_1); -- 
    ca_11334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_11338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2290_store_1_req_1); -- 
    ca_11339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2290_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_11352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_2295_base_resize_req_0); -- 
    base_resize_ack_11353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_11357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_2295_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_2295_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_11365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_2295_addr_0_req_0); -- 
    ra_11366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_11367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2295_addr_0_req_1); -- 
    ca_11368_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_11372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2295_addr_1_req_0); -- 
    ra_11373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_11374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_2295_addr_1_req_1); -- 
    ca_11375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_11379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_2295_addr_2_req_0); -- 
    ra_11380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_11381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_2295_addr_2_req_1); -- 
    ca_11382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_11386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_2295_addr_3_req_0); -- 
    ra_11387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_11388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2295_addr_3_req_1); -- 
    ca_11389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_11399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2295_load_0_req_0); -- 
    ra_11400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_11404_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_2295_load_1_req_0); -- 
    ra_11405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_11409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2295_load_2_req_0); -- 
    ra_11410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_11414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2295_load_3_req_0); -- 
    ra_11415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_11425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2295_load_0_req_1); -- 
    ca_11426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_11430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_2295_load_1_req_1); -- 
    ca_11431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_11435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2295_load_2_req_1); -- 
    ca_11436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_11440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2295_load_3_req_1); -- 
    ca_11441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_11442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_2295_gather_scatter_req_0); -- 
    merge_ack_11443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_2299_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_11453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2299_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_11464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2301_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_2307_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_11477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_11482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_2305_inst_req_0); -- 
    pipe_wack_11483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2305_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2206_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2206_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2206_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2221_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2221_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2221_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_2269 : std_logic_vector(0 downto 0);
    signal ptr_deref_2178_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2178_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2178_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2178_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2178_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2178_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2178_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2178_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2178_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2210_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2210_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2210_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2210_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2210_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2225_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2225_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2225_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2225_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2225_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2283_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2283_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2283_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2290_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2290_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2290_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2295_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2295_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2295_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2295_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2295_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2156_wire : std_logic_vector(31 downto 0);
    signal tmp10_2211 : std_logic_vector(31 downto 0);
    signal tmp11_2215 : std_logic_vector(31 downto 0);
    signal tmp12_2222 : std_logic_vector(31 downto 0);
    signal tmp13_2226 : std_logic_vector(31 downto 0);
    signal tmp14_2230 : std_logic_vector(31 downto 0);
    signal tmp15_2235 : std_logic_vector(31 downto 0);
    signal tmp16_2239 : std_logic_vector(15 downto 0);
    signal tmp17_2245 : std_logic_vector(31 downto 0);
    signal tmp18_2255 : std_logic_vector(15 downto 0);
    signal tmp19_2261 : std_logic_vector(31 downto 0);
    signal tmp1_2162 : std_logic_vector(31 downto 0);
    signal tmp20_2273 : std_logic_vector(15 downto 0);
    signal tmp21_2278 : std_logic_vector(15 downto 0);
    signal tmp22_2281 : std_logic_vector(15 downto 0);
    signal tmp23_2288 : std_logic_vector(15 downto 0);
    signal tmp24_2296 : std_logic_vector(31 downto 0);
    signal tmp25_2300 : std_logic_vector(31 downto 0);
    signal tmp2_2168 : std_logic_vector(31 downto 0);
    signal tmp3_2172 : std_logic_vector(31 downto 0);
    signal tmp4_2176 : std_logic_vector(15 downto 0);
    signal tmp5_2186 : std_logic_vector(31 downto 0);
    signal tmp6_2190 : std_logic_vector(31 downto 0);
    signal tmp7_2196 : std_logic_vector(31 downto 0);
    signal tmp8_2200 : std_logic_vector(31 downto 0);
    signal tmp9_2207 : std_logic_vector(31 downto 0);
    signal tmp_2158 : std_logic_vector(31 downto 0);
    signal type_cast_2166_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2174_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2184_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2194_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2243_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2253_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2259_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2264_wire : std_logic_vector(31 downto 0);
    signal type_cast_2267_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2307_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_2249 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2206_final_offset <= "0000000000010000";
    array_obj_ref_2221_final_offset <= "0000000000001100";
    ptr_deref_2178_word_offset_0 <= "0000000000000000";
    ptr_deref_2178_word_offset_1 <= "0000000000000001";
    ptr_deref_2210_word_offset_0 <= "0000000000000000";
    ptr_deref_2210_word_offset_1 <= "0000000000000001";
    ptr_deref_2210_word_offset_2 <= "0000000000000010";
    ptr_deref_2210_word_offset_3 <= "0000000000000011";
    ptr_deref_2225_word_offset_0 <= "0000000000000000";
    ptr_deref_2225_word_offset_1 <= "0000000000000001";
    ptr_deref_2225_word_offset_2 <= "0000000000000010";
    ptr_deref_2225_word_offset_3 <= "0000000000000011";
    ptr_deref_2283_word_offset_0 <= "0000000000000000";
    ptr_deref_2283_word_offset_1 <= "0000000000000001";
    ptr_deref_2290_word_offset_0 <= "0000000000000000";
    ptr_deref_2290_word_offset_1 <= "0000000000000001";
    ptr_deref_2295_word_offset_0 <= "0000000000000000";
    ptr_deref_2295_word_offset_1 <= "0000000000000001";
    ptr_deref_2295_word_offset_2 <= "0000000000000010";
    ptr_deref_2295_word_offset_3 <= "0000000000000011";
    type_cast_2166_wire_constant <= "11111111111111111111100000000000";
    type_cast_2174_wire_constant <= "0000000000000100";
    type_cast_2184_wire_constant <= "00000000000000000000000000000110";
    type_cast_2194_wire_constant <= "00000000000000000000000000000010";
    type_cast_2243_wire_constant <= "00000000000000000000000000000011";
    type_cast_2253_wire_constant <= "0001111111111111";
    type_cast_2259_wire_constant <= "00000000000000000000000000000111";
    type_cast_2267_wire_constant <= "00000000000000000000000000000000";
    type_cast_2303_wire_constant <= "00000000000000000000000000000011";
    array_obj_ref_2206_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2162, dout => array_obj_ref_2206_resized_base_address, req => array_obj_ref_2206_base_resize_req_0, ack => array_obj_ref_2206_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2206_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2206_root_address, dout => tmp9_2207, req => array_obj_ref_2206_final_reg_req_0, ack => array_obj_ref_2206_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2221_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2162, dout => array_obj_ref_2221_resized_base_address, req => array_obj_ref_2221_base_resize_req_0, ack => array_obj_ref_2221_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2221_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2221_root_address, dout => tmp12_2222, req => array_obj_ref_2221_final_reg_req_0, ack => array_obj_ref_2221_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2178_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2172, dout => ptr_deref_2178_resized_base_address, req => ptr_deref_2178_base_resize_req_0, ack => ptr_deref_2178_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2210_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2207, dout => ptr_deref_2210_resized_base_address, req => ptr_deref_2210_base_resize_req_0, ack => ptr_deref_2210_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2225_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2222, dout => ptr_deref_2225_resized_base_address, req => ptr_deref_2225_base_resize_req_0, ack => ptr_deref_2225_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2283_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2190, dout => ptr_deref_2283_resized_base_address, req => ptr_deref_2283_base_resize_req_0, ack => ptr_deref_2283_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2290_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2200, dout => ptr_deref_2290_resized_base_address, req => ptr_deref_2290_base_resize_req_0, ack => ptr_deref_2290_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2295_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2222, dout => ptr_deref_2295_resized_base_address, req => ptr_deref_2295_base_resize_req_0, ack => ptr_deref_2295_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2157_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2156_wire, dout => tmp_2158, req => type_cast_2157_inst_req_0, ack => type_cast_2157_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2161_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_2158, dout => tmp1_2162, req => type_cast_2161_inst_req_0, ack => type_cast_2161_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2171_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2168, dout => tmp3_2172, req => type_cast_2171_inst_req_0, ack => type_cast_2171_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2189_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2186, dout => tmp6_2190, req => type_cast_2189_inst_req_0, ack => type_cast_2189_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2199_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2196, dout => tmp8_2200, req => type_cast_2199_inst_req_0, ack => type_cast_2199_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2214_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2211, dout => tmp11_2215, req => type_cast_2214_inst_req_0, ack => type_cast_2214_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2229_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2226, dout => tmp14_2230, req => type_cast_2229_inst_req_0, ack => type_cast_2229_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2238_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_2235, dout => tmp16_2239, req => type_cast_2238_inst_req_0, ack => type_cast_2238_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2248_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_2245, dout => xx_xtrx_xi_2249, req => type_cast_2248_inst_req_0, ack => type_cast_2248_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2264_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_2261, dout => type_cast_2264_wire, req => type_cast_2264_inst_req_0, ack => type_cast_2264_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2272_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_2269, dout => tmp20_2273, req => type_cast_2272_inst_req_0, ack => type_cast_2272_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2299_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_2296, dout => tmp25_2300, req => type_cast_2299_inst_req_0, ack => type_cast_2299_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2307_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_2300, dout => type_cast_2307_wire, req => type_cast_2307_inst_req_0, ack => type_cast_2307_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2178_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2178_gather_scatter_ack_0 <= ptr_deref_2178_gather_scatter_req_0;
      aggregated_sig <= tmp4_2176;
      ptr_deref_2178_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2178_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2178_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2178_root_address_inst_ack_0 <= ptr_deref_2178_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2178_resized_base_address;
      ptr_deref_2178_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2210_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2210_gather_scatter_ack_0 <= ptr_deref_2210_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2210_data_3 & ptr_deref_2210_data_2 & ptr_deref_2210_data_1 & ptr_deref_2210_data_0;
      tmp10_2211 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2210_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2210_root_address_inst_ack_0 <= ptr_deref_2210_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2210_resized_base_address;
      ptr_deref_2210_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2225_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2225_gather_scatter_ack_0 <= ptr_deref_2225_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2225_data_3 & ptr_deref_2225_data_2 & ptr_deref_2225_data_1 & ptr_deref_2225_data_0;
      tmp13_2226 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2225_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2225_root_address_inst_ack_0 <= ptr_deref_2225_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2225_resized_base_address;
      ptr_deref_2225_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2283_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2283_gather_scatter_ack_0 <= ptr_deref_2283_gather_scatter_req_0;
      aggregated_sig <= tmp22_2281;
      ptr_deref_2283_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2283_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2283_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2283_root_address_inst_ack_0 <= ptr_deref_2283_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2283_resized_base_address;
      ptr_deref_2283_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2290_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2290_gather_scatter_ack_0 <= ptr_deref_2290_gather_scatter_req_0;
      aggregated_sig <= tmp23_2288;
      ptr_deref_2290_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2290_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2290_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2290_root_address_inst_ack_0 <= ptr_deref_2290_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2290_resized_base_address;
      ptr_deref_2290_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2295_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2295_gather_scatter_ack_0 <= ptr_deref_2295_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2295_data_3 & ptr_deref_2295_data_2 & ptr_deref_2295_data_1 & ptr_deref_2295_data_0;
      tmp24_2296 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2295_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2295_root_address_inst_ack_0 <= ptr_deref_2295_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2295_resized_base_address;
      ptr_deref_2295_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2206_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2206_resized_base_address;
      array_obj_ref_2206_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2206_root_address_inst_req_0,
          ackL => array_obj_ref_2206_root_address_inst_ack_0,
          reqR => array_obj_ref_2206_root_address_inst_req_1,
          ackR => array_obj_ref_2206_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2221_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2221_resized_base_address;
      array_obj_ref_2221_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2221_root_address_inst_req_0,
          ackL => array_obj_ref_2221_root_address_inst_ack_0,
          reqR => array_obj_ref_2221_root_address_inst_req_1,
          ackR => array_obj_ref_2221_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2167_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2158;
      tmp2_2168 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2167_inst_req_0,
          ackL => binary_2167_inst_ack_0,
          reqR => binary_2167_inst_req_1,
          ackR => binary_2167_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2185_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2168;
      tmp5_2186 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2185_inst_req_0,
          ackL => binary_2185_inst_ack_0,
          reqR => binary_2185_inst_req_1,
          ackR => binary_2185_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2195_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2168;
      tmp7_2196 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2195_inst_req_0,
          ackL => binary_2195_inst_ack_0,
          reqR => binary_2195_inst_req_1,
          ackR => binary_2195_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2234_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2215 & tmp14_2230;
      tmp15_2235 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2234_inst_req_0,
          ackL => binary_2234_inst_ack_0,
          reqR => binary_2234_inst_req_1,
          ackR => binary_2234_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2244_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2235;
      tmp17_2245 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2244_inst_req_0,
          ackL => binary_2244_inst_ack_0,
          reqR => binary_2244_inst_req_1,
          ackR => binary_2244_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2254_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_2249;
      tmp18_2255 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2254_inst_req_0,
          ackL => binary_2254_inst_ack_0,
          reqR => binary_2254_inst_req_1,
          ackR => binary_2254_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2260_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2235;
      tmp19_2261 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2260_inst_req_0,
          ackL => binary_2260_inst_ack_0,
          reqR => binary_2260_inst_req_1,
          ackR => binary_2260_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2268_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2264_wire;
      notx_xx_xi_2269 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2268_inst_req_0,
          ackL => binary_2268_inst_ack_0,
          reqR => binary_2268_inst_req_1,
          ackR => binary_2268_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2277_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_2255 & tmp20_2273;
      tmp21_2278 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2277_inst_req_0,
          ackL => binary_2277_inst_ack_0,
          reqR => binary_2277_inst_req_1,
          ackR => binary_2277_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2178_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2178_root_address;
      ptr_deref_2178_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2178_addr_0_req_0,
          ackL => ptr_deref_2178_addr_0_ack_0,
          reqR => ptr_deref_2178_addr_0_req_1,
          ackR => ptr_deref_2178_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2178_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2178_root_address;
      ptr_deref_2178_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2178_addr_1_req_0,
          ackL => ptr_deref_2178_addr_1_ack_0,
          reqR => ptr_deref_2178_addr_1_req_1,
          ackR => ptr_deref_2178_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2210_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2210_root_address;
      ptr_deref_2210_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2210_addr_0_req_0,
          ackL => ptr_deref_2210_addr_0_ack_0,
          reqR => ptr_deref_2210_addr_0_req_1,
          ackR => ptr_deref_2210_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2210_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2210_root_address;
      ptr_deref_2210_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2210_addr_1_req_0,
          ackL => ptr_deref_2210_addr_1_ack_0,
          reqR => ptr_deref_2210_addr_1_req_1,
          ackR => ptr_deref_2210_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2210_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2210_root_address;
      ptr_deref_2210_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2210_addr_2_req_0,
          ackL => ptr_deref_2210_addr_2_ack_0,
          reqR => ptr_deref_2210_addr_2_req_1,
          ackR => ptr_deref_2210_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2210_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2210_root_address;
      ptr_deref_2210_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2210_addr_3_req_0,
          ackL => ptr_deref_2210_addr_3_ack_0,
          reqR => ptr_deref_2210_addr_3_req_1,
          ackR => ptr_deref_2210_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2225_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2225_root_address;
      ptr_deref_2225_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2225_addr_0_req_0,
          ackL => ptr_deref_2225_addr_0_ack_0,
          reqR => ptr_deref_2225_addr_0_req_1,
          ackR => ptr_deref_2225_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2225_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2225_root_address;
      ptr_deref_2225_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2225_addr_1_req_0,
          ackL => ptr_deref_2225_addr_1_ack_0,
          reqR => ptr_deref_2225_addr_1_req_1,
          ackR => ptr_deref_2225_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2225_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2225_root_address;
      ptr_deref_2225_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2225_addr_2_req_0,
          ackL => ptr_deref_2225_addr_2_ack_0,
          reqR => ptr_deref_2225_addr_2_req_1,
          ackR => ptr_deref_2225_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2225_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2225_root_address;
      ptr_deref_2225_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2225_addr_3_req_0,
          ackL => ptr_deref_2225_addr_3_ack_0,
          reqR => ptr_deref_2225_addr_3_req_1,
          ackR => ptr_deref_2225_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2283_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2283_root_address;
      ptr_deref_2283_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2283_addr_0_req_0,
          ackL => ptr_deref_2283_addr_0_ack_0,
          reqR => ptr_deref_2283_addr_0_req_1,
          ackR => ptr_deref_2283_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2283_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2283_root_address;
      ptr_deref_2283_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2283_addr_1_req_0,
          ackL => ptr_deref_2283_addr_1_ack_0,
          reqR => ptr_deref_2283_addr_1_req_1,
          ackR => ptr_deref_2283_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2290_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2290_root_address;
      ptr_deref_2290_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2290_addr_0_req_0,
          ackL => ptr_deref_2290_addr_0_ack_0,
          reqR => ptr_deref_2290_addr_0_req_1,
          ackR => ptr_deref_2290_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2290_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2290_root_address;
      ptr_deref_2290_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2290_addr_1_req_0,
          ackL => ptr_deref_2290_addr_1_ack_0,
          reqR => ptr_deref_2290_addr_1_req_1,
          ackR => ptr_deref_2290_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2295_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2295_root_address;
      ptr_deref_2295_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2295_addr_0_req_0,
          ackL => ptr_deref_2295_addr_0_ack_0,
          reqR => ptr_deref_2295_addr_0_req_1,
          ackR => ptr_deref_2295_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2295_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2295_root_address;
      ptr_deref_2295_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2295_addr_1_req_0,
          ackL => ptr_deref_2295_addr_1_ack_0,
          reqR => ptr_deref_2295_addr_1_req_1,
          ackR => ptr_deref_2295_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2295_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2295_root_address;
      ptr_deref_2295_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2295_addr_2_req_0,
          ackL => ptr_deref_2295_addr_2_ack_0,
          reqR => ptr_deref_2295_addr_2_req_1,
          ackR => ptr_deref_2295_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2295_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2295_root_address;
      ptr_deref_2295_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2295_addr_3_req_0,
          ackL => ptr_deref_2295_addr_3_ack_0,
          reqR => ptr_deref_2295_addr_3_req_1,
          ackR => ptr_deref_2295_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2210_load_0 ptr_deref_2210_load_1 ptr_deref_2210_load_2 ptr_deref_2210_load_3 ptr_deref_2225_load_0 ptr_deref_2225_load_1 ptr_deref_2225_load_2 ptr_deref_2225_load_3 ptr_deref_2295_load_0 ptr_deref_2295_load_1 ptr_deref_2295_load_2 ptr_deref_2295_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2210_load_0_req_0,
        ptr_deref_2210_load_0_ack_0,
        ptr_deref_2210_load_0_req_1,
        ptr_deref_2210_load_0_ack_1,
        "ptr_deref_2210_load_0",
        "memory_space_5" ,
        ptr_deref_2210_data_0,
        ptr_deref_2210_word_address_0,
        "ptr_deref_2210_data_0",
        "ptr_deref_2210_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2210_load_1_req_0,
        ptr_deref_2210_load_1_ack_0,
        ptr_deref_2210_load_1_req_1,
        ptr_deref_2210_load_1_ack_1,
        "ptr_deref_2210_load_1",
        "memory_space_5" ,
        ptr_deref_2210_data_1,
        ptr_deref_2210_word_address_1,
        "ptr_deref_2210_data_1",
        "ptr_deref_2210_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2210_load_2_req_0,
        ptr_deref_2210_load_2_ack_0,
        ptr_deref_2210_load_2_req_1,
        ptr_deref_2210_load_2_ack_1,
        "ptr_deref_2210_load_2",
        "memory_space_5" ,
        ptr_deref_2210_data_2,
        ptr_deref_2210_word_address_2,
        "ptr_deref_2210_data_2",
        "ptr_deref_2210_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2210_load_3_req_0,
        ptr_deref_2210_load_3_ack_0,
        ptr_deref_2210_load_3_req_1,
        ptr_deref_2210_load_3_ack_1,
        "ptr_deref_2210_load_3",
        "memory_space_5" ,
        ptr_deref_2210_data_3,
        ptr_deref_2210_word_address_3,
        "ptr_deref_2210_data_3",
        "ptr_deref_2210_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2225_load_0_req_0,
        ptr_deref_2225_load_0_ack_0,
        ptr_deref_2225_load_0_req_1,
        ptr_deref_2225_load_0_ack_1,
        "ptr_deref_2225_load_0",
        "memory_space_5" ,
        ptr_deref_2225_data_0,
        ptr_deref_2225_word_address_0,
        "ptr_deref_2225_data_0",
        "ptr_deref_2225_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2225_load_1_req_0,
        ptr_deref_2225_load_1_ack_0,
        ptr_deref_2225_load_1_req_1,
        ptr_deref_2225_load_1_ack_1,
        "ptr_deref_2225_load_1",
        "memory_space_5" ,
        ptr_deref_2225_data_1,
        ptr_deref_2225_word_address_1,
        "ptr_deref_2225_data_1",
        "ptr_deref_2225_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2225_load_2_req_0,
        ptr_deref_2225_load_2_ack_0,
        ptr_deref_2225_load_2_req_1,
        ptr_deref_2225_load_2_ack_1,
        "ptr_deref_2225_load_2",
        "memory_space_5" ,
        ptr_deref_2225_data_2,
        ptr_deref_2225_word_address_2,
        "ptr_deref_2225_data_2",
        "ptr_deref_2225_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2225_load_3_req_0,
        ptr_deref_2225_load_3_ack_0,
        ptr_deref_2225_load_3_req_1,
        ptr_deref_2225_load_3_ack_1,
        "ptr_deref_2225_load_3",
        "memory_space_5" ,
        ptr_deref_2225_data_3,
        ptr_deref_2225_word_address_3,
        "ptr_deref_2225_data_3",
        "ptr_deref_2225_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2295_load_0_req_0,
        ptr_deref_2295_load_0_ack_0,
        ptr_deref_2295_load_0_req_1,
        ptr_deref_2295_load_0_ack_1,
        "ptr_deref_2295_load_0",
        "memory_space_5" ,
        ptr_deref_2295_data_0,
        ptr_deref_2295_word_address_0,
        "ptr_deref_2295_data_0",
        "ptr_deref_2295_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2295_load_1_req_0,
        ptr_deref_2295_load_1_ack_0,
        ptr_deref_2295_load_1_req_1,
        ptr_deref_2295_load_1_ack_1,
        "ptr_deref_2295_load_1",
        "memory_space_5" ,
        ptr_deref_2295_data_1,
        ptr_deref_2295_word_address_1,
        "ptr_deref_2295_data_1",
        "ptr_deref_2295_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2295_load_2_req_0,
        ptr_deref_2295_load_2_ack_0,
        ptr_deref_2295_load_2_req_1,
        ptr_deref_2295_load_2_ack_1,
        "ptr_deref_2295_load_2",
        "memory_space_5" ,
        ptr_deref_2295_data_2,
        ptr_deref_2295_word_address_2,
        "ptr_deref_2295_data_2",
        "ptr_deref_2295_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2295_load_3_req_0,
        ptr_deref_2295_load_3_ack_0,
        ptr_deref_2295_load_3_req_1,
        ptr_deref_2295_load_3_ack_1,
        "ptr_deref_2295_load_3",
        "memory_space_5" ,
        ptr_deref_2295_data_3,
        ptr_deref_2295_word_address_3,
        "ptr_deref_2295_data_3",
        "ptr_deref_2295_word_address_3" -- 
      );
      reqL(11) <= ptr_deref_2210_load_0_req_0;
      reqL(10) <= ptr_deref_2210_load_1_req_0;
      reqL(9) <= ptr_deref_2210_load_2_req_0;
      reqL(8) <= ptr_deref_2210_load_3_req_0;
      reqL(7) <= ptr_deref_2225_load_0_req_0;
      reqL(6) <= ptr_deref_2225_load_1_req_0;
      reqL(5) <= ptr_deref_2225_load_2_req_0;
      reqL(4) <= ptr_deref_2225_load_3_req_0;
      reqL(3) <= ptr_deref_2295_load_0_req_0;
      reqL(2) <= ptr_deref_2295_load_1_req_0;
      reqL(1) <= ptr_deref_2295_load_2_req_0;
      reqL(0) <= ptr_deref_2295_load_3_req_0;
      ptr_deref_2210_load_0_ack_0 <= ackL(11);
      ptr_deref_2210_load_1_ack_0 <= ackL(10);
      ptr_deref_2210_load_2_ack_0 <= ackL(9);
      ptr_deref_2210_load_3_ack_0 <= ackL(8);
      ptr_deref_2225_load_0_ack_0 <= ackL(7);
      ptr_deref_2225_load_1_ack_0 <= ackL(6);
      ptr_deref_2225_load_2_ack_0 <= ackL(5);
      ptr_deref_2225_load_3_ack_0 <= ackL(4);
      ptr_deref_2295_load_0_ack_0 <= ackL(3);
      ptr_deref_2295_load_1_ack_0 <= ackL(2);
      ptr_deref_2295_load_2_ack_0 <= ackL(1);
      ptr_deref_2295_load_3_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2210_load_0_req_1;
      reqR(10) <= ptr_deref_2210_load_1_req_1;
      reqR(9) <= ptr_deref_2210_load_2_req_1;
      reqR(8) <= ptr_deref_2210_load_3_req_1;
      reqR(7) <= ptr_deref_2225_load_0_req_1;
      reqR(6) <= ptr_deref_2225_load_1_req_1;
      reqR(5) <= ptr_deref_2225_load_2_req_1;
      reqR(4) <= ptr_deref_2225_load_3_req_1;
      reqR(3) <= ptr_deref_2295_load_0_req_1;
      reqR(2) <= ptr_deref_2295_load_1_req_1;
      reqR(1) <= ptr_deref_2295_load_2_req_1;
      reqR(0) <= ptr_deref_2295_load_3_req_1;
      ptr_deref_2210_load_0_ack_1 <= ackR(11);
      ptr_deref_2210_load_1_ack_1 <= ackR(10);
      ptr_deref_2210_load_2_ack_1 <= ackR(9);
      ptr_deref_2210_load_3_ack_1 <= ackR(8);
      ptr_deref_2225_load_0_ack_1 <= ackR(7);
      ptr_deref_2225_load_1_ack_1 <= ackR(6);
      ptr_deref_2225_load_2_ack_1 <= ackR(5);
      ptr_deref_2225_load_3_ack_1 <= ackR(4);
      ptr_deref_2295_load_0_ack_1 <= ackR(3);
      ptr_deref_2295_load_1_ack_1 <= ackR(2);
      ptr_deref_2295_load_2_ack_1 <= ackR(1);
      ptr_deref_2295_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_2210_word_address_0 & ptr_deref_2210_word_address_1 & ptr_deref_2210_word_address_2 & ptr_deref_2210_word_address_3 & ptr_deref_2225_word_address_0 & ptr_deref_2225_word_address_1 & ptr_deref_2225_word_address_2 & ptr_deref_2225_word_address_3 & ptr_deref_2295_word_address_0 & ptr_deref_2295_word_address_1 & ptr_deref_2295_word_address_2 & ptr_deref_2295_word_address_3;
      ptr_deref_2210_data_0 <= data_out(95 downto 88);
      ptr_deref_2210_data_1 <= data_out(87 downto 80);
      ptr_deref_2210_data_2 <= data_out(79 downto 72);
      ptr_deref_2210_data_3 <= data_out(71 downto 64);
      ptr_deref_2225_data_0 <= data_out(63 downto 56);
      ptr_deref_2225_data_1 <= data_out(55 downto 48);
      ptr_deref_2225_data_2 <= data_out(47 downto 40);
      ptr_deref_2225_data_3 <= data_out(39 downto 32);
      ptr_deref_2295_data_0 <= data_out(31 downto 24);
      ptr_deref_2295_data_1 <= data_out(23 downto 16);
      ptr_deref_2295_data_2 <= data_out(15 downto 8);
      ptr_deref_2295_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2178_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2178_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2178_word_address_0) &  " data ptr_deref_2178_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2178_data_0) severity note; --
        end if;
        if ptr_deref_2178_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2178_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2178_word_address_1) &  " data ptr_deref_2178_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2178_data_1) severity note; --
        end if;
        if ptr_deref_2283_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2283_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2283_word_address_0) &  " data ptr_deref_2283_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2283_data_0) severity note; --
        end if;
        if ptr_deref_2283_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2283_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2283_word_address_1) &  " data ptr_deref_2283_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2283_data_1) severity note; --
        end if;
        if ptr_deref_2290_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2290_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2290_word_address_0) &  " data ptr_deref_2290_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2290_data_0) severity note; --
        end if;
        if ptr_deref_2290_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2290_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2290_word_address_1) &  " data ptr_deref_2290_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2290_data_1) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2178_store_0 ptr_deref_2178_store_1 ptr_deref_2283_store_0 ptr_deref_2283_store_1 ptr_deref_2290_store_0 ptr_deref_2290_store_1 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2178_store_0_req_0;
      reqL(4) <= ptr_deref_2178_store_1_req_0;
      reqL(3) <= ptr_deref_2283_store_0_req_0;
      reqL(2) <= ptr_deref_2283_store_1_req_0;
      reqL(1) <= ptr_deref_2290_store_0_req_0;
      reqL(0) <= ptr_deref_2290_store_1_req_0;
      ptr_deref_2178_store_0_ack_0 <= ackL(5);
      ptr_deref_2178_store_1_ack_0 <= ackL(4);
      ptr_deref_2283_store_0_ack_0 <= ackL(3);
      ptr_deref_2283_store_1_ack_0 <= ackL(2);
      ptr_deref_2290_store_0_ack_0 <= ackL(1);
      ptr_deref_2290_store_1_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2178_store_0_req_1;
      reqR(4) <= ptr_deref_2178_store_1_req_1;
      reqR(3) <= ptr_deref_2283_store_0_req_1;
      reqR(2) <= ptr_deref_2283_store_1_req_1;
      reqR(1) <= ptr_deref_2290_store_0_req_1;
      reqR(0) <= ptr_deref_2290_store_1_req_1;
      ptr_deref_2178_store_0_ack_1 <= ackR(5);
      ptr_deref_2178_store_1_ack_1 <= ackR(4);
      ptr_deref_2283_store_0_ack_1 <= ackR(3);
      ptr_deref_2283_store_1_ack_1 <= ackR(2);
      ptr_deref_2290_store_0_ack_1 <= ackR(1);
      ptr_deref_2290_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2178_word_address_0 & ptr_deref_2178_word_address_1 & ptr_deref_2283_word_address_0 & ptr_deref_2283_word_address_1 & ptr_deref_2290_word_address_0 & ptr_deref_2290_word_address_1;
      data_in <= ptr_deref_2178_data_0 & ptr_deref_2178_data_1 & ptr_deref_2283_data_0 & ptr_deref_2283_data_1 & ptr_deref_2290_data_0 & ptr_deref_2290_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2156_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2156_inst_ack_0 then -- 
            assert false report " ReadPipe to2_in0 to wire simple_obj_ref_2156_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2156_inst_req_0;
      simple_obj_ref_2156_inst_ack_0 <= ack(0);
      simple_obj_ref_2156_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to2_in0_pipe_read_req(0),
          oack => to2_in0_pipe_read_ack(0),
          odata => to2_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2301_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_2303_wire_constant value="  &  convert_slv_to_hex_string(type_cast_2303_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2301_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2301_inst_req_0;
      simple_obj_ref_2301_inst_ack_0 <= ack(0);
      data_in <= type_cast_2303_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2305_inst_ack_0 then -- 
          assert false report " WritePipe tofpga2_out0 from wire type_cast_2307_wire value="  &  convert_slv_to_hex_string(type_cast_2307_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2305_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2305_inst_req_0;
      simple_obj_ref_2305_inst_ack_0 <= ack(0);
      data_in <= type_cast_2307_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga2_out0_pipe_write_req(0),
          oack => tofpga2_out0_pipe_write_ack(0),
          odata => tofpga2_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2176_call call_stmt_2281_call call_stmt_2288_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2176_call_req_0;
      reqL(1) <= call_stmt_2281_call_req_0;
      reqL(0) <= call_stmt_2288_call_req_0;
      call_stmt_2176_call_ack_0 <= ackL(2);
      call_stmt_2281_call_ack_0 <= ackL(1);
      call_stmt_2288_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2176_call_req_1;
      reqR(1) <= call_stmt_2281_call_req_1;
      reqR(0) <= call_stmt_2288_call_req_1;
      call_stmt_2176_call_ack_1 <= ackR(2);
      call_stmt_2281_call_ack_1 <= ackR(1);
      call_stmt_2288_call_ack_1 <= ackR(0);
      data_in <= type_cast_2174_wire_constant & tmp16_2239 & tmp21_2278;
      tmp4_2176 <= data_out(47 downto 32);
      tmp22_2281 <= data_out(31 downto 16);
      tmp23_2288 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to3 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to3_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to3_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to3_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga3_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to3;
architecture Default of ahir_glue_to3 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to3_CP_11492_start: Boolean;
  -- links between control-path and data-path
  signal type_cast_2408_inst_ack_0 : boolean;
  signal ptr_deref_2455_addr_2_ack_0 : boolean;
  signal call_stmt_2441_call_req_0 : boolean;
  signal array_obj_ref_2381_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2455_root_address_inst_req_0 : boolean;
  signal type_cast_2432_inst_req_0 : boolean;
  signal array_obj_ref_2381_root_address_inst_req_0 : boolean;
  signal ptr_deref_2443_store_1_ack_1 : boolean;
  signal binary_2414_inst_req_0 : boolean;
  signal ptr_deref_2443_store_1_req_1 : boolean;
  signal ptr_deref_2443_addr_0_ack_1 : boolean;
  signal array_obj_ref_2381_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2455_load_3_req_0 : boolean;
  signal ptr_deref_2385_load_1_req_1 : boolean;
  signal binary_2404_inst_ack_0 : boolean;
  signal call_stmt_2441_call_ack_1 : boolean;
  signal ptr_deref_2385_addr_2_ack_0 : boolean;
  signal ptr_deref_2450_gather_scatter_req_0 : boolean;
  signal ptr_deref_2443_store_0_ack_1 : boolean;
  signal ptr_deref_2455_addr_0_req_1 : boolean;
  signal array_obj_ref_2381_base_resize_req_0 : boolean;
  signal ptr_deref_2455_addr_2_req_1 : boolean;
  signal ptr_deref_2455_addr_1_ack_0 : boolean;
  signal ptr_deref_2385_load_2_req_1 : boolean;
  signal ptr_deref_2385_addr_3_req_0 : boolean;
  signal ptr_deref_2455_load_3_ack_1 : boolean;
  signal binary_2414_inst_ack_0 : boolean;
  signal ptr_deref_2455_addr_0_ack_1 : boolean;
  signal type_cast_2408_inst_req_0 : boolean;
  signal ptr_deref_2450_addr_0_ack_0 : boolean;
  signal ptr_deref_2450_addr_0_ack_1 : boolean;
  signal ptr_deref_2455_addr_0_ack_0 : boolean;
  signal ptr_deref_2450_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2443_store_0_req_1 : boolean;
  signal call_stmt_2441_call_ack_0 : boolean;
  signal binary_2404_inst_req_0 : boolean;
  signal array_obj_ref_2381_base_resize_ack_0 : boolean;
  signal ptr_deref_2455_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2443_addr_0_ack_0 : boolean;
  signal ptr_deref_2385_load_3_req_0 : boolean;
  signal ptr_deref_2450_store_0_ack_1 : boolean;
  signal ptr_deref_2455_load_1_req_0 : boolean;
  signal ptr_deref_2443_store_1_ack_0 : boolean;
  signal type_cast_2432_inst_ack_0 : boolean;
  signal ptr_deref_2455_load_0_ack_0 : boolean;
  signal ptr_deref_2385_load_0_req_1 : boolean;
  signal ptr_deref_2450_addr_0_req_1 : boolean;
  signal ptr_deref_2443_store_0_req_0 : boolean;
  signal binary_2414_inst_ack_1 : boolean;
  signal ptr_deref_2443_store_0_ack_0 : boolean;
  signal ptr_deref_2455_load_1_ack_0 : boolean;
  signal ptr_deref_2450_store_0_req_1 : boolean;
  signal ptr_deref_2450_root_address_inst_req_0 : boolean;
  signal ptr_deref_2443_addr_0_req_1 : boolean;
  signal binary_2404_inst_req_1 : boolean;
  signal ptr_deref_2450_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2443_store_1_req_0 : boolean;
  signal binary_2414_inst_req_1 : boolean;
  signal binary_2404_inst_ack_1 : boolean;
  signal array_obj_ref_2381_root_address_inst_req_1 : boolean;
  signal ptr_deref_2385_addr_2_ack_1 : boolean;
  signal ptr_deref_2455_addr_1_req_0 : boolean;
  signal ptr_deref_2385_load_2_ack_0 : boolean;
  signal ptr_deref_2385_load_1_ack_1 : boolean;
  signal ptr_deref_2455_load_2_req_0 : boolean;
  signal array_obj_ref_2381_final_reg_req_0 : boolean;
  signal array_obj_ref_2381_final_reg_ack_0 : boolean;
  signal ptr_deref_2455_load_3_req_1 : boolean;
  signal ptr_deref_2385_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2385_load_2_ack_1 : boolean;
  signal ptr_deref_2385_base_resize_req_0 : boolean;
  signal ptr_deref_2385_load_3_ack_0 : boolean;
  signal call_stmt_2441_call_req_1 : boolean;
  signal binary_2437_inst_ack_0 : boolean;
  signal ptr_deref_2455_addr_0_req_0 : boolean;
  signal ptr_deref_2450_base_resize_ack_0 : boolean;
  signal binary_2437_inst_req_0 : boolean;
  signal ptr_deref_2385_addr_2_req_1 : boolean;
  signal ptr_deref_2385_load_0_ack_1 : boolean;
  signal binary_2437_inst_req_1 : boolean;
  signal ptr_deref_2450_addr_1_req_1 : boolean;
  signal ptr_deref_2450_base_resize_req_0 : boolean;
  signal ptr_deref_2385_addr_2_req_0 : boolean;
  signal binary_2437_inst_ack_1 : boolean;
  signal ptr_deref_2385_load_2_req_0 : boolean;
  signal ptr_deref_2455_addr_1_ack_1 : boolean;
  signal ptr_deref_2450_addr_0_req_0 : boolean;
  signal ptr_deref_2455_load_2_req_1 : boolean;
  signal ptr_deref_2455_addr_3_ack_1 : boolean;
  signal ptr_deref_2455_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_2461_inst_ack_0 : boolean;
  signal ptr_deref_2443_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2443_gather_scatter_ack_0 : boolean;
  signal type_cast_2398_inst_ack_0 : boolean;
  signal type_cast_2398_inst_req_0 : boolean;
  signal ptr_deref_2443_gather_scatter_req_0 : boolean;
  signal ptr_deref_2450_store_1_ack_1 : boolean;
  signal type_cast_2389_inst_ack_0 : boolean;
  signal ptr_deref_2443_addr_0_req_0 : boolean;
  signal ptr_deref_2385_addr_1_ack_1 : boolean;
  signal ptr_deref_2385_addr_1_req_1 : boolean;
  signal type_cast_2374_inst_ack_0 : boolean;
  signal ptr_deref_2385_addr_1_ack_0 : boolean;
  signal ptr_deref_2385_addr_1_req_0 : boolean;
  signal ptr_deref_2385_load_1_ack_0 : boolean;
  signal type_cast_2374_inst_req_0 : boolean;
  signal ptr_deref_2450_store_1_req_1 : boolean;
  signal ptr_deref_2385_load_1_req_0 : boolean;
  signal ptr_deref_2443_addr_1_ack_1 : boolean;
  signal ptr_deref_2443_addr_1_req_1 : boolean;
  signal binary_2394_inst_ack_1 : boolean;
  signal ptr_deref_2455_addr_2_req_0 : boolean;
  signal binary_2394_inst_req_1 : boolean;
  signal ptr_deref_2443_addr_1_ack_0 : boolean;
  signal binary_2394_inst_ack_0 : boolean;
  signal binary_2394_inst_req_0 : boolean;
  signal ptr_deref_2450_addr_1_ack_1 : boolean;
  signal ptr_deref_2385_base_resize_ack_0 : boolean;
  signal call_stmt_2448_call_req_0 : boolean;
  signal call_stmt_2448_call_ack_0 : boolean;
  signal ptr_deref_2455_addr_2_ack_1 : boolean;
  signal ptr_deref_2385_load_3_req_1 : boolean;
  signal call_stmt_2448_call_req_1 : boolean;
  signal binary_2420_inst_req_0 : boolean;
  signal binary_2420_inst_ack_0 : boolean;
  signal binary_2420_inst_req_1 : boolean;
  signal call_stmt_2448_call_ack_1 : boolean;
  signal ptr_deref_2443_addr_1_req_0 : boolean;
  signal ptr_deref_2385_root_address_inst_req_0 : boolean;
  signal binary_2420_inst_ack_1 : boolean;
  signal type_cast_2467_inst_req_0 : boolean;
  signal ptr_deref_2385_load_3_ack_1 : boolean;
  signal ptr_deref_2450_addr_1_req_0 : boolean;
  signal ptr_deref_2450_store_0_req_0 : boolean;
  signal simple_obj_ref_2465_inst_req_0 : boolean;
  signal type_cast_2459_inst_req_0 : boolean;
  signal ptr_deref_2385_gather_scatter_req_0 : boolean;
  signal ptr_deref_2455_base_resize_req_0 : boolean;
  signal type_cast_2389_inst_req_0 : boolean;
  signal ptr_deref_2455_load_1_req_1 : boolean;
  signal ptr_deref_2450_addr_1_ack_0 : boolean;
  signal simple_obj_ref_2465_inst_ack_0 : boolean;
  signal ptr_deref_2385_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2450_store_0_ack_0 : boolean;
  signal ptr_deref_2443_base_resize_req_0 : boolean;
  signal ptr_deref_2455_load_1_ack_1 : boolean;
  signal ptr_deref_2455_load_2_ack_0 : boolean;
  signal ptr_deref_2443_base_resize_ack_0 : boolean;
  signal ptr_deref_2455_gather_scatter_req_0 : boolean;
  signal type_cast_2467_inst_ack_0 : boolean;
  signal ptr_deref_2455_addr_1_req_1 : boolean;
  signal ptr_deref_2385_addr_0_req_0 : boolean;
  signal ptr_deref_2455_addr_3_req_0 : boolean;
  signal ptr_deref_2455_load_0_req_1 : boolean;
  signal type_cast_2424_inst_req_0 : boolean;
  signal type_cast_2424_inst_ack_0 : boolean;
  signal ptr_deref_2455_load_0_ack_1 : boolean;
  signal type_cast_2459_inst_ack_0 : boolean;
  signal ptr_deref_2385_addr_0_ack_0 : boolean;
  signal ptr_deref_2385_addr_0_req_1 : boolean;
  signal ptr_deref_2450_store_1_req_0 : boolean;
  signal ptr_deref_2385_addr_0_ack_1 : boolean;
  signal ptr_deref_2450_store_1_ack_0 : boolean;
  signal ptr_deref_2443_root_address_inst_req_0 : boolean;
  signal binary_2428_inst_req_0 : boolean;
  signal binary_2428_inst_ack_0 : boolean;
  signal binary_2428_inst_req_1 : boolean;
  signal ptr_deref_2455_addr_3_ack_0 : boolean;
  signal ptr_deref_2455_base_resize_ack_0 : boolean;
  signal simple_obj_ref_2461_inst_req_0 : boolean;
  signal binary_2428_inst_ack_1 : boolean;
  signal simple_obj_ref_2316_inst_req_0 : boolean;
  signal simple_obj_ref_2316_inst_ack_0 : boolean;
  signal type_cast_2317_inst_req_0 : boolean;
  signal type_cast_2317_inst_ack_0 : boolean;
  signal type_cast_2321_inst_req_0 : boolean;
  signal type_cast_2321_inst_ack_0 : boolean;
  signal binary_2327_inst_req_0 : boolean;
  signal binary_2327_inst_ack_0 : boolean;
  signal binary_2327_inst_req_1 : boolean;
  signal binary_2327_inst_ack_1 : boolean;
  signal type_cast_2331_inst_req_0 : boolean;
  signal type_cast_2331_inst_ack_0 : boolean;
  signal call_stmt_2336_call_req_0 : boolean;
  signal call_stmt_2336_call_ack_0 : boolean;
  signal call_stmt_2336_call_req_1 : boolean;
  signal call_stmt_2336_call_ack_1 : boolean;
  signal ptr_deref_2338_base_resize_req_0 : boolean;
  signal ptr_deref_2338_base_resize_ack_0 : boolean;
  signal ptr_deref_2338_root_address_inst_req_0 : boolean;
  signal ptr_deref_2338_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2385_addr_3_ack_1 : boolean;
  signal ptr_deref_2338_addr_0_req_0 : boolean;
  signal ptr_deref_2338_addr_0_ack_0 : boolean;
  signal ptr_deref_2338_addr_0_req_1 : boolean;
  signal ptr_deref_2338_addr_0_ack_1 : boolean;
  signal ptr_deref_2338_addr_1_req_0 : boolean;
  signal ptr_deref_2338_addr_1_ack_0 : boolean;
  signal ptr_deref_2338_addr_1_req_1 : boolean;
  signal ptr_deref_2338_addr_1_ack_1 : boolean;
  signal ptr_deref_2385_addr_3_req_1 : boolean;
  signal ptr_deref_2385_addr_3_ack_0 : boolean;
  signal ptr_deref_2338_gather_scatter_req_0 : boolean;
  signal ptr_deref_2338_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2338_store_0_req_0 : boolean;
  signal ptr_deref_2338_store_0_ack_0 : boolean;
  signal ptr_deref_2338_store_1_req_0 : boolean;
  signal ptr_deref_2338_store_1_ack_0 : boolean;
  signal ptr_deref_2338_store_0_req_1 : boolean;
  signal ptr_deref_2338_store_0_ack_1 : boolean;
  signal ptr_deref_2338_store_1_req_1 : boolean;
  signal ptr_deref_2338_store_1_ack_1 : boolean;
  signal ptr_deref_2455_load_3_ack_0 : boolean;
  signal ptr_deref_2455_addr_3_req_1 : boolean;
  signal ptr_deref_2455_load_0_req_0 : boolean;
  signal binary_2345_inst_req_0 : boolean;
  signal binary_2345_inst_ack_0 : boolean;
  signal binary_2345_inst_req_1 : boolean;
  signal binary_2345_inst_ack_1 : boolean;
  signal ptr_deref_2455_load_2_ack_1 : boolean;
  signal ptr_deref_2385_load_0_ack_0 : boolean;
  signal ptr_deref_2385_load_0_req_0 : boolean;
  signal type_cast_2349_inst_req_0 : boolean;
  signal type_cast_2349_inst_ack_0 : boolean;
  signal binary_2355_inst_req_0 : boolean;
  signal binary_2355_inst_ack_0 : boolean;
  signal binary_2355_inst_req_1 : boolean;
  signal binary_2355_inst_ack_1 : boolean;
  signal type_cast_2359_inst_req_0 : boolean;
  signal type_cast_2359_inst_ack_0 : boolean;
  signal array_obj_ref_2366_base_resize_req_0 : boolean;
  signal array_obj_ref_2366_base_resize_ack_0 : boolean;
  signal array_obj_ref_2366_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2366_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2366_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2366_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2366_final_reg_req_0 : boolean;
  signal array_obj_ref_2366_final_reg_ack_0 : boolean;
  signal ptr_deref_2370_base_resize_req_0 : boolean;
  signal ptr_deref_2370_base_resize_ack_0 : boolean;
  signal ptr_deref_2370_root_address_inst_req_0 : boolean;
  signal ptr_deref_2370_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2370_addr_0_req_0 : boolean;
  signal ptr_deref_2370_addr_0_ack_0 : boolean;
  signal ptr_deref_2370_addr_0_req_1 : boolean;
  signal ptr_deref_2370_addr_0_ack_1 : boolean;
  signal ptr_deref_2370_addr_1_req_0 : boolean;
  signal ptr_deref_2370_addr_1_ack_0 : boolean;
  signal ptr_deref_2370_addr_1_req_1 : boolean;
  signal ptr_deref_2370_addr_1_ack_1 : boolean;
  signal ptr_deref_2370_addr_2_req_0 : boolean;
  signal ptr_deref_2370_addr_2_ack_0 : boolean;
  signal ptr_deref_2370_addr_2_req_1 : boolean;
  signal ptr_deref_2370_addr_2_ack_1 : boolean;
  signal ptr_deref_2370_addr_3_req_0 : boolean;
  signal ptr_deref_2370_addr_3_ack_0 : boolean;
  signal ptr_deref_2370_addr_3_req_1 : boolean;
  signal ptr_deref_2370_addr_3_ack_1 : boolean;
  signal ptr_deref_2370_load_0_req_0 : boolean;
  signal ptr_deref_2370_load_0_ack_0 : boolean;
  signal ptr_deref_2370_load_1_req_0 : boolean;
  signal ptr_deref_2370_load_1_ack_0 : boolean;
  signal ptr_deref_2370_load_2_req_0 : boolean;
  signal ptr_deref_2370_load_2_ack_0 : boolean;
  signal ptr_deref_2370_load_3_req_0 : boolean;
  signal ptr_deref_2370_load_3_ack_0 : boolean;
  signal ptr_deref_2370_load_0_req_1 : boolean;
  signal ptr_deref_2370_load_0_ack_1 : boolean;
  signal ptr_deref_2370_load_1_req_1 : boolean;
  signal ptr_deref_2370_load_1_ack_1 : boolean;
  signal ptr_deref_2370_load_2_req_1 : boolean;
  signal ptr_deref_2370_load_2_ack_1 : boolean;
  signal ptr_deref_2370_load_3_req_1 : boolean;
  signal ptr_deref_2370_load_3_ack_1 : boolean;
  signal ptr_deref_2370_gather_scatter_req_0 : boolean;
  signal ptr_deref_2370_gather_scatter_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to3_CP_11492: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_11583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2336_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_12108_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2441_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_12406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2461_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_2317_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_11533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_2316_inst_req_0); -- 
    ack_11534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2316_inst_ack_0, ack => cp_elements(8)); -- 
    ack_11539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2317_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2321_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_11552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2321_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2327_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_11562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2327_inst_ack_0, ack => cp_elements(18)); -- 
    cr_11563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2327_inst_req_1); -- 
    ca_11564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2327_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2331_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_11574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_11584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2336_call_ack_0, ack => cp_elements(24)); -- 
    ccr_11588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2336_call_req_1); -- 
    cca_11589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2336_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2338_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_11608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2338_base_resize_req_0); -- 
    base_resize_ack_11609_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_11613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2338_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2338_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_11621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2338_addr_0_req_0); -- 
    ra_11622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_11623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2338_addr_0_req_1); -- 
    ca_11624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_11628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2338_addr_1_req_0); -- 
    ra_11629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_11630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2338_addr_1_req_1); -- 
    ca_11631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2338_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_11643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2338_store_0_req_0); -- 
    ra_11644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_11648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2338_store_1_req_0); -- 
    ra_11649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_11659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2338_store_0_req_1); -- 
    ca_11660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_11664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2338_store_1_req_1); -- 
    ca_11665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2338_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2345_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_11675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2345_inst_ack_0, ack => cp_elements(55)); -- 
    cr_11676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2345_inst_req_1); -- 
    ca_11677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2345_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11686_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2349_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_11687_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2349_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2355_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_11697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2355_inst_ack_0, ack => cp_elements(63)); -- 
    cr_11698_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2355_inst_req_1); -- 
    ca_11699_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2355_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2359_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_11709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2366_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_11720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2366_base_resize_req_0); -- 
    base_resize_ack_11721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2366_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_11726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2366_root_address_inst_req_0); -- 
    plus_base_ra_11727_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2366_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_11728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2366_root_address_inst_req_1); -- 
    plus_base_ca_11729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2366_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2366_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_11747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2370_base_resize_req_0); -- 
    base_resize_ack_11748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_11752_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2370_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2370_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_11760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2370_addr_0_req_0); -- 
    ra_11761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_11762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2370_addr_0_req_1); -- 
    ca_11763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_11767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2370_addr_1_req_0); -- 
    ra_11768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_11769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2370_addr_1_req_1); -- 
    ca_11770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_11774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2370_addr_2_req_0); -- 
    ra_11775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_11776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2370_addr_2_req_1); -- 
    ca_11777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_11781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2370_addr_3_req_0); -- 
    ra_11782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_11783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2370_addr_3_req_1); -- 
    ca_11784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_11794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2370_load_0_req_0); -- 
    ra_11795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_11799_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2370_load_1_req_0); -- 
    ra_11800_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_11804_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2370_load_2_req_0); -- 
    ra_11805_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_11809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2370_load_3_req_0); -- 
    ra_11810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_11820_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2370_load_0_req_1); -- 
    ca_11821_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_11825_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2370_load_1_req_1); -- 
    ca_11826_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_11830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2370_load_2_req_1); -- 
    ca_11831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_11835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2370_load_3_req_1); -- 
    ca_11836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_11837_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2370_gather_scatter_req_0); -- 
    merge_ack_11838_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2370_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2374_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_11848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2374_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11872_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2381_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_11859_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2381_base_resize_req_0); -- 
    base_resize_ack_11860_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2381_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_11865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2381_root_address_inst_req_0); -- 
    plus_base_ra_11866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2381_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_11867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2381_root_address_inst_req_1); -- 
    plus_base_ca_11868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2381_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2381_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_11886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2385_base_resize_req_0); -- 
    base_resize_ack_11887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_11891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2385_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2385_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_11899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2385_addr_0_req_0); -- 
    ra_11900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_11901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2385_addr_0_req_1); -- 
    ca_11902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_11906_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2385_addr_1_req_0); -- 
    ra_11907_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_11908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2385_addr_1_req_1); -- 
    ca_11909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_11913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2385_addr_2_req_0); -- 
    ra_11914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_11915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2385_addr_2_req_1); -- 
    ca_11916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_11920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2385_addr_3_req_0); -- 
    ra_11921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_11922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2385_addr_3_req_1); -- 
    ca_11923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_11933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2385_load_0_req_0); -- 
    ra_11934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_11938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2385_load_1_req_0); -- 
    ra_11939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_11943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2385_load_2_req_0); -- 
    ra_11944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_11948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2385_load_3_req_0); -- 
    ra_11949_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_11959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2385_load_0_req_1); -- 
    ca_11960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_11964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2385_load_1_req_1); -- 
    ca_11965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_11969_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2385_load_2_req_1); -- 
    ca_11970_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_11974_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2385_load_3_req_1); -- 
    ca_11975_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_11976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2385_gather_scatter_req_0); -- 
    merge_ack_11977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2385_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2389_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_11987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11997_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_2394_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_11998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2394_inst_ack_0, ack => cp_elements(162)); -- 
    cr_11999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_2394_inst_req_1); -- 
    cp_elements(163) <= binary_2394_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_2398_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_12010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2398_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_2404_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_12020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2404_inst_ack_0, ack => cp_elements(171)); -- 
    cr_12021_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_2404_inst_req_1); -- 
    ca_12022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2404_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_2408_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_12032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2408_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12041_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2414_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_12042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2414_inst_ack_0, ack => cp_elements(178)); -- 
    cr_12043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_2414_inst_req_1); -- 
    ca_12044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2414_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_2420_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_12054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2420_inst_ack_0, ack => cp_elements(183)); -- 
    cr_12055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2420_inst_req_1); -- 
    ca_12056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2420_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_2428_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12067_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_2424_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_12068_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2424_inst_ack_0, ack => cp_elements(189)); -- 
    ra_12073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2428_inst_ack_0, ack => cp_elements(190)); -- 
    cr_12074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_2428_inst_req_1); -- 
    ca_12075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2428_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_2432_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_12085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_2437_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_12096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2437_inst_ack_0, ack => cp_elements(197)); -- 
    cr_12097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_2437_inst_req_1); -- 
    ca_12098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2437_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_12109_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2441_call_ack_0, ack => cp_elements(200)); -- 
    ccr_12113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_2441_call_req_1); -- 
    cca_12114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2441_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_12160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_2443_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_12133_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_2443_base_resize_req_0); -- 
    base_resize_ack_12134_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_12138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2443_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_2443_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_12146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2443_addr_0_req_0); -- 
    ra_12147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_12148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_2443_addr_0_req_1); -- 
    ca_12149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_12153_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_2443_addr_1_req_0); -- 
    ra_12154_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_12155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2443_addr_1_req_1); -- 
    ca_12156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_2443_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_12168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2443_store_0_req_0); -- 
    ra_12169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_12173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2443_store_1_req_0); -- 
    ra_12174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_12184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_2443_store_0_req_1); -- 
    ca_12185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_12189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_2443_store_1_req_1); -- 
    ca_12190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2443_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_12200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_2448_call_req_0); -- 
    cra_12201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2448_call_ack_0, ack => cp_elements(227)); -- 
    ccr_12205_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_2448_call_req_1); -- 
    cca_12206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2448_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_12252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_2450_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_12225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_2450_base_resize_req_0); -- 
    base_resize_ack_12226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_12230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_2450_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_2450_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_12238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_2450_addr_0_req_0); -- 
    ra_12239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_12240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_2450_addr_0_req_1); -- 
    ca_12241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_12245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_2450_addr_1_req_0); -- 
    ra_12246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_12247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_2450_addr_1_req_1); -- 
    ca_12248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_2450_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_12260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_2450_store_0_req_0); -- 
    ra_12261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_12265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2450_store_1_req_0); -- 
    ra_12266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_12276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_2450_store_0_req_1); -- 
    ca_12277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_12281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2450_store_1_req_1); -- 
    ca_12282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_12295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_2455_base_resize_req_0); -- 
    base_resize_ack_12296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_12300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_2455_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_2455_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_12308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_2455_addr_0_req_0); -- 
    ra_12309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_12310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2455_addr_0_req_1); -- 
    ca_12311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_12315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2455_addr_1_req_0); -- 
    ra_12316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_12317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_2455_addr_1_req_1); -- 
    ca_12318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_12322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_2455_addr_2_req_0); -- 
    ra_12323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_12324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_2455_addr_2_req_1); -- 
    ca_12325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_12329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_2455_addr_3_req_0); -- 
    ra_12330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_12331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2455_addr_3_req_1); -- 
    ca_12332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_12342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2455_load_0_req_0); -- 
    ra_12343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_12347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_2455_load_1_req_0); -- 
    ra_12348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_12352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2455_load_2_req_0); -- 
    ra_12353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_12357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2455_load_3_req_0); -- 
    ra_12358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_12368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2455_load_0_req_1); -- 
    ca_12369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_12373_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_2455_load_1_req_1); -- 
    ca_12374_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_12378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2455_load_2_req_1); -- 
    ca_12379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_12383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2455_load_3_req_1); -- 
    ca_12384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_2455_gather_scatter_req_0); -- 
    merge_ack_12386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_2459_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_12396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2459_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_12407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2461_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_2467_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_12420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2467_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_12425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_2465_inst_req_0); -- 
    pipe_wack_12426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2465_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2366_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2366_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2366_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2381_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2381_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2381_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_2429 : std_logic_vector(0 downto 0);
    signal ptr_deref_2338_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2338_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2338_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2338_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2338_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2338_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2338_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2338_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2338_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2370_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2370_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2370_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2370_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2370_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2385_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2385_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2385_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2385_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2385_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2443_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2443_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2443_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2450_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2450_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2455_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2455_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2455_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2455_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2316_wire : std_logic_vector(31 downto 0);
    signal tmp10_2371 : std_logic_vector(31 downto 0);
    signal tmp11_2375 : std_logic_vector(31 downto 0);
    signal tmp12_2382 : std_logic_vector(31 downto 0);
    signal tmp13_2386 : std_logic_vector(31 downto 0);
    signal tmp14_2390 : std_logic_vector(31 downto 0);
    signal tmp15_2395 : std_logic_vector(31 downto 0);
    signal tmp16_2399 : std_logic_vector(15 downto 0);
    signal tmp17_2405 : std_logic_vector(31 downto 0);
    signal tmp18_2415 : std_logic_vector(15 downto 0);
    signal tmp19_2421 : std_logic_vector(31 downto 0);
    signal tmp1_2322 : std_logic_vector(31 downto 0);
    signal tmp20_2433 : std_logic_vector(15 downto 0);
    signal tmp21_2438 : std_logic_vector(15 downto 0);
    signal tmp22_2441 : std_logic_vector(15 downto 0);
    signal tmp23_2448 : std_logic_vector(15 downto 0);
    signal tmp24_2456 : std_logic_vector(31 downto 0);
    signal tmp25_2460 : std_logic_vector(31 downto 0);
    signal tmp2_2328 : std_logic_vector(31 downto 0);
    signal tmp3_2332 : std_logic_vector(31 downto 0);
    signal tmp4_2336 : std_logic_vector(15 downto 0);
    signal tmp5_2346 : std_logic_vector(31 downto 0);
    signal tmp6_2350 : std_logic_vector(31 downto 0);
    signal tmp7_2356 : std_logic_vector(31 downto 0);
    signal tmp8_2360 : std_logic_vector(31 downto 0);
    signal tmp9_2367 : std_logic_vector(31 downto 0);
    signal tmp_2318 : std_logic_vector(31 downto 0);
    signal type_cast_2326_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2334_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2344_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2354_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2403_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2413_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2424_wire : std_logic_vector(31 downto 0);
    signal type_cast_2427_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2463_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2467_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_2409 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2366_final_offset <= "0000000000010000";
    array_obj_ref_2381_final_offset <= "0000000000001100";
    ptr_deref_2338_word_offset_0 <= "0000000000000000";
    ptr_deref_2338_word_offset_1 <= "0000000000000001";
    ptr_deref_2370_word_offset_0 <= "0000000000000000";
    ptr_deref_2370_word_offset_1 <= "0000000000000001";
    ptr_deref_2370_word_offset_2 <= "0000000000000010";
    ptr_deref_2370_word_offset_3 <= "0000000000000011";
    ptr_deref_2385_word_offset_0 <= "0000000000000000";
    ptr_deref_2385_word_offset_1 <= "0000000000000001";
    ptr_deref_2385_word_offset_2 <= "0000000000000010";
    ptr_deref_2385_word_offset_3 <= "0000000000000011";
    ptr_deref_2443_word_offset_0 <= "0000000000000000";
    ptr_deref_2443_word_offset_1 <= "0000000000000001";
    ptr_deref_2450_word_offset_0 <= "0000000000000000";
    ptr_deref_2450_word_offset_1 <= "0000000000000001";
    ptr_deref_2455_word_offset_0 <= "0000000000000000";
    ptr_deref_2455_word_offset_1 <= "0000000000000001";
    ptr_deref_2455_word_offset_2 <= "0000000000000010";
    ptr_deref_2455_word_offset_3 <= "0000000000000011";
    type_cast_2326_wire_constant <= "11111111111111111111100000000000";
    type_cast_2334_wire_constant <= "0000000000001000";
    type_cast_2344_wire_constant <= "00000000000000000000000000000110";
    type_cast_2354_wire_constant <= "00000000000000000000000000000010";
    type_cast_2403_wire_constant <= "00000000000000000000000000000011";
    type_cast_2413_wire_constant <= "0001111111111111";
    type_cast_2419_wire_constant <= "00000000000000000000000000000111";
    type_cast_2427_wire_constant <= "00000000000000000000000000000000";
    type_cast_2463_wire_constant <= "00000000000000000000000000000100";
    array_obj_ref_2366_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2322, dout => array_obj_ref_2366_resized_base_address, req => array_obj_ref_2366_base_resize_req_0, ack => array_obj_ref_2366_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2366_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2366_root_address, dout => tmp9_2367, req => array_obj_ref_2366_final_reg_req_0, ack => array_obj_ref_2366_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2381_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2322, dout => array_obj_ref_2381_resized_base_address, req => array_obj_ref_2381_base_resize_req_0, ack => array_obj_ref_2381_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2381_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2381_root_address, dout => tmp12_2382, req => array_obj_ref_2381_final_reg_req_0, ack => array_obj_ref_2381_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2338_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2332, dout => ptr_deref_2338_resized_base_address, req => ptr_deref_2338_base_resize_req_0, ack => ptr_deref_2338_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2370_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2367, dout => ptr_deref_2370_resized_base_address, req => ptr_deref_2370_base_resize_req_0, ack => ptr_deref_2370_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2385_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2382, dout => ptr_deref_2385_resized_base_address, req => ptr_deref_2385_base_resize_req_0, ack => ptr_deref_2385_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2443_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2350, dout => ptr_deref_2443_resized_base_address, req => ptr_deref_2443_base_resize_req_0, ack => ptr_deref_2443_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2450_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2360, dout => ptr_deref_2450_resized_base_address, req => ptr_deref_2450_base_resize_req_0, ack => ptr_deref_2450_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2455_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2382, dout => ptr_deref_2455_resized_base_address, req => ptr_deref_2455_base_resize_req_0, ack => ptr_deref_2455_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2317_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2316_wire, dout => tmp_2318, req => type_cast_2317_inst_req_0, ack => type_cast_2317_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2321_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_2318, dout => tmp1_2322, req => type_cast_2321_inst_req_0, ack => type_cast_2321_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2331_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2328, dout => tmp3_2332, req => type_cast_2331_inst_req_0, ack => type_cast_2331_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2349_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2346, dout => tmp6_2350, req => type_cast_2349_inst_req_0, ack => type_cast_2349_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2359_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2356, dout => tmp8_2360, req => type_cast_2359_inst_req_0, ack => type_cast_2359_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2374_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2371, dout => tmp11_2375, req => type_cast_2374_inst_req_0, ack => type_cast_2374_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2389_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2386, dout => tmp14_2390, req => type_cast_2389_inst_req_0, ack => type_cast_2389_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2398_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_2395, dout => tmp16_2399, req => type_cast_2398_inst_req_0, ack => type_cast_2398_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2408_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_2405, dout => xx_xtrx_xi_2409, req => type_cast_2408_inst_req_0, ack => type_cast_2408_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2424_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_2421, dout => type_cast_2424_wire, req => type_cast_2424_inst_req_0, ack => type_cast_2424_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2432_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_2429, dout => tmp20_2433, req => type_cast_2432_inst_req_0, ack => type_cast_2432_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2459_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_2456, dout => tmp25_2460, req => type_cast_2459_inst_req_0, ack => type_cast_2459_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2467_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_2460, dout => type_cast_2467_wire, req => type_cast_2467_inst_req_0, ack => type_cast_2467_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2338_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2338_gather_scatter_ack_0 <= ptr_deref_2338_gather_scatter_req_0;
      aggregated_sig <= tmp4_2336;
      ptr_deref_2338_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2338_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2338_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2338_root_address_inst_ack_0 <= ptr_deref_2338_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2338_resized_base_address;
      ptr_deref_2338_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2370_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2370_gather_scatter_ack_0 <= ptr_deref_2370_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2370_data_3 & ptr_deref_2370_data_2 & ptr_deref_2370_data_1 & ptr_deref_2370_data_0;
      tmp10_2371 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2370_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2370_root_address_inst_ack_0 <= ptr_deref_2370_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2370_resized_base_address;
      ptr_deref_2370_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2385_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2385_gather_scatter_ack_0 <= ptr_deref_2385_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2385_data_3 & ptr_deref_2385_data_2 & ptr_deref_2385_data_1 & ptr_deref_2385_data_0;
      tmp13_2386 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2385_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2385_root_address_inst_ack_0 <= ptr_deref_2385_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2385_resized_base_address;
      ptr_deref_2385_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2443_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2443_gather_scatter_ack_0 <= ptr_deref_2443_gather_scatter_req_0;
      aggregated_sig <= tmp22_2441;
      ptr_deref_2443_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2443_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2443_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2443_root_address_inst_ack_0 <= ptr_deref_2443_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2443_resized_base_address;
      ptr_deref_2443_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2450_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2450_gather_scatter_ack_0 <= ptr_deref_2450_gather_scatter_req_0;
      aggregated_sig <= tmp23_2448;
      ptr_deref_2450_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2450_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2450_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2450_root_address_inst_ack_0 <= ptr_deref_2450_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2450_resized_base_address;
      ptr_deref_2450_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2455_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2455_gather_scatter_ack_0 <= ptr_deref_2455_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2455_data_3 & ptr_deref_2455_data_2 & ptr_deref_2455_data_1 & ptr_deref_2455_data_0;
      tmp24_2456 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2455_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2455_root_address_inst_ack_0 <= ptr_deref_2455_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2455_resized_base_address;
      ptr_deref_2455_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2366_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2366_resized_base_address;
      array_obj_ref_2366_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2366_root_address_inst_req_0,
          ackL => array_obj_ref_2366_root_address_inst_ack_0,
          reqR => array_obj_ref_2366_root_address_inst_req_1,
          ackR => array_obj_ref_2366_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2381_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2381_resized_base_address;
      array_obj_ref_2381_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2381_root_address_inst_req_0,
          ackL => array_obj_ref_2381_root_address_inst_ack_0,
          reqR => array_obj_ref_2381_root_address_inst_req_1,
          ackR => array_obj_ref_2381_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2327_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2318;
      tmp2_2328 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2327_inst_req_0,
          ackL => binary_2327_inst_ack_0,
          reqR => binary_2327_inst_req_1,
          ackR => binary_2327_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2345_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2328;
      tmp5_2346 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2345_inst_req_0,
          ackL => binary_2345_inst_ack_0,
          reqR => binary_2345_inst_req_1,
          ackR => binary_2345_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2355_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2328;
      tmp7_2356 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2355_inst_req_0,
          ackL => binary_2355_inst_ack_0,
          reqR => binary_2355_inst_req_1,
          ackR => binary_2355_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2394_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2375 & tmp14_2390;
      tmp15_2395 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2394_inst_req_0,
          ackL => binary_2394_inst_ack_0,
          reqR => binary_2394_inst_req_1,
          ackR => binary_2394_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2404_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2395;
      tmp17_2405 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2404_inst_req_0,
          ackL => binary_2404_inst_ack_0,
          reqR => binary_2404_inst_req_1,
          ackR => binary_2404_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2414_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_2409;
      tmp18_2415 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2414_inst_req_0,
          ackL => binary_2414_inst_ack_0,
          reqR => binary_2414_inst_req_1,
          ackR => binary_2414_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2420_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2395;
      tmp19_2421 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2420_inst_req_0,
          ackL => binary_2420_inst_ack_0,
          reqR => binary_2420_inst_req_1,
          ackR => binary_2420_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2428_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2424_wire;
      notx_xx_xi_2429 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2428_inst_req_0,
          ackL => binary_2428_inst_ack_0,
          reqR => binary_2428_inst_req_1,
          ackR => binary_2428_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2437_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_2415 & tmp20_2433;
      tmp21_2438 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2437_inst_req_0,
          ackL => binary_2437_inst_ack_0,
          reqR => binary_2437_inst_req_1,
          ackR => binary_2437_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2338_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2338_root_address;
      ptr_deref_2338_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2338_addr_0_req_0,
          ackL => ptr_deref_2338_addr_0_ack_0,
          reqR => ptr_deref_2338_addr_0_req_1,
          ackR => ptr_deref_2338_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2338_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2338_root_address;
      ptr_deref_2338_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2338_addr_1_req_0,
          ackL => ptr_deref_2338_addr_1_ack_0,
          reqR => ptr_deref_2338_addr_1_req_1,
          ackR => ptr_deref_2338_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2370_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2370_root_address;
      ptr_deref_2370_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2370_addr_0_req_0,
          ackL => ptr_deref_2370_addr_0_ack_0,
          reqR => ptr_deref_2370_addr_0_req_1,
          ackR => ptr_deref_2370_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2370_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2370_root_address;
      ptr_deref_2370_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2370_addr_1_req_0,
          ackL => ptr_deref_2370_addr_1_ack_0,
          reqR => ptr_deref_2370_addr_1_req_1,
          ackR => ptr_deref_2370_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2370_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2370_root_address;
      ptr_deref_2370_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2370_addr_2_req_0,
          ackL => ptr_deref_2370_addr_2_ack_0,
          reqR => ptr_deref_2370_addr_2_req_1,
          ackR => ptr_deref_2370_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2370_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2370_root_address;
      ptr_deref_2370_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2370_addr_3_req_0,
          ackL => ptr_deref_2370_addr_3_ack_0,
          reqR => ptr_deref_2370_addr_3_req_1,
          ackR => ptr_deref_2370_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2385_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2385_root_address;
      ptr_deref_2385_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2385_addr_0_req_0,
          ackL => ptr_deref_2385_addr_0_ack_0,
          reqR => ptr_deref_2385_addr_0_req_1,
          ackR => ptr_deref_2385_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2385_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2385_root_address;
      ptr_deref_2385_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2385_addr_1_req_0,
          ackL => ptr_deref_2385_addr_1_ack_0,
          reqR => ptr_deref_2385_addr_1_req_1,
          ackR => ptr_deref_2385_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2385_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2385_root_address;
      ptr_deref_2385_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2385_addr_2_req_0,
          ackL => ptr_deref_2385_addr_2_ack_0,
          reqR => ptr_deref_2385_addr_2_req_1,
          ackR => ptr_deref_2385_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2385_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2385_root_address;
      ptr_deref_2385_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2385_addr_3_req_0,
          ackL => ptr_deref_2385_addr_3_ack_0,
          reqR => ptr_deref_2385_addr_3_req_1,
          ackR => ptr_deref_2385_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2443_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2443_root_address;
      ptr_deref_2443_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2443_addr_0_req_0,
          ackL => ptr_deref_2443_addr_0_ack_0,
          reqR => ptr_deref_2443_addr_0_req_1,
          ackR => ptr_deref_2443_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2443_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2443_root_address;
      ptr_deref_2443_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2443_addr_1_req_0,
          ackL => ptr_deref_2443_addr_1_ack_0,
          reqR => ptr_deref_2443_addr_1_req_1,
          ackR => ptr_deref_2443_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2450_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2450_root_address;
      ptr_deref_2450_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2450_addr_0_req_0,
          ackL => ptr_deref_2450_addr_0_ack_0,
          reqR => ptr_deref_2450_addr_0_req_1,
          ackR => ptr_deref_2450_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2450_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2450_root_address;
      ptr_deref_2450_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2450_addr_1_req_0,
          ackL => ptr_deref_2450_addr_1_ack_0,
          reqR => ptr_deref_2450_addr_1_req_1,
          ackR => ptr_deref_2450_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2455_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2455_root_address;
      ptr_deref_2455_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2455_addr_0_req_0,
          ackL => ptr_deref_2455_addr_0_ack_0,
          reqR => ptr_deref_2455_addr_0_req_1,
          ackR => ptr_deref_2455_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2455_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2455_root_address;
      ptr_deref_2455_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2455_addr_1_req_0,
          ackL => ptr_deref_2455_addr_1_ack_0,
          reqR => ptr_deref_2455_addr_1_req_1,
          ackR => ptr_deref_2455_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2455_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2455_root_address;
      ptr_deref_2455_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2455_addr_2_req_0,
          ackL => ptr_deref_2455_addr_2_ack_0,
          reqR => ptr_deref_2455_addr_2_req_1,
          ackR => ptr_deref_2455_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2455_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2455_root_address;
      ptr_deref_2455_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2455_addr_3_req_0,
          ackL => ptr_deref_2455_addr_3_ack_0,
          reqR => ptr_deref_2455_addr_3_req_1,
          ackR => ptr_deref_2455_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2370_load_0 ptr_deref_2370_load_1 ptr_deref_2370_load_2 ptr_deref_2370_load_3 ptr_deref_2385_load_0 ptr_deref_2385_load_1 ptr_deref_2385_load_2 ptr_deref_2385_load_3 ptr_deref_2455_load_0 ptr_deref_2455_load_1 ptr_deref_2455_load_2 ptr_deref_2455_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2370_load_0_req_0,
        ptr_deref_2370_load_0_ack_0,
        ptr_deref_2370_load_0_req_1,
        ptr_deref_2370_load_0_ack_1,
        "ptr_deref_2370_load_0",
        "memory_space_5" ,
        ptr_deref_2370_data_0,
        ptr_deref_2370_word_address_0,
        "ptr_deref_2370_data_0",
        "ptr_deref_2370_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2370_load_1_req_0,
        ptr_deref_2370_load_1_ack_0,
        ptr_deref_2370_load_1_req_1,
        ptr_deref_2370_load_1_ack_1,
        "ptr_deref_2370_load_1",
        "memory_space_5" ,
        ptr_deref_2370_data_1,
        ptr_deref_2370_word_address_1,
        "ptr_deref_2370_data_1",
        "ptr_deref_2370_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2370_load_2_req_0,
        ptr_deref_2370_load_2_ack_0,
        ptr_deref_2370_load_2_req_1,
        ptr_deref_2370_load_2_ack_1,
        "ptr_deref_2370_load_2",
        "memory_space_5" ,
        ptr_deref_2370_data_2,
        ptr_deref_2370_word_address_2,
        "ptr_deref_2370_data_2",
        "ptr_deref_2370_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2370_load_3_req_0,
        ptr_deref_2370_load_3_ack_0,
        ptr_deref_2370_load_3_req_1,
        ptr_deref_2370_load_3_ack_1,
        "ptr_deref_2370_load_3",
        "memory_space_5" ,
        ptr_deref_2370_data_3,
        ptr_deref_2370_word_address_3,
        "ptr_deref_2370_data_3",
        "ptr_deref_2370_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2385_load_0_req_0,
        ptr_deref_2385_load_0_ack_0,
        ptr_deref_2385_load_0_req_1,
        ptr_deref_2385_load_0_ack_1,
        "ptr_deref_2385_load_0",
        "memory_space_5" ,
        ptr_deref_2385_data_0,
        ptr_deref_2385_word_address_0,
        "ptr_deref_2385_data_0",
        "ptr_deref_2385_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2385_load_1_req_0,
        ptr_deref_2385_load_1_ack_0,
        ptr_deref_2385_load_1_req_1,
        ptr_deref_2385_load_1_ack_1,
        "ptr_deref_2385_load_1",
        "memory_space_5" ,
        ptr_deref_2385_data_1,
        ptr_deref_2385_word_address_1,
        "ptr_deref_2385_data_1",
        "ptr_deref_2385_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2385_load_2_req_0,
        ptr_deref_2385_load_2_ack_0,
        ptr_deref_2385_load_2_req_1,
        ptr_deref_2385_load_2_ack_1,
        "ptr_deref_2385_load_2",
        "memory_space_5" ,
        ptr_deref_2385_data_2,
        ptr_deref_2385_word_address_2,
        "ptr_deref_2385_data_2",
        "ptr_deref_2385_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2385_load_3_req_0,
        ptr_deref_2385_load_3_ack_0,
        ptr_deref_2385_load_3_req_1,
        ptr_deref_2385_load_3_ack_1,
        "ptr_deref_2385_load_3",
        "memory_space_5" ,
        ptr_deref_2385_data_3,
        ptr_deref_2385_word_address_3,
        "ptr_deref_2385_data_3",
        "ptr_deref_2385_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2455_load_0_req_0,
        ptr_deref_2455_load_0_ack_0,
        ptr_deref_2455_load_0_req_1,
        ptr_deref_2455_load_0_ack_1,
        "ptr_deref_2455_load_0",
        "memory_space_5" ,
        ptr_deref_2455_data_0,
        ptr_deref_2455_word_address_0,
        "ptr_deref_2455_data_0",
        "ptr_deref_2455_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2455_load_1_req_0,
        ptr_deref_2455_load_1_ack_0,
        ptr_deref_2455_load_1_req_1,
        ptr_deref_2455_load_1_ack_1,
        "ptr_deref_2455_load_1",
        "memory_space_5" ,
        ptr_deref_2455_data_1,
        ptr_deref_2455_word_address_1,
        "ptr_deref_2455_data_1",
        "ptr_deref_2455_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2455_load_2_req_0,
        ptr_deref_2455_load_2_ack_0,
        ptr_deref_2455_load_2_req_1,
        ptr_deref_2455_load_2_ack_1,
        "ptr_deref_2455_load_2",
        "memory_space_5" ,
        ptr_deref_2455_data_2,
        ptr_deref_2455_word_address_2,
        "ptr_deref_2455_data_2",
        "ptr_deref_2455_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2455_load_3_req_0,
        ptr_deref_2455_load_3_ack_0,
        ptr_deref_2455_load_3_req_1,
        ptr_deref_2455_load_3_ack_1,
        "ptr_deref_2455_load_3",
        "memory_space_5" ,
        ptr_deref_2455_data_3,
        ptr_deref_2455_word_address_3,
        "ptr_deref_2455_data_3",
        "ptr_deref_2455_word_address_3" -- 
      );
      reqL(11) <= ptr_deref_2370_load_0_req_0;
      reqL(10) <= ptr_deref_2370_load_1_req_0;
      reqL(9) <= ptr_deref_2370_load_2_req_0;
      reqL(8) <= ptr_deref_2370_load_3_req_0;
      reqL(7) <= ptr_deref_2385_load_0_req_0;
      reqL(6) <= ptr_deref_2385_load_1_req_0;
      reqL(5) <= ptr_deref_2385_load_2_req_0;
      reqL(4) <= ptr_deref_2385_load_3_req_0;
      reqL(3) <= ptr_deref_2455_load_0_req_0;
      reqL(2) <= ptr_deref_2455_load_1_req_0;
      reqL(1) <= ptr_deref_2455_load_2_req_0;
      reqL(0) <= ptr_deref_2455_load_3_req_0;
      ptr_deref_2370_load_0_ack_0 <= ackL(11);
      ptr_deref_2370_load_1_ack_0 <= ackL(10);
      ptr_deref_2370_load_2_ack_0 <= ackL(9);
      ptr_deref_2370_load_3_ack_0 <= ackL(8);
      ptr_deref_2385_load_0_ack_0 <= ackL(7);
      ptr_deref_2385_load_1_ack_0 <= ackL(6);
      ptr_deref_2385_load_2_ack_0 <= ackL(5);
      ptr_deref_2385_load_3_ack_0 <= ackL(4);
      ptr_deref_2455_load_0_ack_0 <= ackL(3);
      ptr_deref_2455_load_1_ack_0 <= ackL(2);
      ptr_deref_2455_load_2_ack_0 <= ackL(1);
      ptr_deref_2455_load_3_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2370_load_0_req_1;
      reqR(10) <= ptr_deref_2370_load_1_req_1;
      reqR(9) <= ptr_deref_2370_load_2_req_1;
      reqR(8) <= ptr_deref_2370_load_3_req_1;
      reqR(7) <= ptr_deref_2385_load_0_req_1;
      reqR(6) <= ptr_deref_2385_load_1_req_1;
      reqR(5) <= ptr_deref_2385_load_2_req_1;
      reqR(4) <= ptr_deref_2385_load_3_req_1;
      reqR(3) <= ptr_deref_2455_load_0_req_1;
      reqR(2) <= ptr_deref_2455_load_1_req_1;
      reqR(1) <= ptr_deref_2455_load_2_req_1;
      reqR(0) <= ptr_deref_2455_load_3_req_1;
      ptr_deref_2370_load_0_ack_1 <= ackR(11);
      ptr_deref_2370_load_1_ack_1 <= ackR(10);
      ptr_deref_2370_load_2_ack_1 <= ackR(9);
      ptr_deref_2370_load_3_ack_1 <= ackR(8);
      ptr_deref_2385_load_0_ack_1 <= ackR(7);
      ptr_deref_2385_load_1_ack_1 <= ackR(6);
      ptr_deref_2385_load_2_ack_1 <= ackR(5);
      ptr_deref_2385_load_3_ack_1 <= ackR(4);
      ptr_deref_2455_load_0_ack_1 <= ackR(3);
      ptr_deref_2455_load_1_ack_1 <= ackR(2);
      ptr_deref_2455_load_2_ack_1 <= ackR(1);
      ptr_deref_2455_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_2370_word_address_0 & ptr_deref_2370_word_address_1 & ptr_deref_2370_word_address_2 & ptr_deref_2370_word_address_3 & ptr_deref_2385_word_address_0 & ptr_deref_2385_word_address_1 & ptr_deref_2385_word_address_2 & ptr_deref_2385_word_address_3 & ptr_deref_2455_word_address_0 & ptr_deref_2455_word_address_1 & ptr_deref_2455_word_address_2 & ptr_deref_2455_word_address_3;
      ptr_deref_2370_data_0 <= data_out(95 downto 88);
      ptr_deref_2370_data_1 <= data_out(87 downto 80);
      ptr_deref_2370_data_2 <= data_out(79 downto 72);
      ptr_deref_2370_data_3 <= data_out(71 downto 64);
      ptr_deref_2385_data_0 <= data_out(63 downto 56);
      ptr_deref_2385_data_1 <= data_out(55 downto 48);
      ptr_deref_2385_data_2 <= data_out(47 downto 40);
      ptr_deref_2385_data_3 <= data_out(39 downto 32);
      ptr_deref_2455_data_0 <= data_out(31 downto 24);
      ptr_deref_2455_data_1 <= data_out(23 downto 16);
      ptr_deref_2455_data_2 <= data_out(15 downto 8);
      ptr_deref_2455_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2338_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2338_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2338_word_address_0) &  " data ptr_deref_2338_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2338_data_0) severity note; --
        end if;
        if ptr_deref_2338_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2338_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2338_word_address_1) &  " data ptr_deref_2338_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2338_data_1) severity note; --
        end if;
        if ptr_deref_2443_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2443_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2443_word_address_0) &  " data ptr_deref_2443_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2443_data_0) severity note; --
        end if;
        if ptr_deref_2443_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2443_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2443_word_address_1) &  " data ptr_deref_2443_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2443_data_1) severity note; --
        end if;
        if ptr_deref_2450_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2450_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2450_word_address_0) &  " data ptr_deref_2450_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2450_data_0) severity note; --
        end if;
        if ptr_deref_2450_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2450_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2450_word_address_1) &  " data ptr_deref_2450_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2450_data_1) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2338_store_0 ptr_deref_2338_store_1 ptr_deref_2443_store_0 ptr_deref_2443_store_1 ptr_deref_2450_store_0 ptr_deref_2450_store_1 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2338_store_0_req_0;
      reqL(4) <= ptr_deref_2338_store_1_req_0;
      reqL(3) <= ptr_deref_2443_store_0_req_0;
      reqL(2) <= ptr_deref_2443_store_1_req_0;
      reqL(1) <= ptr_deref_2450_store_0_req_0;
      reqL(0) <= ptr_deref_2450_store_1_req_0;
      ptr_deref_2338_store_0_ack_0 <= ackL(5);
      ptr_deref_2338_store_1_ack_0 <= ackL(4);
      ptr_deref_2443_store_0_ack_0 <= ackL(3);
      ptr_deref_2443_store_1_ack_0 <= ackL(2);
      ptr_deref_2450_store_0_ack_0 <= ackL(1);
      ptr_deref_2450_store_1_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2338_store_0_req_1;
      reqR(4) <= ptr_deref_2338_store_1_req_1;
      reqR(3) <= ptr_deref_2443_store_0_req_1;
      reqR(2) <= ptr_deref_2443_store_1_req_1;
      reqR(1) <= ptr_deref_2450_store_0_req_1;
      reqR(0) <= ptr_deref_2450_store_1_req_1;
      ptr_deref_2338_store_0_ack_1 <= ackR(5);
      ptr_deref_2338_store_1_ack_1 <= ackR(4);
      ptr_deref_2443_store_0_ack_1 <= ackR(3);
      ptr_deref_2443_store_1_ack_1 <= ackR(2);
      ptr_deref_2450_store_0_ack_1 <= ackR(1);
      ptr_deref_2450_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2338_word_address_0 & ptr_deref_2338_word_address_1 & ptr_deref_2443_word_address_0 & ptr_deref_2443_word_address_1 & ptr_deref_2450_word_address_0 & ptr_deref_2450_word_address_1;
      data_in <= ptr_deref_2338_data_0 & ptr_deref_2338_data_1 & ptr_deref_2443_data_0 & ptr_deref_2443_data_1 & ptr_deref_2450_data_0 & ptr_deref_2450_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2316_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2316_inst_ack_0 then -- 
            assert false report " ReadPipe to3_in0 to wire simple_obj_ref_2316_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2316_inst_req_0;
      simple_obj_ref_2316_inst_ack_0 <= ack(0);
      simple_obj_ref_2316_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to3_in0_pipe_read_req(0),
          oack => to3_in0_pipe_read_ack(0),
          odata => to3_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2461_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_2463_wire_constant value="  &  convert_slv_to_hex_string(type_cast_2463_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2461_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2461_inst_req_0;
      simple_obj_ref_2461_inst_ack_0 <= ack(0);
      data_in <= type_cast_2463_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2465_inst_ack_0 then -- 
          assert false report " WritePipe tofpga3_out0 from wire type_cast_2467_wire value="  &  convert_slv_to_hex_string(type_cast_2467_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2465_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2465_inst_req_0;
      simple_obj_ref_2465_inst_ack_0 <= ack(0);
      data_in <= type_cast_2467_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga3_out0_pipe_write_req(0),
          oack => tofpga3_out0_pipe_write_ack(0),
          odata => tofpga3_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2336_call call_stmt_2441_call call_stmt_2448_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2336_call_req_0;
      reqL(1) <= call_stmt_2441_call_req_0;
      reqL(0) <= call_stmt_2448_call_req_0;
      call_stmt_2336_call_ack_0 <= ackL(2);
      call_stmt_2441_call_ack_0 <= ackL(1);
      call_stmt_2448_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2336_call_req_1;
      reqR(1) <= call_stmt_2441_call_req_1;
      reqR(0) <= call_stmt_2448_call_req_1;
      call_stmt_2336_call_ack_1 <= ackR(2);
      call_stmt_2441_call_ack_1 <= ackR(1);
      call_stmt_2448_call_ack_1 <= ackR(0);
      data_in <= type_cast_2334_wire_constant & tmp16_2399 & tmp21_2438;
      tmp4_2336 <= data_out(47 downto 32);
      tmp22_2441 <= data_out(31 downto 16);
      tmp23_2448 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_packet_free is -- 
  generic (tag_length : integer); 
  port ( -- 
    pkt : in  std_logic_vector(31 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_packet_free;
architecture Default of ahir_packet_free is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_packet_free_CP_1029_start: Boolean;
  -- links between control-path and data-path
  signal binary_2478_inst_req_0 : boolean;
  signal binary_2478_inst_ack_0 : boolean;
  signal binary_2478_inst_req_1 : boolean;
  signal binary_2478_inst_ack_1 : boolean;
  signal simple_obj_ref_2475_inst_req_0 : boolean;
  signal simple_obj_ref_2475_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_packet_free_CP_1029: Block -- control-path 
    signal cp_elements: BooleanArray(6 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(6);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(6), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cpelement_group_1 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(3));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => binary_2478_inst_req_0); -- 
    cp_elements(2) <= cp_elements(0);
    cp_elements(3) <= cp_elements(0);
    ra_1044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2478_inst_ack_0, ack => cp_elements(4)); -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => binary_2478_inst_req_1); -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2478_inst_ack_1, ack => cp_elements(5)); -- 
    pipe_wreq_1051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => simple_obj_ref_2475_inst_req_0); -- 
    pipe_wack_1052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2475_inst_ack_0, ack => cp_elements(6)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal binary_2478_wire : std_logic_vector(31 downto 0);
    signal expr_2477_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    expr_2477_wire_constant <= "11111111111111111111100000000000";
    -- shared split operator group (0) : binary_2478_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= pkt;
      binary_2478_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2478_inst_req_0,
          ackL => binary_2478_inst_ack_0,
          reqR => binary_2478_inst_req_1,
          ackR => binary_2478_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2475_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_2478_wire value="  &  convert_slv_to_hex_string(binary_2478_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2475_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2475_inst_req_0;
      simple_obj_ref_2475_inst_ack_0 <= ack(0);
      data_in <= binary_2478_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_packet_get is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf : out  std_logic_vector(31 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    free_queue_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_packet_get;
architecture Default of ahir_packet_get is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal buf_buffer :  std_logic_vector(31 downto 0);
  signal ahir_packet_get_CP_12435_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_2484_inst_req_0 : boolean;
  signal simple_obj_ref_2484_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  buf <= buf_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_packet_get_CP_12435: Block -- control-path 
    signal cp_elements: BooleanArray(1 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    req_12447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => simple_obj_ref_2484_inst_req_0); -- 
    ack_12448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2484_inst_ack_0, ack => cp_elements(1)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared inport operator group (0) : simple_obj_ref_2484_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2484_inst_ack_0 then -- 
            assert false report " ReadPipe free_queue_pipe to wire buf value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2484_inst_req_0;
      simple_obj_ref_2484_inst_ack_0 <= ack(0);
      buf_buffer <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_pipe_pipe_read_req(0),
          oack => free_queue_pipe_pipe_read_ack(0),
          odata => free_queue_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity analyze_packet is -- 
  generic (tag_length : integer); 
  port ( -- 
    pkt : in  std_logic_vector(31 downto 0);
    buf : out  std_logic_vector(31 downto 0);
    wlen : out  std_logic_vector(15 downto 0);
    blen : out  std_logic_vector(15 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity analyze_packet;
architecture Default of analyze_packet is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal buf_buffer :  std_logic_vector(31 downto 0);
  signal wlen_buffer :  std_logic_vector(15 downto 0);
  signal blen_buffer :  std_logic_vector(15 downto 0);
  signal analyze_packet_CP_12449_start: Boolean;
  -- links between control-path and data-path
  signal binary_2500_inst_ack_0 : boolean;
  signal binary_2500_inst_req_1 : boolean;
  signal binary_2500_inst_ack_1 : boolean;
  signal array_obj_ref_2516_base_resize_req_0 : boolean;
  signal simple_obj_ref_2510_inst_req_0 : boolean;
  signal type_cast_2494_inst_req_0 : boolean;
  signal type_cast_2494_inst_ack_0 : boolean;
  signal simple_obj_ref_2510_inst_ack_0 : boolean;
  signal type_cast_2504_inst_req_0 : boolean;
  signal binary_2500_inst_req_0 : boolean;
  signal type_cast_2504_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal array_obj_ref_2516_base_resize_ack_0 : boolean;
  signal array_obj_ref_2516_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2516_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2516_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2516_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2516_final_reg_req_0 : boolean;
  signal array_obj_ref_2516_final_reg_ack_0 : boolean;
  signal ptr_deref_2520_base_resize_req_0 : boolean;
  signal ptr_deref_2520_base_resize_ack_0 : boolean;
  signal ptr_deref_2520_root_address_inst_req_0 : boolean;
  signal ptr_deref_2520_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2520_addr_0_req_0 : boolean;
  signal ptr_deref_2520_addr_0_ack_0 : boolean;
  signal ptr_deref_2520_addr_0_req_1 : boolean;
  signal ptr_deref_2520_addr_0_ack_1 : boolean;
  signal ptr_deref_2520_addr_1_req_0 : boolean;
  signal ptr_deref_2520_addr_1_ack_0 : boolean;
  signal ptr_deref_2520_addr_1_req_1 : boolean;
  signal ptr_deref_2520_addr_1_ack_1 : boolean;
  signal ptr_deref_2520_load_0_req_0 : boolean;
  signal ptr_deref_2520_load_0_ack_0 : boolean;
  signal ptr_deref_2520_load_1_req_0 : boolean;
  signal ptr_deref_2520_load_1_ack_0 : boolean;
  signal ptr_deref_2520_load_0_req_1 : boolean;
  signal ptr_deref_2520_load_0_ack_1 : boolean;
  signal ptr_deref_2520_load_1_req_1 : boolean;
  signal ptr_deref_2520_load_1_ack_1 : boolean;
  signal ptr_deref_2520_gather_scatter_req_0 : boolean;
  signal ptr_deref_2520_gather_scatter_ack_0 : boolean;
  signal type_cast_2524_inst_req_0 : boolean;
  signal type_cast_2524_inst_ack_0 : boolean;
  signal array_obj_ref_2529_base_resize_req_0 : boolean;
  signal array_obj_ref_2529_base_resize_ack_0 : boolean;
  signal array_obj_ref_2529_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2529_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2529_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2529_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2529_final_reg_req_0 : boolean;
  signal array_obj_ref_2529_final_reg_ack_0 : boolean;
  signal ptr_deref_2533_base_resize_req_0 : boolean;
  signal ptr_deref_2533_base_resize_ack_0 : boolean;
  signal ptr_deref_2533_root_address_inst_req_0 : boolean;
  signal ptr_deref_2533_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2533_addr_0_req_0 : boolean;
  signal ptr_deref_2533_addr_0_ack_0 : boolean;
  signal ptr_deref_2533_addr_0_req_1 : boolean;
  signal ptr_deref_2533_addr_0_ack_1 : boolean;
  signal ptr_deref_2533_addr_1_req_0 : boolean;
  signal ptr_deref_2533_addr_1_ack_0 : boolean;
  signal ptr_deref_2533_addr_1_req_1 : boolean;
  signal ptr_deref_2533_addr_1_ack_1 : boolean;
  signal ptr_deref_2533_load_0_req_0 : boolean;
  signal ptr_deref_2533_load_0_ack_0 : boolean;
  signal ptr_deref_2533_load_1_req_0 : boolean;
  signal ptr_deref_2533_load_1_ack_0 : boolean;
  signal ptr_deref_2533_load_0_req_1 : boolean;
  signal ptr_deref_2533_load_0_ack_1 : boolean;
  signal ptr_deref_2533_load_1_req_1 : boolean;
  signal ptr_deref_2533_load_1_ack_1 : boolean;
  signal ptr_deref_2533_gather_scatter_req_0 : boolean;
  signal ptr_deref_2533_gather_scatter_ack_0 : boolean;
  signal type_cast_2537_inst_req_0 : boolean;
  signal type_cast_2537_inst_ack_0 : boolean;
  signal binary_2543_inst_req_0 : boolean;
  signal binary_2543_inst_ack_0 : boolean;
  signal binary_2543_inst_req_1 : boolean;
  signal binary_2543_inst_ack_1 : boolean;
  signal type_cast_2547_inst_req_0 : boolean;
  signal type_cast_2547_inst_ack_0 : boolean;
  signal type_cast_2551_inst_req_0 : boolean;
  signal type_cast_2551_inst_ack_0 : boolean;
  signal binary_2555_inst_req_0 : boolean;
  signal binary_2555_inst_ack_0 : boolean;
  signal binary_2555_inst_req_1 : boolean;
  signal binary_2555_inst_ack_1 : boolean;
  signal type_cast_2556_inst_req_0 : boolean;
  signal type_cast_2556_inst_ack_0 : boolean;
  signal binary_2561_inst_req_0 : boolean;
  signal binary_2561_inst_ack_0 : boolean;
  signal binary_2561_inst_req_1 : boolean;
  signal binary_2561_inst_ack_1 : boolean;
  signal type_cast_2565_inst_req_0 : boolean;
  signal type_cast_2565_inst_ack_0 : boolean;
  signal type_cast_2569_inst_req_0 : boolean;
  signal type_cast_2569_inst_ack_0 : boolean;
  signal array_obj_ref_2574_base_resize_req_0 : boolean;
  signal array_obj_ref_2574_base_resize_ack_0 : boolean;
  signal array_obj_ref_2574_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2574_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2574_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2574_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2574_final_reg_req_0 : boolean;
  signal array_obj_ref_2574_final_reg_ack_0 : boolean;
  signal ptr_deref_2578_base_resize_req_0 : boolean;
  signal ptr_deref_2578_base_resize_ack_0 : boolean;
  signal ptr_deref_2578_root_address_inst_req_0 : boolean;
  signal ptr_deref_2578_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2578_addr_0_req_0 : boolean;
  signal ptr_deref_2578_addr_0_ack_0 : boolean;
  signal ptr_deref_2578_addr_0_req_1 : boolean;
  signal ptr_deref_2578_addr_0_ack_1 : boolean;
  signal ptr_deref_2578_addr_1_req_0 : boolean;
  signal ptr_deref_2578_addr_1_ack_0 : boolean;
  signal ptr_deref_2578_addr_1_req_1 : boolean;
  signal ptr_deref_2578_addr_1_ack_1 : boolean;
  signal ptr_deref_2578_load_0_req_0 : boolean;
  signal ptr_deref_2578_load_0_ack_0 : boolean;
  signal ptr_deref_2578_load_1_req_0 : boolean;
  signal ptr_deref_2578_load_1_ack_0 : boolean;
  signal ptr_deref_2578_load_0_req_1 : boolean;
  signal ptr_deref_2578_load_0_ack_1 : boolean;
  signal ptr_deref_2578_load_1_req_1 : boolean;
  signal ptr_deref_2578_load_1_ack_1 : boolean;
  signal ptr_deref_2578_gather_scatter_req_0 : boolean;
  signal ptr_deref_2578_gather_scatter_ack_0 : boolean;
  signal type_cast_2582_inst_req_0 : boolean;
  signal type_cast_2582_inst_ack_0 : boolean;
  signal array_obj_ref_2587_base_resize_req_0 : boolean;
  signal array_obj_ref_2587_base_resize_ack_0 : boolean;
  signal array_obj_ref_2587_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2587_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2587_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2587_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2587_final_reg_req_0 : boolean;
  signal array_obj_ref_2587_final_reg_ack_0 : boolean;
  signal ptr_deref_2591_base_resize_req_0 : boolean;
  signal ptr_deref_2591_base_resize_ack_0 : boolean;
  signal ptr_deref_2591_root_address_inst_req_0 : boolean;
  signal ptr_deref_2591_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2591_addr_0_req_0 : boolean;
  signal ptr_deref_2591_addr_0_ack_0 : boolean;
  signal ptr_deref_2591_addr_0_req_1 : boolean;
  signal ptr_deref_2591_addr_0_ack_1 : boolean;
  signal ptr_deref_2591_addr_1_req_0 : boolean;
  signal ptr_deref_2591_addr_1_ack_0 : boolean;
  signal ptr_deref_2591_addr_1_req_1 : boolean;
  signal ptr_deref_2591_addr_1_ack_1 : boolean;
  signal ptr_deref_2591_load_0_req_0 : boolean;
  signal ptr_deref_2591_load_0_ack_0 : boolean;
  signal ptr_deref_2591_load_1_req_0 : boolean;
  signal ptr_deref_2591_load_1_ack_0 : boolean;
  signal ptr_deref_2591_load_0_req_1 : boolean;
  signal ptr_deref_2591_load_0_ack_1 : boolean;
  signal ptr_deref_2591_load_1_req_1 : boolean;
  signal ptr_deref_2591_load_1_ack_1 : boolean;
  signal ptr_deref_2591_gather_scatter_req_0 : boolean;
  signal ptr_deref_2591_gather_scatter_ack_0 : boolean;
  signal type_cast_2595_inst_req_0 : boolean;
  signal type_cast_2595_inst_ack_0 : boolean;
  signal binary_2601_inst_req_0 : boolean;
  signal binary_2601_inst_ack_0 : boolean;
  signal binary_2601_inst_req_1 : boolean;
  signal binary_2601_inst_ack_1 : boolean;
  signal type_cast_2605_inst_req_0 : boolean;
  signal type_cast_2605_inst_ack_0 : boolean;
  signal type_cast_2609_inst_req_0 : boolean;
  signal type_cast_2609_inst_ack_0 : boolean;
  signal binary_2613_inst_req_0 : boolean;
  signal binary_2613_inst_ack_0 : boolean;
  signal binary_2613_inst_req_1 : boolean;
  signal binary_2613_inst_ack_1 : boolean;
  signal type_cast_2614_inst_req_0 : boolean;
  signal type_cast_2614_inst_ack_0 : boolean;
  signal binary_2619_inst_req_0 : boolean;
  signal binary_2619_inst_ack_0 : boolean;
  signal binary_2619_inst_req_1 : boolean;
  signal binary_2619_inst_ack_1 : boolean;
  signal type_cast_2623_inst_req_0 : boolean;
  signal type_cast_2623_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  buf <= buf_buffer; 
  wlen <= wlen_buffer; 
  blen <= blen_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  analyze_packet_CP_12449: Block -- control-path 
    signal cp_elements: BooleanArray(198 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(198);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(198), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cpelement_group_1 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(3));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => type_cast_2494_inst_req_0); -- 
    cp_elements(2) <= cp_elements(0);
    cp_elements(3) <= cp_elements(0);
    ack_12464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2494_inst_ack_0, ack => cp_elements(4)); -- 
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(4) & cp_elements(6));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12473_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => binary_2500_inst_req_0); -- 
    cp_elements(6) <= cp_elements(0);
    ra_12474_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2500_inst_ack_0, ack => cp_elements(7)); -- 
    cr_12475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => binary_2500_inst_req_1); -- 
    cp_elements(8) <= binary_2500_inst_ack_1;
    cpelement_group_9 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(10) & cp_elements(11));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(9),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => type_cast_2504_inst_req_0); -- 
    cp_elements(10) <= cp_elements(0);
    cp_elements(11) <= cp_elements(8);
    cp_elements(12) <= type_cast_2504_inst_ack_0;
    cpelement_group_13 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(15));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(13),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => type_cast_2508_inst_req_0); -- 
    cp_elements(14) <= cp_elements(0);
    cp_elements(15) <= cp_elements(8);
    ack_12496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => cp_elements(16)); -- 
    base_resize_req_12515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_2516_base_resize_req_0); -- 
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(19));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(18) <= cp_elements(12);
    req_12503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => simple_obj_ref_2510_inst_req_0); -- 
    ack_12504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2510_inst_ack_0, ack => cp_elements(19)); -- 
    cp_elements(20) <= cp_elements(0);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(20) & cp_elements(24));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_2516_final_reg_req_0); -- 
    base_resize_ack_12516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2516_base_resize_ack_0, ack => cp_elements(22)); -- 
    plus_base_rr_12521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_2516_root_address_inst_req_0); -- 
    plus_base_ra_12522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2516_root_address_inst_ack_0, ack => cp_elements(23)); -- 
    plus_base_cr_12523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => array_obj_ref_2516_root_address_inst_req_1); -- 
    plus_base_ca_12524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2516_root_address_inst_ack_1, ack => cp_elements(24)); -- 
    cp_elements(25) <= array_obj_ref_2516_final_reg_ack_0;
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(25) & cp_elements(36));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(27) <= cp_elements(25);
    base_resize_req_12542_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => ptr_deref_2520_base_resize_req_0); -- 
    base_resize_ack_12543_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_base_resize_ack_0, ack => cp_elements(28)); -- 
    sum_rename_req_12547_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2520_root_address_inst_req_0); -- 
    cp_elements(29) <= ptr_deref_2520_root_address_inst_ack_0;
    cp_elements(30) <= cp_elements(29);
    rr_12555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2520_addr_0_req_0); -- 
    ra_12556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_addr_0_ack_0, ack => cp_elements(31)); -- 
    cr_12557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2520_addr_0_req_1); -- 
    ca_12558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_addr_0_ack_1, ack => cp_elements(32)); -- 
    cp_elements(33) <= cp_elements(29);
    rr_12562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2520_addr_1_req_0); -- 
    ra_12563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_addr_1_ack_0, ack => cp_elements(34)); -- 
    cr_12564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2520_addr_1_req_1); -- 
    ca_12565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_addr_1_ack_1, ack => cp_elements(35)); -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(35));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(37) <= cp_elements(26);
    rr_12575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2520_load_0_req_0); -- 
    ra_12576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_load_0_ack_0, ack => cp_elements(38)); -- 
    cp_elements(39) <= cp_elements(26);
    rr_12580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => ptr_deref_2520_load_1_req_0); -- 
    ra_12581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_load_1_ack_0, ack => cp_elements(40)); -- 
    cpelement_group_41 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(38) & cp_elements(40));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(41),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(42) <= cp_elements(41);
    cr_12591_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_2520_load_0_req_1); -- 
    ca_12592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_load_0_ack_1, ack => cp_elements(43)); -- 
    cp_elements(44) <= cp_elements(41);
    cr_12596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_2520_load_1_req_1); -- 
    ca_12597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_load_1_ack_1, ack => cp_elements(45)); -- 
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(43) & cp_elements(45));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12598_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_2520_gather_scatter_req_0); -- 
    merge_ack_12599_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2520_gather_scatter_ack_0, ack => cp_elements(47)); -- 
    cpelement_group_48 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(49) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(48),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => type_cast_2524_inst_req_0); -- 
    cp_elements(49) <= cp_elements(0);
    cp_elements(50) <= cp_elements(17);
    ack_12609_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2524_inst_ack_0, ack => cp_elements(51)); -- 
    base_resize_req_12620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_2529_base_resize_req_0); -- 
    cp_elements(52) <= cp_elements(0);
    cpelement_group_53 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(52) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(53),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_2529_final_reg_req_0); -- 
    base_resize_ack_12621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2529_base_resize_ack_0, ack => cp_elements(54)); -- 
    plus_base_rr_12626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => array_obj_ref_2529_root_address_inst_req_0); -- 
    plus_base_ra_12627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2529_root_address_inst_ack_0, ack => cp_elements(55)); -- 
    plus_base_cr_12628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => array_obj_ref_2529_root_address_inst_req_1); -- 
    plus_base_ca_12629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2529_root_address_inst_ack_1, ack => cp_elements(56)); -- 
    cp_elements(57) <= array_obj_ref_2529_final_reg_ack_0;
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(57) & cp_elements(68));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(59) <= cp_elements(57);
    base_resize_req_12647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => ptr_deref_2533_base_resize_req_0); -- 
    base_resize_ack_12648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_base_resize_ack_0, ack => cp_elements(60)); -- 
    sum_rename_req_12652_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => ptr_deref_2533_root_address_inst_req_0); -- 
    cp_elements(61) <= ptr_deref_2533_root_address_inst_ack_0;
    cp_elements(62) <= cp_elements(61);
    rr_12660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_2533_addr_0_req_0); -- 
    ra_12661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_addr_0_ack_0, ack => cp_elements(63)); -- 
    cr_12662_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_2533_addr_0_req_1); -- 
    ca_12663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_addr_0_ack_1, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(61);
    rr_12667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_2533_addr_1_req_0); -- 
    ra_12668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_addr_1_ack_0, ack => cp_elements(66)); -- 
    cr_12669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => ptr_deref_2533_addr_1_req_1); -- 
    ca_12670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_addr_1_ack_1, ack => cp_elements(67)); -- 
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(67));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(69) <= cp_elements(58);
    rr_12680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_2533_load_0_req_0); -- 
    ra_12681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_load_0_ack_0, ack => cp_elements(70)); -- 
    cp_elements(71) <= cp_elements(58);
    rr_12685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => ptr_deref_2533_load_1_req_0); -- 
    ra_12686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_load_1_ack_0, ack => cp_elements(72)); -- 
    cpelement_group_73 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(72));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(73),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(74) <= cp_elements(73);
    cr_12696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_2533_load_0_req_1); -- 
    ca_12697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_load_0_ack_1, ack => cp_elements(75)); -- 
    cp_elements(76) <= cp_elements(73);
    cr_12701_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2533_load_1_req_1); -- 
    ca_12702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_load_1_ack_1, ack => cp_elements(77)); -- 
    cpelement_group_78 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(77));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(78),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => ptr_deref_2533_gather_scatter_req_0); -- 
    merge_ack_12704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2533_gather_scatter_ack_0, ack => cp_elements(79)); -- 
    cpelement_group_80 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(79) & cp_elements(81));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(80),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => type_cast_2537_inst_req_0); -- 
    cp_elements(81) <= cp_elements(0);
    ack_12714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2537_inst_ack_0, ack => cp_elements(82)); -- 
    cpelement_group_83 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(83),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => binary_2543_inst_req_0); -- 
    cp_elements(84) <= cp_elements(0);
    ra_12724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2543_inst_ack_0, ack => cp_elements(85)); -- 
    cr_12725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => binary_2543_inst_req_1); -- 
    ca_12726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2543_inst_ack_1, ack => cp_elements(86)); -- 
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(47) & cp_elements(88));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => type_cast_2547_inst_req_0); -- 
    cp_elements(88) <= cp_elements(0);
    ack_12736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2547_inst_ack_0, ack => cp_elements(89)); -- 
    cpelement_group_90 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(98));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(90),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => type_cast_2556_inst_req_0); -- 
    cp_elements(91) <= cp_elements(0);
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(96));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => binary_2555_inst_req_0); -- 
    cp_elements(93) <= cp_elements(0);
    cpelement_group_94 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(95));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(94),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => type_cast_2551_inst_req_0); -- 
    cp_elements(95) <= cp_elements(0);
    ack_12750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2551_inst_ack_0, ack => cp_elements(96)); -- 
    ra_12755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2555_inst_ack_0, ack => cp_elements(97)); -- 
    cr_12756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => binary_2555_inst_req_1); -- 
    ca_12757_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2555_inst_ack_1, ack => cp_elements(98)); -- 
    ack_12762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2556_inst_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(86) & cp_elements(99) & cp_elements(101));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => binary_2561_inst_req_0); -- 
    cp_elements(101) <= cp_elements(0);
    ra_12773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2561_inst_ack_0, ack => cp_elements(102)); -- 
    cr_12774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => binary_2561_inst_req_1); -- 
    ca_12775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2561_inst_ack_1, ack => cp_elements(103)); -- 
    cpelement_group_104 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(103) & cp_elements(105));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(104),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => type_cast_2565_inst_req_0); -- 
    cp_elements(105) <= cp_elements(0);
    ack_12785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_0, ack => cp_elements(106)); -- 
    cpelement_group_107 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(108) & cp_elements(109));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => type_cast_2569_inst_req_0); -- 
    cp_elements(108) <= cp_elements(0);
    cp_elements(109) <= cp_elements(17);
    ack_12795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2569_inst_ack_0, ack => cp_elements(110)); -- 
    base_resize_req_12806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => array_obj_ref_2574_base_resize_req_0); -- 
    cp_elements(111) <= cp_elements(0);
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(111) & cp_elements(115));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => array_obj_ref_2574_final_reg_req_0); -- 
    base_resize_ack_12807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2574_base_resize_ack_0, ack => cp_elements(113)); -- 
    plus_base_rr_12812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => array_obj_ref_2574_root_address_inst_req_0); -- 
    plus_base_ra_12813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2574_root_address_inst_ack_0, ack => cp_elements(114)); -- 
    plus_base_cr_12814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => array_obj_ref_2574_root_address_inst_req_1); -- 
    plus_base_ca_12815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2574_root_address_inst_ack_1, ack => cp_elements(115)); -- 
    cp_elements(116) <= array_obj_ref_2574_final_reg_ack_0;
    cpelement_group_117 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(116) & cp_elements(127));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(118) <= cp_elements(116);
    base_resize_req_12833_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => ptr_deref_2578_base_resize_req_0); -- 
    base_resize_ack_12834_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_base_resize_ack_0, ack => cp_elements(119)); -- 
    sum_rename_req_12838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_2578_root_address_inst_req_0); -- 
    cp_elements(120) <= ptr_deref_2578_root_address_inst_ack_0;
    cp_elements(121) <= cp_elements(120);
    rr_12846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => ptr_deref_2578_addr_0_req_0); -- 
    ra_12847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_addr_0_ack_0, ack => cp_elements(122)); -- 
    cr_12848_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2578_addr_0_req_1); -- 
    ca_12849_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_addr_0_ack_1, ack => cp_elements(123)); -- 
    cp_elements(124) <= cp_elements(120);
    rr_12853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => ptr_deref_2578_addr_1_req_0); -- 
    ra_12854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_addr_1_ack_0, ack => cp_elements(125)); -- 
    cr_12855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2578_addr_1_req_1); -- 
    ca_12856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_addr_1_ack_1, ack => cp_elements(126)); -- 
    cpelement_group_127 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(123) & cp_elements(126));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(127),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(128) <= cp_elements(117);
    rr_12866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2578_load_0_req_0); -- 
    ra_12867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_load_0_ack_0, ack => cp_elements(129)); -- 
    cp_elements(130) <= cp_elements(117);
    rr_12871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => ptr_deref_2578_load_1_req_0); -- 
    ra_12872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_load_1_ack_0, ack => cp_elements(131)); -- 
    cpelement_group_132 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(129) & cp_elements(131));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(132),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(133) <= cp_elements(132);
    cr_12882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => ptr_deref_2578_load_0_req_1); -- 
    ca_12883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_load_0_ack_1, ack => cp_elements(134)); -- 
    cp_elements(135) <= cp_elements(132);
    cr_12887_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2578_load_1_req_1); -- 
    ca_12888_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_load_1_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(137), ack => ptr_deref_2578_gather_scatter_req_0); -- 
    merge_ack_12890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2578_gather_scatter_ack_0, ack => cp_elements(138)); -- 
    cpelement_group_139 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(140) & cp_elements(141));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(139),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => type_cast_2582_inst_req_0); -- 
    cp_elements(140) <= cp_elements(0);
    cp_elements(141) <= cp_elements(17);
    ack_12900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_0, ack => cp_elements(142)); -- 
    base_resize_req_12911_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => array_obj_ref_2587_base_resize_req_0); -- 
    cp_elements(143) <= cp_elements(0);
    cpelement_group_144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(147));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => array_obj_ref_2587_final_reg_req_0); -- 
    base_resize_ack_12912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2587_base_resize_ack_0, ack => cp_elements(145)); -- 
    plus_base_rr_12917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => array_obj_ref_2587_root_address_inst_req_0); -- 
    plus_base_ra_12918_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2587_root_address_inst_ack_0, ack => cp_elements(146)); -- 
    plus_base_cr_12919_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(146), ack => array_obj_ref_2587_root_address_inst_req_1); -- 
    plus_base_ca_12920_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2587_root_address_inst_ack_1, ack => cp_elements(147)); -- 
    cp_elements(148) <= array_obj_ref_2587_final_reg_ack_0;
    cpelement_group_149 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(159));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(149),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(150) <= cp_elements(148);
    base_resize_req_12938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(150), ack => ptr_deref_2591_base_resize_req_0); -- 
    base_resize_ack_12939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_base_resize_ack_0, ack => cp_elements(151)); -- 
    sum_rename_req_12943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2591_root_address_inst_req_0); -- 
    cp_elements(152) <= ptr_deref_2591_root_address_inst_ack_0;
    cp_elements(153) <= cp_elements(152);
    rr_12951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2591_addr_0_req_0); -- 
    ra_12952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_addr_0_ack_0, ack => cp_elements(154)); -- 
    cr_12953_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => ptr_deref_2591_addr_0_req_1); -- 
    ca_12954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_addr_0_ack_1, ack => cp_elements(155)); -- 
    cp_elements(156) <= cp_elements(152);
    rr_12958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => ptr_deref_2591_addr_1_req_0); -- 
    ra_12959_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_addr_1_ack_0, ack => cp_elements(157)); -- 
    cr_12960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => ptr_deref_2591_addr_1_req_1); -- 
    ca_12961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_addr_1_ack_1, ack => cp_elements(158)); -- 
    cpelement_group_159 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(155) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(159),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(160) <= cp_elements(149);
    rr_12971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => ptr_deref_2591_load_0_req_0); -- 
    ra_12972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_load_0_ack_0, ack => cp_elements(161)); -- 
    cp_elements(162) <= cp_elements(149);
    rr_12976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => ptr_deref_2591_load_1_req_0); -- 
    ra_12977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_load_1_ack_0, ack => cp_elements(163)); -- 
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(161) & cp_elements(163));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(165) <= cp_elements(164);
    cr_12987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => ptr_deref_2591_load_0_req_1); -- 
    ca_12988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_load_0_ack_1, ack => cp_elements(166)); -- 
    cp_elements(167) <= cp_elements(164);
    cr_12992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => ptr_deref_2591_load_1_req_1); -- 
    ca_12993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_load_1_ack_1, ack => cp_elements(168)); -- 
    cpelement_group_169 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(166) & cp_elements(168));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(169),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => ptr_deref_2591_gather_scatter_req_0); -- 
    merge_ack_12995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2591_gather_scatter_ack_0, ack => cp_elements(170)); -- 
    cpelement_group_171 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(170) & cp_elements(172));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(171),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => type_cast_2595_inst_req_0); -- 
    cp_elements(172) <= cp_elements(0);
    ack_13005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2595_inst_ack_0, ack => cp_elements(173)); -- 
    cpelement_group_174 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(173) & cp_elements(175));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(174),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(174), ack => binary_2601_inst_req_0); -- 
    cp_elements(175) <= cp_elements(0);
    ra_13015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2601_inst_ack_0, ack => cp_elements(176)); -- 
    cr_13016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2601_inst_req_1); -- 
    ca_13017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2601_inst_ack_1, ack => cp_elements(177)); -- 
    cpelement_group_178 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(138) & cp_elements(179));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(178),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => type_cast_2605_inst_req_0); -- 
    cp_elements(179) <= cp_elements(0);
    ack_13027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2605_inst_ack_0, ack => cp_elements(180)); -- 
    cpelement_group_181 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(182) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(181),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => type_cast_2614_inst_req_0); -- 
    cp_elements(182) <= cp_elements(0);
    cpelement_group_183 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(187));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(183),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2613_inst_req_0); -- 
    cp_elements(184) <= cp_elements(0);
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(180) & cp_elements(186));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => type_cast_2609_inst_req_0); -- 
    cp_elements(186) <= cp_elements(0);
    ack_13041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_0, ack => cp_elements(187)); -- 
    ra_13046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2613_inst_ack_0, ack => cp_elements(188)); -- 
    cr_13047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => binary_2613_inst_req_1); -- 
    ca_13048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2613_inst_ack_1, ack => cp_elements(189)); -- 
    ack_13053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_0, ack => cp_elements(190)); -- 
    cpelement_group_191 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(177) & cp_elements(190) & cp_elements(192));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(191),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => binary_2619_inst_req_0); -- 
    cp_elements(192) <= cp_elements(0);
    ra_13064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2619_inst_ack_0, ack => cp_elements(193)); -- 
    cr_13065_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => binary_2619_inst_req_1); -- 
    ca_13066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2619_inst_ack_1, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => type_cast_2623_inst_req_0); -- 
    cp_elements(196) <= cp_elements(0);
    ack_13076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2623_inst_ack_0, ack => cp_elements(197)); -- 
    cpelement_group_198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(106) & cp_elements(197));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addx_xptr16_2530 : std_logic_vector(31 downto 0);
    signal addx_xptr25_2575 : std_logic_vector(31 downto 0);
    signal addx_xptr29_2588 : std_logic_vector(31 downto 0);
    signal addx_xptr_2517 : std_logic_vector(31 downto 0);
    signal and_2501 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2516_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2516_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2516_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2529_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2529_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2529_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2574_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2574_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2574_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2587_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2587_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2587_root_address : std_logic_vector(15 downto 0);
    signal binary_2555_wire : std_logic_vector(31 downto 0);
    signal binary_2613_wire : std_logic_vector(31 downto 0);
    signal blen_h_2579 : std_logic_vector(15 downto 0);
    signal blen_l_2592 : std_logic_vector(15 downto 0);
    signal conv21_2548 : std_logic_vector(31 downto 0);
    signal conv33_2596 : std_logic_vector(31 downto 0);
    signal conv36_2606 : std_logic_vector(31 downto 0);
    signal conv_2538 : std_logic_vector(31 downto 0);
    signal iNsTr_11_2525 : std_logic_vector(31 downto 0);
    signal iNsTr_14_2570 : std_logic_vector(31 downto 0);
    signal iNsTr_16_2583 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2495 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2505 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2509 : std_logic_vector(31 downto 0);
    signal or38_2620 : std_logic_vector(31 downto 0);
    signal or_2562 : std_logic_vector(31 downto 0);
    signal ptr_deref_2520_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2520_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2520_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2520_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2520_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2520_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2520_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2520_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2533_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2533_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2533_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2533_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2533_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2533_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2533_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2533_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2578_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2578_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2578_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2578_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2578_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2578_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2578_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2578_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2591_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2591_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2591_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2591_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2591_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2591_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2591_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2591_word_offset_1 : std_logic_vector(15 downto 0);
    signal shl34_2602 : std_logic_vector(31 downto 0);
    signal shl_2544 : std_logic_vector(31 downto 0);
    signal shr37_2615 : std_logic_vector(31 downto 0);
    signal shr_2557 : std_logic_vector(31 downto 0);
    signal type_cast_2499_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2542_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2551_wire : std_logic_vector(31 downto 0);
    signal type_cast_2554_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2600_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2609_wire : std_logic_vector(31 downto 0);
    signal type_cast_2612_wire_constant : std_logic_vector(31 downto 0);
    signal wlen_h_2521 : std_logic_vector(15 downto 0);
    signal wlen_l_2534 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2516_final_offset <= "0000000000000010";
    array_obj_ref_2529_final_offset <= "0000000000000010";
    array_obj_ref_2574_final_offset <= "0000000000000110";
    array_obj_ref_2587_final_offset <= "0000000000000110";
    ptr_deref_2520_word_offset_0 <= "0000000000000000";
    ptr_deref_2520_word_offset_1 <= "0000000000000001";
    ptr_deref_2533_word_offset_0 <= "0000000000000000";
    ptr_deref_2533_word_offset_1 <= "0000000000000001";
    ptr_deref_2578_word_offset_0 <= "0000000000000000";
    ptr_deref_2578_word_offset_1 <= "0000000000000001";
    ptr_deref_2591_word_offset_0 <= "0000000000000000";
    ptr_deref_2591_word_offset_1 <= "0000000000000001";
    type_cast_2499_wire_constant <= "11111111111111111111100000000000";
    type_cast_2542_wire_constant <= "00000000000000000000000000001000";
    type_cast_2554_wire_constant <= "00000000000000000000000000001000";
    type_cast_2600_wire_constant <= "00000000000000000000000000001000";
    type_cast_2612_wire_constant <= "00000000000000000000000000001000";
    array_obj_ref_2516_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_9_2509, dout => array_obj_ref_2516_resized_base_address, req => array_obj_ref_2516_base_resize_req_0, ack => array_obj_ref_2516_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2516_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2516_root_address, dout => addx_xptr_2517, req => array_obj_ref_2516_final_reg_req_0, ack => array_obj_ref_2516_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2529_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_11_2525, dout => array_obj_ref_2529_resized_base_address, req => array_obj_ref_2529_base_resize_req_0, ack => array_obj_ref_2529_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2529_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2529_root_address, dout => addx_xptr16_2530, req => array_obj_ref_2529_final_reg_req_0, ack => array_obj_ref_2529_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2574_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_14_2570, dout => array_obj_ref_2574_resized_base_address, req => array_obj_ref_2574_base_resize_req_0, ack => array_obj_ref_2574_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2574_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2574_root_address, dout => addx_xptr25_2575, req => array_obj_ref_2574_final_reg_req_0, ack => array_obj_ref_2574_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2587_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_16_2583, dout => array_obj_ref_2587_resized_base_address, req => array_obj_ref_2587_base_resize_req_0, ack => array_obj_ref_2587_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2587_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2587_root_address, dout => addx_xptr29_2588, req => array_obj_ref_2587_final_reg_req_0, ack => array_obj_ref_2587_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2520_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr_2517, dout => ptr_deref_2520_resized_base_address, req => ptr_deref_2520_base_resize_req_0, ack => ptr_deref_2520_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2533_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr16_2530, dout => ptr_deref_2533_resized_base_address, req => ptr_deref_2533_base_resize_req_0, ack => ptr_deref_2533_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2578_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr25_2575, dout => ptr_deref_2578_resized_base_address, req => ptr_deref_2578_base_resize_req_0, ack => ptr_deref_2578_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2591_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr29_2588, dout => ptr_deref_2591_resized_base_address, req => ptr_deref_2591_base_resize_req_0, ack => ptr_deref_2591_base_resize_ack_0, clk => clk, reset => reset); -- 
    simple_obj_ref_2510_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_7_2505, dout => buf_buffer, req => simple_obj_ref_2510_inst_req_0, ack => simple_obj_ref_2510_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2494_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => pkt, dout => iNsTr_6_2495, req => type_cast_2494_inst_req_0, ack => type_cast_2494_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2504_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => and_2501, dout => iNsTr_7_2505, req => type_cast_2504_inst_req_0, ack => type_cast_2504_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2508_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => and_2501, dout => iNsTr_9_2509, req => type_cast_2508_inst_req_0, ack => type_cast_2508_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2524_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_buffer, dout => iNsTr_11_2525, req => type_cast_2524_inst_req_0, ack => type_cast_2524_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2537_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => wlen_l_2534, dout => conv_2538, req => type_cast_2537_inst_req_0, ack => type_cast_2537_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2547_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => wlen_h_2521, dout => conv21_2548, req => type_cast_2547_inst_req_0, ack => type_cast_2547_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2551_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => conv21_2548, dout => type_cast_2551_wire, req => type_cast_2551_inst_req_0, ack => type_cast_2551_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2556_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => binary_2555_wire, dout => shr_2557, req => type_cast_2556_inst_req_0, ack => type_cast_2556_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2565_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => or_2562, dout => wlen_buffer, req => type_cast_2565_inst_req_0, ack => type_cast_2565_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2569_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_buffer, dout => iNsTr_14_2570, req => type_cast_2569_inst_req_0, ack => type_cast_2569_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2582_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_buffer, dout => iNsTr_16_2583, req => type_cast_2582_inst_req_0, ack => type_cast_2582_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2595_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => blen_l_2592, dout => conv33_2596, req => type_cast_2595_inst_req_0, ack => type_cast_2595_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2605_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => blen_h_2579, dout => conv36_2606, req => type_cast_2605_inst_req_0, ack => type_cast_2605_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2609_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => conv36_2606, dout => type_cast_2609_wire, req => type_cast_2609_inst_req_0, ack => type_cast_2609_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2614_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => binary_2613_wire, dout => shr37_2615, req => type_cast_2614_inst_req_0, ack => type_cast_2614_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2623_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => or38_2620, dout => blen_buffer, req => type_cast_2623_inst_req_0, ack => type_cast_2623_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2520_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2520_gather_scatter_ack_0 <= ptr_deref_2520_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2520_data_1 & ptr_deref_2520_data_0;
      wlen_h_2521 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2520_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2520_root_address_inst_ack_0 <= ptr_deref_2520_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2520_resized_base_address;
      ptr_deref_2520_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2533_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2533_gather_scatter_ack_0 <= ptr_deref_2533_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2533_data_1 & ptr_deref_2533_data_0;
      wlen_l_2534 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2533_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2533_root_address_inst_ack_0 <= ptr_deref_2533_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2533_resized_base_address;
      ptr_deref_2533_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2578_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2578_gather_scatter_ack_0 <= ptr_deref_2578_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2578_data_1 & ptr_deref_2578_data_0;
      blen_h_2579 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2578_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2578_root_address_inst_ack_0 <= ptr_deref_2578_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2578_resized_base_address;
      ptr_deref_2578_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2591_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2591_gather_scatter_ack_0 <= ptr_deref_2591_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2591_data_1 & ptr_deref_2591_data_0;
      blen_l_2592 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2591_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2591_root_address_inst_ack_0 <= ptr_deref_2591_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2591_resized_base_address;
      ptr_deref_2591_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2516_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2516_resized_base_address;
      array_obj_ref_2516_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2516_root_address_inst_req_0,
          ackL => array_obj_ref_2516_root_address_inst_ack_0,
          reqR => array_obj_ref_2516_root_address_inst_req_1,
          ackR => array_obj_ref_2516_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2529_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2529_resized_base_address;
      array_obj_ref_2529_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2529_root_address_inst_req_0,
          ackL => array_obj_ref_2529_root_address_inst_ack_0,
          reqR => array_obj_ref_2529_root_address_inst_req_1,
          ackR => array_obj_ref_2529_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_2574_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2574_resized_base_address;
      array_obj_ref_2574_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2574_root_address_inst_req_0,
          ackL => array_obj_ref_2574_root_address_inst_ack_0,
          reqR => array_obj_ref_2574_root_address_inst_req_1,
          ackR => array_obj_ref_2574_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_2587_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2587_resized_base_address;
      array_obj_ref_2587_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2587_root_address_inst_req_0,
          ackL => array_obj_ref_2587_root_address_inst_ack_0,
          reqR => array_obj_ref_2587_root_address_inst_req_1,
          ackR => array_obj_ref_2587_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2500_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_6_2495;
      and_2501 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2500_inst_req_0,
          ackL => binary_2500_inst_ack_0,
          reqR => binary_2500_inst_req_1,
          ackR => binary_2500_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2543_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= conv_2538;
      shl_2544 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2543_inst_req_0,
          ackL => binary_2543_inst_ack_0,
          reqR => binary_2543_inst_req_1,
          ackR => binary_2543_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2555_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2551_wire;
      binary_2555_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntASHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2555_inst_req_0,
          ackL => binary_2555_inst_ack_0,
          reqR => binary_2555_inst_req_1,
          ackR => binary_2555_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2561_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= shl_2544 & shr_2557;
      or_2562 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2561_inst_req_0,
          ackL => binary_2561_inst_ack_0,
          reqR => binary_2561_inst_req_1,
          ackR => binary_2561_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2601_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= conv33_2596;
      shl34_2602 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2601_inst_req_0,
          ackL => binary_2601_inst_ack_0,
          reqR => binary_2601_inst_req_1,
          ackR => binary_2601_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2613_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2609_wire;
      binary_2613_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntASHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2613_inst_req_0,
          ackL => binary_2613_inst_ack_0,
          reqR => binary_2613_inst_req_1,
          ackR => binary_2613_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2619_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= shl34_2602 & shr37_2615;
      or38_2620 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2619_inst_req_0,
          ackL => binary_2619_inst_ack_0,
          reqR => binary_2619_inst_req_1,
          ackR => binary_2619_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2520_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2520_root_address;
      ptr_deref_2520_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2520_addr_0_req_0,
          ackL => ptr_deref_2520_addr_0_ack_0,
          reqR => ptr_deref_2520_addr_0_req_1,
          ackR => ptr_deref_2520_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2520_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2520_root_address;
      ptr_deref_2520_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2520_addr_1_req_0,
          ackL => ptr_deref_2520_addr_1_ack_0,
          reqR => ptr_deref_2520_addr_1_req_1,
          ackR => ptr_deref_2520_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2533_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2533_root_address;
      ptr_deref_2533_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2533_addr_0_req_0,
          ackL => ptr_deref_2533_addr_0_ack_0,
          reqR => ptr_deref_2533_addr_0_req_1,
          ackR => ptr_deref_2533_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2533_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2533_root_address;
      ptr_deref_2533_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2533_addr_1_req_0,
          ackL => ptr_deref_2533_addr_1_ack_0,
          reqR => ptr_deref_2533_addr_1_req_1,
          ackR => ptr_deref_2533_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2578_addr_0 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2578_root_address;
      ptr_deref_2578_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2578_addr_0_req_0,
          ackL => ptr_deref_2578_addr_0_ack_0,
          reqR => ptr_deref_2578_addr_0_req_1,
          ackR => ptr_deref_2578_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2578_addr_1 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2578_root_address;
      ptr_deref_2578_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2578_addr_1_req_0,
          ackL => ptr_deref_2578_addr_1_ack_0,
          reqR => ptr_deref_2578_addr_1_req_1,
          ackR => ptr_deref_2578_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2591_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2591_root_address;
      ptr_deref_2591_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2591_addr_0_req_0,
          ackL => ptr_deref_2591_addr_0_ack_0,
          reqR => ptr_deref_2591_addr_0_req_1,
          ackR => ptr_deref_2591_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2591_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2591_root_address;
      ptr_deref_2591_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2591_addr_1_req_0,
          ackL => ptr_deref_2591_addr_1_ack_0,
          reqR => ptr_deref_2591_addr_1_req_1,
          ackR => ptr_deref_2591_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared load operator group (0) : ptr_deref_2591_load_1 ptr_deref_2520_load_0 ptr_deref_2533_load_1 ptr_deref_2533_load_0 ptr_deref_2520_load_1 ptr_deref_2591_load_0 ptr_deref_2578_load_0 ptr_deref_2578_load_1 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2591_load_1_req_0,
        ptr_deref_2591_load_1_ack_0,
        ptr_deref_2591_load_1_req_1,
        ptr_deref_2591_load_1_ack_1,
        "ptr_deref_2591_load_1",
        "memory_space_5" ,
        ptr_deref_2591_data_1,
        ptr_deref_2591_word_address_1,
        "ptr_deref_2591_data_1",
        "ptr_deref_2591_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2520_load_0_req_0,
        ptr_deref_2520_load_0_ack_0,
        ptr_deref_2520_load_0_req_1,
        ptr_deref_2520_load_0_ack_1,
        "ptr_deref_2520_load_0",
        "memory_space_5" ,
        ptr_deref_2520_data_0,
        ptr_deref_2520_word_address_0,
        "ptr_deref_2520_data_0",
        "ptr_deref_2520_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2533_load_1_req_0,
        ptr_deref_2533_load_1_ack_0,
        ptr_deref_2533_load_1_req_1,
        ptr_deref_2533_load_1_ack_1,
        "ptr_deref_2533_load_1",
        "memory_space_5" ,
        ptr_deref_2533_data_1,
        ptr_deref_2533_word_address_1,
        "ptr_deref_2533_data_1",
        "ptr_deref_2533_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2533_load_0_req_0,
        ptr_deref_2533_load_0_ack_0,
        ptr_deref_2533_load_0_req_1,
        ptr_deref_2533_load_0_ack_1,
        "ptr_deref_2533_load_0",
        "memory_space_5" ,
        ptr_deref_2533_data_0,
        ptr_deref_2533_word_address_0,
        "ptr_deref_2533_data_0",
        "ptr_deref_2533_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2520_load_1_req_0,
        ptr_deref_2520_load_1_ack_0,
        ptr_deref_2520_load_1_req_1,
        ptr_deref_2520_load_1_ack_1,
        "ptr_deref_2520_load_1",
        "memory_space_5" ,
        ptr_deref_2520_data_1,
        ptr_deref_2520_word_address_1,
        "ptr_deref_2520_data_1",
        "ptr_deref_2520_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2591_load_0_req_0,
        ptr_deref_2591_load_0_ack_0,
        ptr_deref_2591_load_0_req_1,
        ptr_deref_2591_load_0_ack_1,
        "ptr_deref_2591_load_0",
        "memory_space_5" ,
        ptr_deref_2591_data_0,
        ptr_deref_2591_word_address_0,
        "ptr_deref_2591_data_0",
        "ptr_deref_2591_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2578_load_0_req_0,
        ptr_deref_2578_load_0_ack_0,
        ptr_deref_2578_load_0_req_1,
        ptr_deref_2578_load_0_ack_1,
        "ptr_deref_2578_load_0",
        "memory_space_5" ,
        ptr_deref_2578_data_0,
        ptr_deref_2578_word_address_0,
        "ptr_deref_2578_data_0",
        "ptr_deref_2578_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2578_load_1_req_0,
        ptr_deref_2578_load_1_ack_0,
        ptr_deref_2578_load_1_req_1,
        ptr_deref_2578_load_1_ack_1,
        "ptr_deref_2578_load_1",
        "memory_space_5" ,
        ptr_deref_2578_data_1,
        ptr_deref_2578_word_address_1,
        "ptr_deref_2578_data_1",
        "ptr_deref_2578_word_address_1" -- 
      );
      reqL(7) <= ptr_deref_2591_load_1_req_0;
      reqL(6) <= ptr_deref_2520_load_0_req_0;
      reqL(5) <= ptr_deref_2533_load_1_req_0;
      reqL(4) <= ptr_deref_2533_load_0_req_0;
      reqL(3) <= ptr_deref_2520_load_1_req_0;
      reqL(2) <= ptr_deref_2591_load_0_req_0;
      reqL(1) <= ptr_deref_2578_load_0_req_0;
      reqL(0) <= ptr_deref_2578_load_1_req_0;
      ptr_deref_2591_load_1_ack_0 <= ackL(7);
      ptr_deref_2520_load_0_ack_0 <= ackL(6);
      ptr_deref_2533_load_1_ack_0 <= ackL(5);
      ptr_deref_2533_load_0_ack_0 <= ackL(4);
      ptr_deref_2520_load_1_ack_0 <= ackL(3);
      ptr_deref_2591_load_0_ack_0 <= ackL(2);
      ptr_deref_2578_load_0_ack_0 <= ackL(1);
      ptr_deref_2578_load_1_ack_0 <= ackL(0);
      reqR(7) <= ptr_deref_2591_load_1_req_1;
      reqR(6) <= ptr_deref_2520_load_0_req_1;
      reqR(5) <= ptr_deref_2533_load_1_req_1;
      reqR(4) <= ptr_deref_2533_load_0_req_1;
      reqR(3) <= ptr_deref_2520_load_1_req_1;
      reqR(2) <= ptr_deref_2591_load_0_req_1;
      reqR(1) <= ptr_deref_2578_load_0_req_1;
      reqR(0) <= ptr_deref_2578_load_1_req_1;
      ptr_deref_2591_load_1_ack_1 <= ackR(7);
      ptr_deref_2520_load_0_ack_1 <= ackR(6);
      ptr_deref_2533_load_1_ack_1 <= ackR(5);
      ptr_deref_2533_load_0_ack_1 <= ackR(4);
      ptr_deref_2520_load_1_ack_1 <= ackR(3);
      ptr_deref_2591_load_0_ack_1 <= ackR(2);
      ptr_deref_2578_load_0_ack_1 <= ackR(1);
      ptr_deref_2578_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_2591_word_address_1 & ptr_deref_2520_word_address_0 & ptr_deref_2533_word_address_1 & ptr_deref_2533_word_address_0 & ptr_deref_2520_word_address_1 & ptr_deref_2591_word_address_0 & ptr_deref_2578_word_address_0 & ptr_deref_2578_word_address_1;
      ptr_deref_2591_data_1 <= data_out(63 downto 56);
      ptr_deref_2520_data_0 <= data_out(55 downto 48);
      ptr_deref_2533_data_1 <= data_out(47 downto 40);
      ptr_deref_2533_data_0 <= data_out(39 downto 32);
      ptr_deref_2520_data_1 <= data_out(31 downto 24);
      ptr_deref_2591_data_0 <= data_out(23 downto 16);
      ptr_deref_2578_data_0 <= data_out(15 downto 8);
      ptr_deref_2578_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 8,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 8,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity click_bc_storage_initializer_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    GV_15_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity click_bc_storage_initializer_x;
architecture Default of click_bc_storage_initializer_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal click_bc_storage_initializer_x_xCP_13077_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_2628_call_req_0 : boolean;
  signal call_stmt_2628_call_ack_0 : boolean;
  signal call_stmt_2628_call_req_1 : boolean;
  signal call_stmt_2628_call_ack_1 : boolean;
  signal call_stmt_2629_call_req_0 : boolean;
  signal call_stmt_2629_call_ack_0 : boolean;
  signal call_stmt_2629_call_req_1 : boolean;
  signal call_stmt_2629_call_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  click_bc_storage_initializer_x_xCP_13077: Block -- control-path 
    signal cp_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(7);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(7), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    crr_13091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2628_call_req_0); -- 
    cra_13092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2628_call_ack_0, ack => cp_elements(2)); -- 
    ccr_13096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2628_call_req_1); -- 
    cca_13097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2628_call_ack_1, ack => cp_elements(3)); -- 
    cp_elements(4) <= cp_elements(0);
    crr_13108_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => call_stmt_2629_call_req_0); -- 
    cra_13109_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2629_call_ack_0, ack => cp_elements(5)); -- 
    ccr_13113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => call_stmt_2629_call_req_1); -- 
    cca_13114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2629_call_ack_1, ack => cp_elements(6)); -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(6));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_2628_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_2628_call_req_0;
      call_stmt_2628_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_2628_call_req_1;
      call_stmt_2628_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => GV_15_initializer_in_click_bc_call_reqs(0),
          ackR => GV_15_initializer_in_click_bc_call_acks(0),
          tagR => GV_15_initializer_in_click_bc_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => GV_15_initializer_in_click_bc_return_acks(0), -- cross-over
          ackL => GV_15_initializer_in_click_bc_return_reqs(0), -- cross-over
          tagL => GV_15_initializer_in_click_bc_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2629_call 
    CallGroup1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_2629_call_req_0;
      call_stmt_2629_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_2629_call_req_1;
      call_stmt_2629_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => GV_16_initializer_in_click_bc_call_reqs(0),
          ackR => GV_16_initializer_in_click_bc_call_acks(0),
          tagR => GV_16_initializer_in_click_bc_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => GV_16_initializer_in_click_bc_return_acks(0), -- cross-over
          ackL => GV_16_initializer_in_click_bc_return_reqs(0), -- cross-over
          tagL => GV_16_initializer_in_click_bc_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_init is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity free_queue_init;
architecture Default of free_queue_init is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal free_queue_init_CP_13117_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_2640_base_resize_req_0 : boolean;
  signal ptr_deref_2640_base_resize_ack_0 : boolean;
  signal ptr_deref_2640_root_address_inst_req_0 : boolean;
  signal ptr_deref_2640_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2640_addr_0_req_0 : boolean;
  signal ptr_deref_2640_addr_0_ack_0 : boolean;
  signal ptr_deref_2640_gather_scatter_req_0 : boolean;
  signal ptr_deref_2640_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2640_store_0_req_0 : boolean;
  signal ptr_deref_2640_store_0_ack_0 : boolean;
  signal ptr_deref_2640_store_0_req_1 : boolean;
  signal ptr_deref_2640_store_0_ack_1 : boolean;
  signal ptr_deref_2648_base_resize_req_0 : boolean;
  signal ptr_deref_2648_base_resize_ack_0 : boolean;
  signal ptr_deref_2648_root_address_inst_req_0 : boolean;
  signal ptr_deref_2648_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2648_addr_0_req_0 : boolean;
  signal ptr_deref_2648_addr_0_ack_0 : boolean;
  signal ptr_deref_2648_load_0_req_0 : boolean;
  signal ptr_deref_2648_load_0_ack_0 : boolean;
  signal ptr_deref_2648_load_0_req_1 : boolean;
  signal ptr_deref_2648_load_0_ack_1 : boolean;
  signal ptr_deref_2648_gather_scatter_req_0 : boolean;
  signal ptr_deref_2648_gather_scatter_ack_0 : boolean;
  signal type_cast_2652_inst_req_0 : boolean;
  signal type_cast_2652_inst_ack_0 : boolean;
  signal binary_2656_inst_req_0 : boolean;
  signal binary_2656_inst_ack_0 : boolean;
  signal binary_2656_inst_req_1 : boolean;
  signal binary_2656_inst_ack_1 : boolean;
  signal if_stmt_2658_branch_req_0 : boolean;
  signal if_stmt_2658_branch_ack_1 : boolean;
  signal if_stmt_2658_branch_ack_0 : boolean;
  signal ptr_deref_2667_base_resize_req_0 : boolean;
  signal ptr_deref_2667_base_resize_ack_0 : boolean;
  signal ptr_deref_2667_root_address_inst_req_0 : boolean;
  signal ptr_deref_2667_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2667_addr_0_req_0 : boolean;
  signal ptr_deref_2667_addr_0_ack_0 : boolean;
  signal ptr_deref_2667_load_0_req_0 : boolean;
  signal ptr_deref_2667_load_0_ack_0 : boolean;
  signal ptr_deref_2667_load_0_req_1 : boolean;
  signal ptr_deref_2667_load_0_ack_1 : boolean;
  signal ptr_deref_2667_gather_scatter_req_0 : boolean;
  signal ptr_deref_2667_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2671_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2671_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2671_index_0_scale_req_0 : boolean;
  signal array_obj_ref_2671_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_2671_index_0_scale_req_1 : boolean;
  signal array_obj_ref_2671_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_2671_offset_inst_req_0 : boolean;
  signal array_obj_ref_2671_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2671_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2671_root_address_inst_ack_0 : boolean;
  signal addr_of_2672_final_reg_req_0 : boolean;
  signal addr_of_2672_final_reg_ack_0 : boolean;
  signal array_obj_ref_2679_base_resize_req_0 : boolean;
  signal array_obj_ref_2679_base_resize_ack_0 : boolean;
  signal array_obj_ref_2679_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2679_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2679_final_reg_req_0 : boolean;
  signal array_obj_ref_2679_final_reg_ack_0 : boolean;
  signal array_obj_ref_2686_base_resize_req_0 : boolean;
  signal array_obj_ref_2686_base_resize_ack_0 : boolean;
  signal array_obj_ref_2686_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2686_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2686_final_reg_req_0 : boolean;
  signal array_obj_ref_2686_final_reg_ack_0 : boolean;
  signal type_cast_2690_inst_req_0 : boolean;
  signal type_cast_2690_inst_ack_0 : boolean;
  signal simple_obj_ref_2692_inst_req_0 : boolean;
  signal simple_obj_ref_2692_inst_ack_0 : boolean;
  signal ptr_deref_2699_base_resize_req_0 : boolean;
  signal ptr_deref_2699_base_resize_ack_0 : boolean;
  signal ptr_deref_2699_root_address_inst_req_0 : boolean;
  signal ptr_deref_2699_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2699_addr_0_req_0 : boolean;
  signal ptr_deref_2699_addr_0_ack_0 : boolean;
  signal ptr_deref_2699_load_0_req_0 : boolean;
  signal ptr_deref_2699_load_0_ack_0 : boolean;
  signal ptr_deref_2699_load_0_req_1 : boolean;
  signal ptr_deref_2699_load_0_ack_1 : boolean;
  signal ptr_deref_2699_gather_scatter_req_0 : boolean;
  signal ptr_deref_2699_gather_scatter_ack_0 : boolean;
  signal binary_2705_inst_req_0 : boolean;
  signal binary_2705_inst_ack_0 : boolean;
  signal binary_2705_inst_req_1 : boolean;
  signal binary_2705_inst_ack_1 : boolean;
  signal ptr_deref_2708_base_resize_req_0 : boolean;
  signal ptr_deref_2708_base_resize_ack_0 : boolean;
  signal ptr_deref_2708_root_address_inst_req_0 : boolean;
  signal ptr_deref_2708_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2708_addr_0_req_0 : boolean;
  signal ptr_deref_2708_addr_0_ack_0 : boolean;
  signal ptr_deref_2708_gather_scatter_req_0 : boolean;
  signal ptr_deref_2708_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2708_store_0_req_0 : boolean;
  signal ptr_deref_2708_store_0_ack_0 : boolean;
  signal ptr_deref_2708_store_0_req_1 : boolean;
  signal ptr_deref_2708_store_0_ack_1 : boolean;
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(1 downto 0);
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  free_queue_init_CP_13117: Block -- control-path 
    signal cp_elements: BooleanArray(98 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(38);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(38), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(36) & cp_elements(98));
    cp_elements(2) <= cp_elements(0);
    cp_elements(3) <= cp_elements(2);
    cpelement_group_4 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(5) & cp_elements(9));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(4),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_13177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => ptr_deref_2640_gather_scatter_req_0); -- 
    cp_elements(5) <= cp_elements(2);
    cp_elements(6) <= cp_elements(5);
    base_resize_req_13162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => ptr_deref_2640_base_resize_req_0); -- 
    base_resize_ack_13163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_base_resize_ack_0, ack => cp_elements(7)); -- 
    sum_rename_req_13167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_2640_root_address_inst_req_0); -- 
    sum_rename_ack_13168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_root_address_inst_ack_0, ack => cp_elements(8)); -- 
    root_rename_req_13172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => ptr_deref_2640_addr_0_req_0); -- 
    root_rename_ack_13173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_addr_0_ack_0, ack => cp_elements(9)); -- 
    split_ack_13178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_gather_scatter_ack_0, ack => cp_elements(10)); -- 
    rr_13185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_2640_store_0_req_0); -- 
    ra_13186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_store_0_ack_0, ack => cp_elements(11)); -- 
    cr_13196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => ptr_deref_2640_store_0_req_1); -- 
    ca_13197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_store_0_ack_1, ack => cp_elements(12)); -- 
    cp_elements(13) <= cp_elements(96);
    cpelement_group_14 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(15) & cp_elements(19));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(14),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13234_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => ptr_deref_2648_load_0_req_0); -- 
    cp_elements(15) <= cp_elements(13);
    cp_elements(16) <= cp_elements(15);
    base_resize_req_13213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_2648_base_resize_req_0); -- 
    base_resize_ack_13214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_base_resize_ack_0, ack => cp_elements(17)); -- 
    sum_rename_req_13218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_2648_root_address_inst_req_0); -- 
    sum_rename_ack_13219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_root_address_inst_ack_0, ack => cp_elements(18)); -- 
    root_rename_req_13223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_2648_addr_0_req_0); -- 
    root_rename_ack_13224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_addr_0_ack_0, ack => cp_elements(19)); -- 
    ra_13235_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_load_0_ack_0, ack => cp_elements(20)); -- 
    cr_13245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_2648_load_0_req_1); -- 
    ca_13246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_load_0_ack_1, ack => cp_elements(21)); -- 
    merge_req_13247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => ptr_deref_2648_gather_scatter_req_0); -- 
    merge_ack_13248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(24) & cp_elements(27));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => binary_2656_inst_req_0); -- 
    cp_elements(24) <= cp_elements(13);
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(26));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13259_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => type_cast_2652_inst_req_0); -- 
    cp_elements(26) <= cp_elements(13);
    ack_13260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2652_inst_ack_0, ack => cp_elements(27)); -- 
    ra_13265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2656_inst_ack_0, ack => cp_elements(28)); -- 
    cr_13266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => binary_2656_inst_req_1); -- 
    ca_13267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2656_inst_ack_1, ack => cp_elements(29)); -- 
    cp_elements(30) <= cp_elements(29);
    cp_elements(31) <= false;
    cp_elements(32) <= cp_elements(31);
    cp_elements(33) <= cp_elements(29);
    branch_req_13275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => if_stmt_2658_branch_req_0); -- 
    cp_elements(34) <= cp_elements(33);
    cp_elements(35) <= cp_elements(34);
    if_choice_transition_13280_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2658_branch_ack_1, ack => cp_elements(36)); -- 
    cp_elements(37) <= cp_elements(34);
    else_choice_transition_13284_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2658_branch_ack_0, ack => cp_elements(38)); -- 
    cp_elements(39) <= cp_elements(1);
    cpelement_group_40 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(41) & cp_elements(45));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(40),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_2667_load_0_req_0); -- 
    cp_elements(41) <= cp_elements(39);
    cp_elements(42) <= cp_elements(41);
    base_resize_req_13302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_2667_base_resize_req_0); -- 
    base_resize_ack_13303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_base_resize_ack_0, ack => cp_elements(43)); -- 
    sum_rename_req_13307_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2667_root_address_inst_req_0); -- 
    sum_rename_ack_13308_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_root_address_inst_ack_0, ack => cp_elements(44)); -- 
    root_rename_req_13312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_2667_addr_0_req_0); -- 
    root_rename_ack_13313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_addr_0_ack_0, ack => cp_elements(45)); -- 
    ra_13324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_load_0_ack_0, ack => cp_elements(46)); -- 
    cr_13334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_2667_load_0_req_1); -- 
    ca_13335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_load_0_ack_1, ack => cp_elements(47)); -- 
    merge_req_13336_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2667_gather_scatter_req_0); -- 
    merge_ack_13337_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_gather_scatter_ack_0, ack => cp_elements(48)); -- 
    index_resize_req_13351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => array_obj_ref_2671_index_0_resize_req_0); -- 
    cpelement_group_49 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(55));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(49),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_13373_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => addr_of_2672_final_reg_req_0); -- 
    cp_elements(50) <= cp_elements(39);
    index_resize_ack_13352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_index_0_resize_ack_0, ack => cp_elements(51)); -- 
    scale_rr_13356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_2671_index_0_scale_req_0); -- 
    scale_ra_13357_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_index_0_scale_ack_0, ack => cp_elements(52)); -- 
    scale_cr_13358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => array_obj_ref_2671_index_0_scale_req_1); -- 
    scale_ca_13359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_index_0_scale_ack_1, ack => cp_elements(53)); -- 
    final_index_req_13363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_2671_offset_inst_req_0); -- 
    final_index_ack_13364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_offset_inst_ack_0, ack => cp_elements(54)); -- 
    sum_rename_req_13368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => array_obj_ref_2671_root_address_inst_req_0); -- 
    sum_rename_ack_13369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_root_address_inst_ack_0, ack => cp_elements(55)); -- 
    final_reg_ack_13374_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2672_final_reg_ack_0, ack => cp_elements(56)); -- 
    base_resize_req_13385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => array_obj_ref_2679_base_resize_req_0); -- 
    cp_elements(57) <= cp_elements(39);
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(57) & cp_elements(60));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_13395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => array_obj_ref_2679_final_reg_req_0); -- 
    base_resize_ack_13386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2679_base_resize_ack_0, ack => cp_elements(59)); -- 
    sum_rename_req_13390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => array_obj_ref_2679_root_address_inst_req_0); -- 
    sum_rename_ack_13391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2679_root_address_inst_ack_0, ack => cp_elements(60)); -- 
    final_reg_ack_13396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2679_final_reg_ack_0, ack => cp_elements(61)); -- 
    base_resize_req_13407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => array_obj_ref_2686_base_resize_req_0); -- 
    cp_elements(62) <= cp_elements(39);
    cpelement_group_63 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(62) & cp_elements(65));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(63),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_13417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => array_obj_ref_2686_final_reg_req_0); -- 
    base_resize_ack_13408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2686_base_resize_ack_0, ack => cp_elements(64)); -- 
    sum_rename_req_13412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => array_obj_ref_2686_root_address_inst_req_0); -- 
    sum_rename_ack_13413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2686_root_address_inst_ack_0, ack => cp_elements(65)); -- 
    final_reg_ack_13418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2686_final_reg_ack_0, ack => cp_elements(66)); -- 
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(68));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13427_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => type_cast_2690_inst_req_0); -- 
    cp_elements(68) <= cp_elements(39);
    ack_13428_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_0, ack => cp_elements(69)); -- 
    pipe_wreq_13439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => simple_obj_ref_2692_inst_req_0); -- 
    pipe_wack_13440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2692_inst_ack_0, ack => cp_elements(70)); -- 
    cp_elements(71) <= cp_elements(70);
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(73) & cp_elements(77));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_2699_load_0_req_0); -- 
    cp_elements(73) <= cp_elements(71);
    cp_elements(74) <= cp_elements(73);
    base_resize_req_13456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_2699_base_resize_req_0); -- 
    base_resize_ack_13457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2699_base_resize_ack_0, ack => cp_elements(75)); -- 
    sum_rename_req_13461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => ptr_deref_2699_root_address_inst_req_0); -- 
    sum_rename_ack_13462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2699_root_address_inst_ack_0, ack => cp_elements(76)); -- 
    root_rename_req_13466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2699_addr_0_req_0); -- 
    root_rename_ack_13467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2699_addr_0_ack_0, ack => cp_elements(77)); -- 
    cp_elements(78) <= ptr_deref_2699_load_0_ack_0;
    cp_elements(79) <= cp_elements(78);
    cr_13488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2699_load_0_req_1); -- 
    ca_13489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2699_load_0_ack_1, ack => cp_elements(80)); -- 
    merge_req_13490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2699_gather_scatter_req_0); -- 
    merge_ack_13491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2699_gather_scatter_ack_0, ack => cp_elements(81)); -- 
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(83));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => binary_2705_inst_req_0); -- 
    cp_elements(83) <= cp_elements(71);
    ra_13501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2705_inst_ack_0, ack => cp_elements(84)); -- 
    cr_13502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => binary_2705_inst_req_1); -- 
    ca_13503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2705_inst_ack_1, ack => cp_elements(85)); -- 
    cpelement_group_86 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(85) & cp_elements(87) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(86),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_13532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2708_gather_scatter_req_0); -- 
    cp_elements(87) <= cp_elements(71);
    cp_elements(88) <= cp_elements(87);
    base_resize_req_13517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2708_base_resize_req_0); -- 
    base_resize_ack_13518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2708_base_resize_ack_0, ack => cp_elements(89)); -- 
    sum_rename_req_13522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2708_root_address_inst_req_0); -- 
    sum_rename_ack_13523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2708_root_address_inst_ack_0, ack => cp_elements(90)); -- 
    root_rename_req_13527_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => ptr_deref_2708_addr_0_req_0); -- 
    root_rename_ack_13528_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2708_addr_0_ack_0, ack => cp_elements(91)); -- 
    split_ack_13533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2708_gather_scatter_ack_0, ack => cp_elements(92)); -- 
    rr_13540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2708_store_0_req_0); -- 
    ra_13541_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2708_store_0_ack_0, ack => cp_elements(93)); -- 
    cr_13551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_2708_store_0_req_1); -- 
    ca_13552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2708_store_0_ack_1, ack => cp_elements(94)); -- 
    cp_elements(95) <= OrReduce(cp_elements(12) & cp_elements(94));
    cp_elements(96) <= cp_elements(95);
    cp_elements(97) <= false;
    cp_elements(98) <= cp_elements(97);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2671_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2671_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2671_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2671_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2679_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2679_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2686_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2686_root_address : std_logic_vector(15 downto 0);
    signal iNsTr_14_2700 : std_logic_vector(31 downto 0);
    signal iNsTr_15_2706 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2649 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2657 : std_logic_vector(0 downto 0);
    signal iNsTr_5_2668 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2673 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2680 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2687 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2691 : std_logic_vector(31 downto 0);
    signal i_2638 : std_logic_vector(31 downto 0);
    signal ptr_deref_2640_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2640_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2640_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2640_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2640_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2640_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2648_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2648_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2648_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2648_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2648_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2667_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2667_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2667_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2667_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2667_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2699_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2699_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2699_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2699_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2699_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2708_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2708_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2708_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2708_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2708_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2708_word_offset_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_2670_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2670_scaled : std_logic_vector(15 downto 0);
    signal type_cast_2642_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2652_wire : std_logic_vector(31 downto 0);
    signal type_cast_2655_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2704_wire_constant : std_logic_vector(31 downto 0);
    signal xxfree_queue_initxxbodyxxi_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_2671_offset_scale_factor_0 <= "0000100000000000";
    array_obj_ref_2671_resized_base_address <= "0000000000000000";
    i_2638 <= "00000000000000000000000000000000";
    ptr_deref_2640_word_offset_0 <= "0";
    ptr_deref_2648_word_offset_0 <= "0";
    ptr_deref_2667_word_offset_0 <= "0";
    ptr_deref_2699_word_offset_0 <= "0";
    ptr_deref_2708_word_offset_0 <= "0";
    type_cast_2642_wire_constant <= "00000000000000000000000000000000";
    type_cast_2655_wire_constant <= "00000000000000000000000000010000";
    type_cast_2704_wire_constant <= "00000000000000000000000000000001";
    xxfree_queue_initxxbodyxxi_alloc_base_address <= "0";
    addr_of_2672_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2671_root_address, dout => iNsTr_6_2673, req => addr_of_2672_final_reg_req_0, ack => addr_of_2672_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2671_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_5_2668, dout => simple_obj_ref_2670_resized, req => array_obj_ref_2671_index_0_resize_req_0, ack => array_obj_ref_2671_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2671_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_2670_scaled, dout => array_obj_ref_2671_final_offset, req => array_obj_ref_2671_offset_inst_req_0, ack => array_obj_ref_2671_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2679_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_6_2673, dout => array_obj_ref_2679_resized_base_address, req => array_obj_ref_2679_base_resize_req_0, ack => array_obj_ref_2679_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2679_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2679_root_address, dout => iNsTr_7_2680, req => array_obj_ref_2679_final_reg_req_0, ack => array_obj_ref_2679_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2686_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_7_2680, dout => array_obj_ref_2686_resized_base_address, req => array_obj_ref_2686_base_resize_req_0, ack => array_obj_ref_2686_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2686_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2686_root_address, dout => iNsTr_8_2687, req => array_obj_ref_2686_final_reg_req_0, ack => array_obj_ref_2686_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2640_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_2638, dout => ptr_deref_2640_resized_base_address, req => ptr_deref_2640_base_resize_req_0, ack => ptr_deref_2640_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2648_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_2638, dout => ptr_deref_2648_resized_base_address, req => ptr_deref_2648_base_resize_req_0, ack => ptr_deref_2648_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2667_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_2638, dout => ptr_deref_2667_resized_base_address, req => ptr_deref_2667_base_resize_req_0, ack => ptr_deref_2667_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2699_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_2638, dout => ptr_deref_2699_resized_base_address, req => ptr_deref_2699_base_resize_req_0, ack => ptr_deref_2699_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2708_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_2638, dout => ptr_deref_2708_resized_base_address, req => ptr_deref_2708_base_resize_req_0, ack => ptr_deref_2708_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2652_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_2_2649, dout => type_cast_2652_wire, req => type_cast_2652_inst_req_0, ack => type_cast_2652_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2690_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_8_2687, dout => iNsTr_9_2691, req => type_cast_2690_inst_req_0, ack => type_cast_2690_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2671_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_2671_root_address_inst_ack_0 <= array_obj_ref_2671_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2671_final_offset;
      array_obj_ref_2671_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_2679_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_2679_root_address_inst_ack_0 <= array_obj_ref_2679_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2679_resized_base_address;
      array_obj_ref_2679_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_2686_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_2686_root_address_inst_ack_0 <= array_obj_ref_2686_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2686_resized_base_address;
      array_obj_ref_2686_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2640_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2640_addr_0_ack_0 <= ptr_deref_2640_addr_0_req_0;
      aggregated_sig <= ptr_deref_2640_root_address;
      ptr_deref_2640_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2640_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2640_gather_scatter_ack_0 <= ptr_deref_2640_gather_scatter_req_0;
      aggregated_sig <= type_cast_2642_wire_constant;
      ptr_deref_2640_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2640_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2640_root_address_inst_ack_0 <= ptr_deref_2640_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2640_resized_base_address;
      ptr_deref_2640_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2648_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2648_addr_0_ack_0 <= ptr_deref_2648_addr_0_req_0;
      aggregated_sig <= ptr_deref_2648_root_address;
      ptr_deref_2648_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2648_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2648_gather_scatter_ack_0 <= ptr_deref_2648_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2648_data_0;
      iNsTr_2_2649 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2648_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2648_root_address_inst_ack_0 <= ptr_deref_2648_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2648_resized_base_address;
      ptr_deref_2648_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2667_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2667_addr_0_ack_0 <= ptr_deref_2667_addr_0_req_0;
      aggregated_sig <= ptr_deref_2667_root_address;
      ptr_deref_2667_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2667_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2667_gather_scatter_ack_0 <= ptr_deref_2667_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2667_data_0;
      iNsTr_5_2668 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2667_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2667_root_address_inst_ack_0 <= ptr_deref_2667_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2667_resized_base_address;
      ptr_deref_2667_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2699_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2699_addr_0_ack_0 <= ptr_deref_2699_addr_0_req_0;
      aggregated_sig <= ptr_deref_2699_root_address;
      ptr_deref_2699_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2699_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2699_gather_scatter_ack_0 <= ptr_deref_2699_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2699_data_0;
      iNsTr_14_2700 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2699_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2699_root_address_inst_ack_0 <= ptr_deref_2699_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2699_resized_base_address;
      ptr_deref_2699_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2708_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2708_addr_0_ack_0 <= ptr_deref_2708_addr_0_req_0;
      aggregated_sig <= ptr_deref_2708_root_address;
      ptr_deref_2708_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_2708_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2708_gather_scatter_ack_0 <= ptr_deref_2708_gather_scatter_req_0;
      aggregated_sig <= iNsTr_15_2706;
      ptr_deref_2708_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2708_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_2708_root_address_inst_ack_0 <= ptr_deref_2708_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2708_resized_base_address;
      ptr_deref_2708_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    if_stmt_2658_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_2657;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2658_branch_req_0,
          ack0 => if_stmt_2658_branch_ack_0,
          ack1 => if_stmt_2658_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_2671_index_0_scale 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2670_resized;
      simple_obj_ref_2670_scaled <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000100000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2671_index_0_scale_req_0,
          ackL => array_obj_ref_2671_index_0_scale_ack_0,
          reqR => array_obj_ref_2671_index_0_scale_req_1,
          ackR => array_obj_ref_2671_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_2656_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2652_wire;
      iNsTr_3_2657 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2656_inst_req_0,
          ackL => binary_2656_inst_ack_0,
          reqR => binary_2656_inst_req_1,
          ackR => binary_2656_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2705_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_14_2700;
      iNsTr_15_2706 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2705_inst_req_0,
          ackL => binary_2705_inst_ack_0,
          reqR => binary_2705_inst_req_1,
          ackR => binary_2705_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : ptr_deref_2699_load_0 ptr_deref_2648_load_0 ptr_deref_2667_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2699_load_0_req_0,
        ptr_deref_2699_load_0_ack_0,
        ptr_deref_2699_load_0_req_1,
        ptr_deref_2699_load_0_ack_1,
        "ptr_deref_2699_load_0",
        "memory_space_6" ,
        ptr_deref_2699_data_0,
        ptr_deref_2699_word_address_0,
        "ptr_deref_2699_data_0",
        "ptr_deref_2699_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2648_load_0_req_0,
        ptr_deref_2648_load_0_ack_0,
        ptr_deref_2648_load_0_req_1,
        ptr_deref_2648_load_0_ack_1,
        "ptr_deref_2648_load_0",
        "memory_space_6" ,
        ptr_deref_2648_data_0,
        ptr_deref_2648_word_address_0,
        "ptr_deref_2648_data_0",
        "ptr_deref_2648_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2667_load_0_req_0,
        ptr_deref_2667_load_0_ack_0,
        ptr_deref_2667_load_0_req_1,
        ptr_deref_2667_load_0_ack_1,
        "ptr_deref_2667_load_0",
        "memory_space_6" ,
        ptr_deref_2667_data_0,
        ptr_deref_2667_word_address_0,
        "ptr_deref_2667_data_0",
        "ptr_deref_2667_word_address_0" -- 
      );
      reqL(2) <= ptr_deref_2699_load_0_req_0;
      reqL(1) <= ptr_deref_2648_load_0_req_0;
      reqL(0) <= ptr_deref_2667_load_0_req_0;
      ptr_deref_2699_load_0_ack_0 <= ackL(2);
      ptr_deref_2648_load_0_ack_0 <= ackL(1);
      ptr_deref_2667_load_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_2699_load_0_req_1;
      reqR(1) <= ptr_deref_2648_load_0_req_1;
      reqR(0) <= ptr_deref_2667_load_0_req_1;
      ptr_deref_2699_load_0_ack_1 <= ackR(2);
      ptr_deref_2648_load_0_ack_1 <= ackR(1);
      ptr_deref_2667_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2699_word_address_0 & ptr_deref_2648_word_address_0 & ptr_deref_2667_word_address_0;
      ptr_deref_2699_data_0 <= data_out(95 downto 64);
      ptr_deref_2648_data_0 <= data_out(63 downto 32);
      ptr_deref_2667_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2708_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_6 address ptr_deref_2708_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2708_word_address_0) &  " data ptr_deref_2708_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2708_data_0) severity note; --
        end if;
        if ptr_deref_2640_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_6 address ptr_deref_2640_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2640_word_address_0) &  " data ptr_deref_2640_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2640_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2708_store_0 ptr_deref_2640_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2708_store_0_req_0;
      reqL(0) <= ptr_deref_2640_store_0_req_0;
      ptr_deref_2708_store_0_ack_0 <= ackL(1);
      ptr_deref_2640_store_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2708_store_0_req_1;
      reqR(0) <= ptr_deref_2640_store_0_req_1;
      ptr_deref_2708_store_0_ack_1 <= ackR(1);
      ptr_deref_2640_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2708_word_address_0 & ptr_deref_2640_word_address_0;
      data_in <= ptr_deref_2708_data_0 & ptr_deref_2640_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(31 downto 0),
          mtag => memory_space_6_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2692_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire iNsTr_9_2691 value="  &  convert_slv_to_hex_string(iNsTr_9_2691) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2692_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2692_inst_req_0;
      simple_obj_ref_2692_inst_ack_0 <= ack(0);
      data_in <= iNsTr_9_2691;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity global_storage_initializer_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    click_bc_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity global_storage_initializer_x;
architecture Default of global_storage_initializer_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal global_storage_initializer_x_xCP_13600_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_2719_call_req_0 : boolean;
  signal call_stmt_2719_call_ack_0 : boolean;
  signal call_stmt_2719_call_req_1 : boolean;
  signal call_stmt_2719_call_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  global_storage_initializer_x_xCP_13600: Block -- control-path 
    signal cp_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    crr_13614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => call_stmt_2719_call_req_0); -- 
    cra_13615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2719_call_ack_0, ack => cp_elements(1)); -- 
    ccr_13619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2719_call_req_1); -- 
    cca_13620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2719_call_ack_1, ack => cp_elements(2)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_2719_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_2719_call_req_0;
      call_stmt_2719_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_2719_call_req_1;
      call_stmt_2719_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => click_bc_storage_initializer_x_call_reqs(0),
          ackR => click_bc_storage_initializer_x_call_acks(0),
          tagR => click_bc_storage_initializer_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => click_bc_storage_initializer_x_return_acks(0), -- cross-over
          ackL => click_bc_storage_initializer_x_return_reqs(0), -- cross-over
          tagL => click_bc_storage_initializer_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity receive_packet_pipeline is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    receive_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
    swapped_in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    swapped_in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    swapped_in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    receive_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
    swapped_in_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    swapped_in_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    swapped_in_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    receive_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_packet_get_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_get_call_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_get_call_tag  :  out  std_logic_vector(0 downto 0);
    ahir_packet_get_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_get_return_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_get_return_data : in   std_logic_vector(31 downto 0);
    ahir_packet_get_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity receive_packet_pipeline;
architecture Default of receive_packet_pipeline is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal receive_packet_pipeline_CP_13792_start: Boolean;
  -- links between control-path and data-path
  signal binary_2744_inst_req_0 : boolean;
  signal binary_2751_inst_req_1 : boolean;
  signal binary_2751_inst_ack_0 : boolean;
  signal binary_2773_inst_ack_1 : boolean;
  signal binary_2772_inst_req_0 : boolean;
  signal binary_2753_inst_req_0 : boolean;
  signal simple_obj_ref_2807_inst_req_0 : boolean;
  signal binary_2773_inst_req_0 : boolean;
  signal type_cast_2762_inst_ack_0 : boolean;
  signal binary_2772_inst_ack_0 : boolean;
  signal type_cast_2752_inst_ack_0 : boolean;
  signal array_obj_ref_2792_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_2824_inst_ack_0 : boolean;
  signal binary_2763_inst_req_0 : boolean;
  signal binary_2753_inst_req_1 : boolean;
  signal simple_obj_ref_2798_inst_req_0 : boolean;
  signal binary_2753_inst_ack_0 : boolean;
  signal type_cast_2809_inst_req_0 : boolean;
  signal binary_2751_inst_ack_1 : boolean;
  signal binary_2751_inst_req_0 : boolean;
  signal binary_2754_inst_ack_1 : boolean;
  signal binary_2773_inst_req_1 : boolean;
  signal binary_2744_inst_req_1 : boolean;
  signal array_obj_ref_2792_root_address_inst_ack_1 : boolean;
  signal type_cast_2739_inst_ack_0 : boolean;
  signal simple_obj_ref_2798_inst_ack_0 : boolean;
  signal type_cast_2752_inst_req_0 : boolean;
  signal binary_2774_inst_req_1 : boolean;
  signal binary_2744_inst_ack_1 : boolean;
  signal simple_obj_ref_2737_inst_req_0 : boolean;
  signal simple_obj_ref_2737_inst_ack_0 : boolean;
  signal binary_2754_inst_ack_0 : boolean;
  signal simple_obj_ref_2833_inst_ack_0 : boolean;
  signal simple_obj_ref_2804_inst_ack_0 : boolean;
  signal binary_2774_inst_req_0 : boolean;
  signal binary_2754_inst_req_0 : boolean;
  signal binary_2773_inst_ack_0 : boolean;
  signal simple_obj_ref_2735_inst_ack_0 : boolean;
  signal binary_2774_inst_ack_0 : boolean;
  signal binary_2754_inst_req_1 : boolean;
  signal binary_2753_inst_ack_1 : boolean;
  signal simple_obj_ref_2824_inst_req_0 : boolean;
  signal type_cast_2739_inst_req_0 : boolean;
  signal binary_2744_inst_ack_0 : boolean;
  signal array_obj_ref_2792_root_address_inst_req_1 : boolean;
  signal simple_obj_ref_2836_inst_ack_0 : boolean;
  signal type_cast_2788_inst_req_0 : boolean;
  signal simple_obj_ref_2804_inst_req_0 : boolean;
  signal binary_2772_inst_req_1 : boolean;
  signal simple_obj_ref_2735_inst_req_0 : boolean;
  signal binary_2772_inst_ack_1 : boolean;
  signal array_obj_ref_2792_root_address_inst_req_0 : boolean;
  signal type_cast_2788_inst_ack_0 : boolean;
  signal simple_obj_ref_2807_inst_ack_0 : boolean;
  signal binary_2774_inst_ack_1 : boolean;
  signal simple_obj_ref_2821_inst_ack_0 : boolean;
  signal simple_obj_ref_2827_inst_ack_0 : boolean;
  signal type_cast_2771_inst_ack_0 : boolean;
  signal type_cast_2771_inst_req_0 : boolean;
  signal type_cast_2784_inst_ack_0 : boolean;
  signal binary_2770_inst_ack_1 : boolean;
  signal binary_2770_inst_req_1 : boolean;
  signal type_cast_2784_inst_req_0 : boolean;
  signal binary_2770_inst_ack_0 : boolean;
  signal binary_2770_inst_req_0 : boolean;
  signal type_cast_2758_inst_ack_0 : boolean;
  signal binary_2761_inst_ack_1 : boolean;
  signal simple_obj_ref_2801_inst_ack_0 : boolean;
  signal type_cast_2758_inst_req_0 : boolean;
  signal type_cast_2762_inst_req_0 : boolean;
  signal type_cast_2767_inst_ack_0 : boolean;
  signal binary_2757_inst_ack_1 : boolean;
  signal type_cast_2748_inst_ack_0 : boolean;
  signal type_cast_2748_inst_req_0 : boolean;
  signal binary_2757_inst_req_1 : boolean;
  signal type_cast_2767_inst_req_0 : boolean;
  signal simple_obj_ref_2801_inst_req_0 : boolean;
  signal binary_2761_inst_req_0 : boolean;
  signal array_obj_ref_2792_base_resize_req_0 : boolean;
  signal array_obj_ref_2792_base_resize_ack_0 : boolean;
  signal simple_obj_ref_2833_inst_req_0 : boolean;
  signal type_cast_2809_inst_ack_0 : boolean;
  signal binary_2761_inst_ack_0 : boolean;
  signal binary_2761_inst_req_1 : boolean;
  signal binary_2742_inst_req_0 : boolean;
  signal simple_obj_ref_2827_inst_req_0 : boolean;
  signal binary_2742_inst_ack_0 : boolean;
  signal binary_2742_inst_req_1 : boolean;
  signal binary_2742_inst_ack_1 : boolean;
  signal call_stmt_2781_call_req_0 : boolean;
  signal call_stmt_2781_call_ack_0 : boolean;
  signal type_cast_2743_inst_req_0 : boolean;
  signal call_stmt_2781_call_req_1 : boolean;
  signal call_stmt_2781_call_ack_1 : boolean;
  signal binary_2757_inst_req_0 : boolean;
  signal binary_2757_inst_ack_0 : boolean;
  signal type_cast_2743_inst_ack_0 : boolean;
  signal binary_2747_inst_ack_1 : boolean;
  signal binary_2766_inst_ack_1 : boolean;
  signal binary_2747_inst_req_1 : boolean;
  signal binary_2766_inst_req_1 : boolean;
  signal binary_2766_inst_ack_0 : boolean;
  signal binary_2766_inst_req_0 : boolean;
  signal binary_2747_inst_ack_0 : boolean;
  signal binary_2747_inst_req_0 : boolean;
  signal array_obj_ref_2792_final_reg_ack_0 : boolean;
  signal simple_obj_ref_2836_inst_req_0 : boolean;
  signal array_obj_ref_2792_final_reg_req_0 : boolean;
  signal simple_obj_ref_2818_inst_ack_0 : boolean;
  signal simple_obj_ref_2818_inst_req_0 : boolean;
  signal binary_2763_inst_ack_1 : boolean;
  signal simple_obj_ref_2794_inst_ack_0 : boolean;
  signal simple_obj_ref_2821_inst_req_0 : boolean;
  signal binary_2763_inst_req_1 : boolean;
  signal simple_obj_ref_2794_inst_req_0 : boolean;
  signal binary_2763_inst_ack_0 : boolean;
  signal binary_2842_inst_req_0 : boolean;
  signal binary_2842_inst_ack_0 : boolean;
  signal binary_2842_inst_req_1 : boolean;
  signal binary_2842_inst_ack_1 : boolean;
  signal if_stmt_2839_branch_req_0 : boolean;
  signal if_stmt_2839_branch_ack_1 : boolean;
  signal if_stmt_2839_branch_ack_0 : boolean;
  signal simple_obj_ref_2846_inst_req_0 : boolean;
  signal simple_obj_ref_2846_inst_ack_0 : boolean;
  signal simple_obj_ref_2849_inst_req_0 : boolean;
  signal simple_obj_ref_2849_inst_ack_0 : boolean;
  signal simple_obj_ref_2852_inst_req_0 : boolean;
  signal simple_obj_ref_2852_inst_ack_0 : boolean;
  signal simple_obj_ref_2865_inst_req_0 : boolean;
  signal simple_obj_ref_2865_inst_ack_0 : boolean;
  signal simple_obj_ref_2868_inst_req_0 : boolean;
  signal simple_obj_ref_2868_inst_ack_0 : boolean;
  signal binary_2873_inst_req_0 : boolean;
  signal binary_2873_inst_ack_0 : boolean;
  signal binary_2873_inst_req_1 : boolean;
  signal binary_2873_inst_ack_1 : boolean;
  signal simple_obj_ref_2877_inst_req_0 : boolean;
  signal simple_obj_ref_2877_inst_ack_0 : boolean;
  signal array_obj_ref_2882_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2882_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2882_index_0_scale_req_0 : boolean;
  signal array_obj_ref_2882_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_2882_index_0_scale_req_1 : boolean;
  signal array_obj_ref_2882_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_2882_offset_inst_req_0 : boolean;
  signal array_obj_ref_2882_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2882_base_resize_req_0 : boolean;
  signal array_obj_ref_2882_base_resize_ack_0 : boolean;
  signal array_obj_ref_2882_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2882_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2882_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2882_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2882_final_reg_req_0 : boolean;
  signal array_obj_ref_2882_final_reg_ack_0 : boolean;
  signal simple_obj_ref_2880_inst_req_0 : boolean;
  signal simple_obj_ref_2880_inst_ack_0 : boolean;
  signal binary_2887_inst_req_0 : boolean;
  signal binary_2887_inst_ack_0 : boolean;
  signal binary_2887_inst_req_1 : boolean;
  signal binary_2887_inst_ack_1 : boolean;
  signal ternary_2890_inst_req_0 : boolean;
  signal ternary_2890_inst_ack_0 : boolean;
  signal simple_obj_ref_2884_inst_req_0 : boolean;
  signal simple_obj_ref_2884_inst_ack_0 : boolean;
  signal binary_2896_inst_req_0 : boolean;
  signal binary_2896_inst_ack_0 : boolean;
  signal binary_2896_inst_req_1 : boolean;
  signal binary_2896_inst_ack_1 : boolean;
  signal if_stmt_2893_branch_req_0 : boolean;
  signal if_stmt_2893_branch_ack_1 : boolean;
  signal if_stmt_2893_branch_ack_0 : boolean;
  signal phi_stmt_2857_req_0 : boolean;
  signal phi_stmt_2857_req_1 : boolean;
  signal phi_stmt_2857_ack_0 : boolean;
  signal simple_obj_ref_2905_inst_req_0 : boolean;
  signal simple_obj_ref_2905_inst_ack_0 : boolean;
  signal simple_obj_ref_2903_inst_req_0 : boolean;
  signal simple_obj_ref_2903_inst_ack_0 : boolean;
  signal ptr_deref_2904_base_resize_req_0 : boolean;
  signal ptr_deref_2904_base_resize_ack_0 : boolean;
  signal ptr_deref_2904_root_address_inst_req_0 : boolean;
  signal ptr_deref_2904_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2904_addr_0_req_0 : boolean;
  signal ptr_deref_2904_addr_0_ack_0 : boolean;
  signal ptr_deref_2904_addr_0_req_1 : boolean;
  signal ptr_deref_2904_addr_0_ack_1 : boolean;
  signal ptr_deref_2904_addr_1_req_0 : boolean;
  signal ptr_deref_2904_addr_1_ack_0 : boolean;
  signal ptr_deref_2904_addr_1_req_1 : boolean;
  signal ptr_deref_2904_addr_1_ack_1 : boolean;
  signal ptr_deref_2904_addr_2_req_0 : boolean;
  signal ptr_deref_2904_addr_2_ack_0 : boolean;
  signal ptr_deref_2904_addr_2_req_1 : boolean;
  signal ptr_deref_2904_addr_2_ack_1 : boolean;
  signal ptr_deref_2904_addr_3_req_0 : boolean;
  signal ptr_deref_2904_addr_3_ack_0 : boolean;
  signal ptr_deref_2904_addr_3_req_1 : boolean;
  signal ptr_deref_2904_addr_3_ack_1 : boolean;
  signal ptr_deref_2904_addr_4_req_0 : boolean;
  signal ptr_deref_2904_addr_4_ack_0 : boolean;
  signal ptr_deref_2904_addr_4_req_1 : boolean;
  signal ptr_deref_2904_addr_4_ack_1 : boolean;
  signal ptr_deref_2904_addr_5_req_0 : boolean;
  signal ptr_deref_2904_addr_5_ack_0 : boolean;
  signal ptr_deref_2904_addr_5_req_1 : boolean;
  signal ptr_deref_2904_addr_5_ack_1 : boolean;
  signal ptr_deref_2904_addr_6_req_0 : boolean;
  signal ptr_deref_2904_addr_6_ack_0 : boolean;
  signal ptr_deref_2904_addr_6_req_1 : boolean;
  signal ptr_deref_2904_addr_6_ack_1 : boolean;
  signal ptr_deref_2904_addr_7_req_0 : boolean;
  signal ptr_deref_2904_addr_7_ack_0 : boolean;
  signal ptr_deref_2904_addr_7_req_1 : boolean;
  signal ptr_deref_2904_addr_7_ack_1 : boolean;
  signal ptr_deref_2904_gather_scatter_req_0 : boolean;
  signal ptr_deref_2904_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2904_store_0_req_0 : boolean;
  signal ptr_deref_2904_store_0_ack_0 : boolean;
  signal ptr_deref_2904_store_1_req_0 : boolean;
  signal ptr_deref_2904_store_1_ack_0 : boolean;
  signal ptr_deref_2904_store_2_req_0 : boolean;
  signal ptr_deref_2904_store_2_ack_0 : boolean;
  signal ptr_deref_2904_store_3_req_0 : boolean;
  signal ptr_deref_2904_store_3_ack_0 : boolean;
  signal ptr_deref_2904_store_4_req_0 : boolean;
  signal ptr_deref_2904_store_4_ack_0 : boolean;
  signal ptr_deref_2904_store_5_req_0 : boolean;
  signal ptr_deref_2904_store_5_ack_0 : boolean;
  signal ptr_deref_2904_store_6_req_0 : boolean;
  signal ptr_deref_2904_store_6_ack_0 : boolean;
  signal ptr_deref_2904_store_7_req_0 : boolean;
  signal ptr_deref_2904_store_7_ack_0 : boolean;
  signal ptr_deref_2904_store_0_req_1 : boolean;
  signal ptr_deref_2904_store_0_ack_1 : boolean;
  signal ptr_deref_2904_store_1_req_1 : boolean;
  signal ptr_deref_2904_store_1_ack_1 : boolean;
  signal ptr_deref_2904_store_2_req_1 : boolean;
  signal ptr_deref_2904_store_2_ack_1 : boolean;
  signal ptr_deref_2904_store_3_req_1 : boolean;
  signal ptr_deref_2904_store_3_ack_1 : boolean;
  signal ptr_deref_2904_store_4_req_1 : boolean;
  signal ptr_deref_2904_store_4_ack_1 : boolean;
  signal ptr_deref_2904_store_5_req_1 : boolean;
  signal ptr_deref_2904_store_5_ack_1 : boolean;
  signal ptr_deref_2904_store_6_req_1 : boolean;
  signal ptr_deref_2904_store_6_ack_1 : boolean;
  signal ptr_deref_2904_store_7_req_1 : boolean;
  signal ptr_deref_2904_store_7_ack_1 : boolean;
  signal simple_obj_ref_2908_inst_req_0 : boolean;
  signal simple_obj_ref_2908_inst_ack_0 : boolean;
  signal binary_2910_inst_req_0 : boolean;
  signal binary_2910_inst_ack_0 : boolean;
  signal binary_2910_inst_req_1 : boolean;
  signal binary_2910_inst_ack_1 : boolean;
  signal if_stmt_2907_branch_req_0 : boolean;
  signal if_stmt_2907_branch_ack_1 : boolean;
  signal if_stmt_2907_branch_ack_0 : boolean;
  signal simple_obj_ref_2912_inst_req_0 : boolean;
  signal simple_obj_ref_2912_inst_ack_0 : boolean;
  signal type_cast_2913_inst_req_0 : boolean;
  signal type_cast_2913_inst_ack_0 : boolean;
  signal simple_obj_ref_2911_inst_req_0 : boolean;
  signal simple_obj_ref_2911_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  receive_packet_pipeline_CP_13792: Block -- control-path 
    signal cp_elements: BooleanArray(361 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(361);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(361), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    cp_elements(2) <= false; 
    cp_elements(3) <= OrReduce(cp_elements(97) & cp_elements(100));
    req_13819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2735_inst_req_0); -- 
    ack_13820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2735_inst_ack_0, ack => cp_elements(4)); -- 
    cp_elements(5) <= cp_elements(4);
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(7) & cp_elements(47) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => binary_2774_inst_req_0); -- 
    cp_elements(7) <= cp_elements(5);
    cpelement_group_8 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(9) & cp_elements(25) & cp_elements(45));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(8),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => binary_2754_inst_req_0); -- 
    cp_elements(9) <= cp_elements(5);
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(15) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => binary_2744_inst_req_0); -- 
    cp_elements(11) <= cp_elements(5);
    cpelement_group_12 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(13) & cp_elements(14));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(12),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => type_cast_2739_inst_req_0); -- 
    cp_elements(13) <= cp_elements(5);
    cp_elements(14) <= cp_elements(5);
    ack_13839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_0, ack => cp_elements(15)); -- 
    cpelement_group_16 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(17) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(16),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => type_cast_2743_inst_req_0); -- 
    cp_elements(17) <= cp_elements(5);
    cpelement_group_18 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(20));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(18),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13848_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2742_inst_req_0); -- 
    cp_elements(19) <= cp_elements(5);
    cp_elements(20) <= cp_elements(5);
    ra_13849_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2742_inst_ack_0, ack => cp_elements(21)); -- 
    cr_13850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => binary_2742_inst_req_1); -- 
    ca_13851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2742_inst_ack_1, ack => cp_elements(22)); -- 
    ack_13856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2743_inst_ack_0, ack => cp_elements(23)); -- 
    ra_13861_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2744_inst_ack_0, ack => cp_elements(24)); -- 
    cr_13862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => binary_2744_inst_req_1); -- 
    ca_13863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2744_inst_ack_1, ack => cp_elements(25)); -- 
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(35) & cp_elements(43));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => binary_2753_inst_req_0); -- 
    cp_elements(27) <= cp_elements(5);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(29) & cp_elements(34));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => type_cast_2748_inst_req_0); -- 
    cp_elements(29) <= cp_elements(5);
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(31) & cp_elements(32));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => binary_2747_inst_req_0); -- 
    cp_elements(31) <= cp_elements(5);
    cp_elements(32) <= cp_elements(5);
    ra_13875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2747_inst_ack_0, ack => cp_elements(33)); -- 
    cr_13876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => binary_2747_inst_req_1); -- 
    ca_13877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2747_inst_ack_1, ack => cp_elements(34)); -- 
    ack_13882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2748_inst_ack_0, ack => cp_elements(35)); -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(37) & cp_elements(42));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => type_cast_2752_inst_req_0); -- 
    cp_elements(37) <= cp_elements(5);
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(39) & cp_elements(40));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => binary_2751_inst_req_0); -- 
    cp_elements(39) <= cp_elements(5);
    cp_elements(40) <= cp_elements(5);
    ra_13892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2751_inst_ack_0, ack => cp_elements(41)); -- 
    cr_13893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => binary_2751_inst_req_1); -- 
    ca_13894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2751_inst_ack_1, ack => cp_elements(42)); -- 
    ack_13899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2752_inst_ack_0, ack => cp_elements(43)); -- 
    ra_13904_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2753_inst_ack_0, ack => cp_elements(44)); -- 
    cr_13905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => binary_2753_inst_req_1); -- 
    ca_13906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2753_inst_ack_1, ack => cp_elements(45)); -- 
    ra_13911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2754_inst_ack_0, ack => cp_elements(46)); -- 
    cr_13912_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => binary_2754_inst_req_1); -- 
    ca_13913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2754_inst_ack_1, ack => cp_elements(47)); -- 
    cpelement_group_48 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(49) & cp_elements(69) & cp_elements(89));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(48),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => binary_2773_inst_req_0); -- 
    cp_elements(49) <= cp_elements(5);
    cpelement_group_50 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(50),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => binary_2763_inst_req_0); -- 
    cp_elements(51) <= cp_elements(5);
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => type_cast_2758_inst_req_0); -- 
    cp_elements(53) <= cp_elements(5);
    cpelement_group_54 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(55) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(54),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => binary_2757_inst_req_0); -- 
    cp_elements(55) <= cp_elements(5);
    cp_elements(56) <= cp_elements(5);
    ra_13927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2757_inst_ack_0, ack => cp_elements(57)); -- 
    cr_13928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => binary_2757_inst_req_1); -- 
    ca_13929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2757_inst_ack_1, ack => cp_elements(58)); -- 
    ack_13934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => type_cast_2762_inst_req_0); -- 
    cp_elements(61) <= cp_elements(5);
    cpelement_group_62 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(63) & cp_elements(64));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(62),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => binary_2761_inst_req_0); -- 
    cp_elements(63) <= cp_elements(5);
    cp_elements(64) <= cp_elements(5);
    ra_13944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2761_inst_ack_0, ack => cp_elements(65)); -- 
    cr_13945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => binary_2761_inst_req_1); -- 
    ca_13946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2761_inst_ack_1, ack => cp_elements(66)); -- 
    ack_13951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_0, ack => cp_elements(67)); -- 
    ra_13956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2763_inst_ack_0, ack => cp_elements(68)); -- 
    cr_13957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => binary_2763_inst_req_1); -- 
    ca_13958_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2763_inst_ack_1, ack => cp_elements(69)); -- 
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(79) & cp_elements(87));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => binary_2772_inst_req_0); -- 
    cp_elements(71) <= cp_elements(5);
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(73) & cp_elements(78));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => type_cast_2767_inst_req_0); -- 
    cp_elements(73) <= cp_elements(5);
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(76));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13969_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => binary_2766_inst_req_0); -- 
    cp_elements(75) <= cp_elements(5);
    cp_elements(76) <= cp_elements(5);
    ra_13970_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2766_inst_ack_0, ack => cp_elements(77)); -- 
    cr_13971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => binary_2766_inst_req_1); -- 
    ca_13972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2766_inst_ack_1, ack => cp_elements(78)); -- 
    ack_13977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_0, ack => cp_elements(79)); -- 
    cpelement_group_80 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(86));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(80),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => type_cast_2771_inst_req_0); -- 
    cp_elements(81) <= cp_elements(5);
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => binary_2770_inst_req_0); -- 
    cp_elements(83) <= cp_elements(5);
    cp_elements(84) <= cp_elements(5);
    ra_13987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2770_inst_ack_0, ack => cp_elements(85)); -- 
    cr_13988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => binary_2770_inst_req_1); -- 
    ca_13989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2770_inst_ack_1, ack => cp_elements(86)); -- 
    ack_13994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_0, ack => cp_elements(87)); -- 
    ra_13999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2772_inst_ack_0, ack => cp_elements(88)); -- 
    cr_14000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => binary_2772_inst_req_1); -- 
    ca_14001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2772_inst_ack_1, ack => cp_elements(89)); -- 
    ra_14006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2773_inst_ack_0, ack => cp_elements(90)); -- 
    cr_14007_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => binary_2773_inst_req_1); -- 
    ca_14008_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2773_inst_ack_1, ack => cp_elements(91)); -- 
    ra_14013_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2774_inst_ack_0, ack => cp_elements(92)); -- 
    cr_14014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => binary_2774_inst_req_1); -- 
    ca_14015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2774_inst_ack_1, ack => cp_elements(93)); -- 
    pipe_wreq_14020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => simple_obj_ref_2737_inst_req_0); -- 
    pipe_wack_14021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2737_inst_ack_0, ack => cp_elements(94)); -- 
    cp_elements(95) <= cp_elements(1);
    cp_elements(96) <= false;
    cp_elements(97) <= cp_elements(96);
    cp_elements(98) <= cp_elements(1);
    cp_elements(99) <= OrReduce(cp_elements(94) & cp_elements(98));
    cp_elements(100) <= cp_elements(99);
    cp_elements(101) <= cp_elements(0);
    cp_elements(102) <= false; 
    cp_elements(103) <= OrReduce(cp_elements(141) & cp_elements(144));
    crr_14061_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => call_stmt_2781_call_req_0); -- 
    cp_elements(104) <= cp_elements(123);
    pipe_wreq_14128_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => simple_obj_ref_2794_inst_req_0); -- 
    cp_elements(105) <= cp_elements(138);
    cra_14062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2781_call_ack_0, ack => cp_elements(106)); -- 
    ccr_14066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => call_stmt_2781_call_req_1); -- 
    cca_14067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2781_call_ack_1, ack => cp_elements(107)); -- 
    cp_elements(108) <= cp_elements(107);
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(111));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => type_cast_2784_inst_req_0); -- 
    cp_elements(110) <= cp_elements(108);
    cp_elements(111) <= cp_elements(108);
    ack_14082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2784_inst_ack_0, ack => cp_elements(112)); -- 
    base_resize_req_14103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => array_obj_ref_2792_base_resize_req_0); -- 
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(115));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => type_cast_2788_inst_req_0); -- 
    cp_elements(114) <= cp_elements(108);
    cp_elements(115) <= cp_elements(108);
    ack_14092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2788_inst_ack_0, ack => cp_elements(116)); -- 
    cp_elements(117) <= cp_elements(108);
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(117) & cp_elements(121));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_14116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2792_final_reg_req_0); -- 
    base_resize_ack_14104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2792_base_resize_ack_0, ack => cp_elements(119)); -- 
    plus_base_rr_14109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => array_obj_ref_2792_root_address_inst_req_0); -- 
    plus_base_ra_14110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2792_root_address_inst_ack_0, ack => cp_elements(120)); -- 
    plus_base_cr_14111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => array_obj_ref_2792_root_address_inst_req_1); -- 
    plus_base_ca_14112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2792_root_address_inst_ack_1, ack => cp_elements(121)); -- 
    final_reg_ack_14117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2792_final_reg_ack_0, ack => cp_elements(122)); -- 
    cpelement_group_123 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(116) & cp_elements(122));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(123),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_14129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2794_inst_ack_0, ack => cp_elements(124)); -- 
    cp_elements(125) <= cp_elements(124);
    cp_elements(126) <= cp_elements(125);
    pipe_wreq_14143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => simple_obj_ref_2798_inst_req_0); -- 
    pipe_wack_14144_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2798_inst_ack_0, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(125);
    pipe_wreq_14155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => simple_obj_ref_2801_inst_req_0); -- 
    pipe_wack_14156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2801_inst_ack_0, ack => cp_elements(129)); -- 
    cp_elements(130) <= cp_elements(125);
    pipe_wreq_14167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => simple_obj_ref_2804_inst_req_0); -- 
    pipe_wack_14168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2804_inst_ack_0, ack => cp_elements(131)); -- 
    cp_elements(132) <= cp_elements(125);
    cpelement_group_133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(135));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => type_cast_2809_inst_req_0); -- 
    cp_elements(134) <= cp_elements(132);
    cp_elements(135) <= cp_elements(132);
    ack_14181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_0, ack => cp_elements(136)); -- 
    pipe_wreq_14186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => simple_obj_ref_2807_inst_req_0); -- 
    pipe_wack_14187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2807_inst_ack_0, ack => cp_elements(137)); -- 
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(129) & cp_elements(131) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(139) <= cp_elements(101);
    cp_elements(140) <= false;
    cp_elements(141) <= cp_elements(140);
    cp_elements(142) <= cp_elements(101);
    cp_elements(143) <= OrReduce(cp_elements(105) & cp_elements(142));
    cp_elements(144) <= cp_elements(143);
    cp_elements(145) <= cp_elements(0);
    cp_elements(146) <= false; 
    cp_elements(147) <= OrReduce(cp_elements(246) & cp_elements(249));
    cp_elements(148) <= cp_elements(166);
    cp_elements(149) <= OrReduce(cp_elements(252) & cp_elements(255));
    cp_elements(150) <= cp_elements(172);
    cp_elements(151) <= OrReduce(cp_elements(175) & cp_elements(183));
    cp_elements(152) <= cp_elements(191);
    cp_elements(153) <= OrReduce(cp_elements(258) & cp_elements(262));
    cp_elements(154) <= cp_elements(203);
    cp_elements(155) <= cp_elements(232);
    cp_elements(156) <= OrReduce(cp_elements(235) & cp_elements(243));
    cp_elements(157) <= cp_elements(147);
    cp_elements(158) <= cp_elements(157);
    req_14241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => simple_obj_ref_2818_inst_req_0); -- 
    ack_14242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2818_inst_ack_0, ack => cp_elements(159)); -- 
    cp_elements(160) <= cp_elements(157);
    req_14252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => simple_obj_ref_2821_inst_req_0); -- 
    ack_14253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2821_inst_ack_0, ack => cp_elements(161)); -- 
    cp_elements(162) <= cp_elements(157);
    req_14263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => simple_obj_ref_2824_inst_req_0); -- 
    ack_14264_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2824_inst_ack_0, ack => cp_elements(163)); -- 
    cp_elements(164) <= cp_elements(157);
    req_14274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => simple_obj_ref_2827_inst_req_0); -- 
    ack_14275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2827_inst_ack_0, ack => cp_elements(165)); -- 
    cpelement_group_166 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(159) & cp_elements(161) & cp_elements(163) & cp_elements(165));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(167) <= cp_elements(149);
    cp_elements(168) <= cp_elements(167);
    req_14288_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => simple_obj_ref_2833_inst_req_0); -- 
    ack_14289_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2833_inst_ack_0, ack => cp_elements(169)); -- 
    cp_elements(170) <= cp_elements(167);
    req_14299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => simple_obj_ref_2836_inst_req_0); -- 
    ack_14300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2836_inst_ack_0, ack => cp_elements(171)); -- 
    cpelement_group_172 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(171));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(172),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(173) <= cp_elements(150);
    cp_elements(174) <= false;
    cp_elements(175) <= cp_elements(174);
    cp_elements(176) <= cp_elements(150);
    rr_14314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2842_inst_req_0); -- 
    ra_14315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2842_inst_ack_0, ack => cp_elements(177)); -- 
    cr_14316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => binary_2842_inst_req_1); -- 
    ca_14317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2842_inst_ack_1, ack => cp_elements(178)); -- 
    branch_req_14318_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => if_stmt_2839_branch_req_0); -- 
    cp_elements(179) <= cp_elements(178);
    cp_elements(180) <= cp_elements(179);
    if_choice_transition_14323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2839_branch_ack_1, ack => cp_elements(181)); -- 
    cp_elements(182) <= cp_elements(179);
    else_choice_transition_14327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2839_branch_ack_0, ack => cp_elements(183)); -- 
    cp_elements(184) <= cp_elements(151);
    cp_elements(185) <= cp_elements(184);
    pipe_wreq_14342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => simple_obj_ref_2846_inst_req_0); -- 
    pipe_wack_14343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2846_inst_ack_0, ack => cp_elements(186)); -- 
    cp_elements(187) <= cp_elements(184);
    pipe_wreq_14353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => simple_obj_ref_2849_inst_req_0); -- 
    pipe_wack_14354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2849_inst_ack_0, ack => cp_elements(188)); -- 
    cp_elements(189) <= cp_elements(184);
    pipe_wreq_14365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => simple_obj_ref_2852_inst_req_0); -- 
    pipe_wack_14366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2852_inst_ack_0, ack => cp_elements(190)); -- 
    cpelement_group_191 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(188) & cp_elements(190));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(191),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(192) <= cp_elements(153);
    cp_elements(193) <= cp_elements(192);
    req_14379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => simple_obj_ref_2865_inst_req_0); -- 
    ack_14380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2865_inst_ack_0, ack => cp_elements(194)); -- 
    cp_elements(195) <= cp_elements(192);
    req_14390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => simple_obj_ref_2868_inst_req_0); -- 
    ack_14391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2868_inst_ack_0, ack => cp_elements(196)); -- 
    cp_elements(197) <= cp_elements(192);
    cpelement_group_198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(199) & cp_elements(200));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => binary_2873_inst_req_0); -- 
    cp_elements(199) <= cp_elements(197);
    cp_elements(200) <= cp_elements(197);
    ra_14404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2873_inst_ack_0, ack => cp_elements(201)); -- 
    cr_14405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => binary_2873_inst_req_1); -- 
    ca_14406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2873_inst_ack_1, ack => cp_elements(202)); -- 
    cpelement_group_203 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(194) & cp_elements(196) & cp_elements(202));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(203),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(204) <= cp_elements(154);
    cp_elements(205) <= cp_elements(204);
    pipe_wreq_14420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => simple_obj_ref_2877_inst_req_0); -- 
    pipe_wack_14421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2877_inst_ack_0, ack => cp_elements(206)); -- 
    cp_elements(207) <= cp_elements(204);
    cp_elements(208) <= cp_elements(207);
    cpelement_group_209 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(208) & cp_elements(219));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(209),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_14470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => array_obj_ref_2882_final_reg_req_0); -- 
    cp_elements(210) <= cp_elements(207);
    base_resize_req_14457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => array_obj_ref_2882_base_resize_req_0); -- 
    cp_elements(211) <= cp_elements(207);
    index_resize_req_14439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => array_obj_ref_2882_index_0_resize_req_0); -- 
    index_resize_ack_14440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_index_0_resize_ack_0, ack => cp_elements(212)); -- 
    scale_rr_14444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => array_obj_ref_2882_index_0_scale_req_0); -- 
    scale_ra_14445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_index_0_scale_ack_0, ack => cp_elements(213)); -- 
    scale_cr_14446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => array_obj_ref_2882_index_0_scale_req_1); -- 
    scale_ca_14447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_index_0_scale_ack_1, ack => cp_elements(214)); -- 
    final_index_req_14451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => array_obj_ref_2882_offset_inst_req_0); -- 
    final_index_ack_14452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_offset_inst_ack_0, ack => cp_elements(215)); -- 
    base_resize_ack_14458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_base_resize_ack_0, ack => cp_elements(216)); -- 
    cpelement_group_217 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(215) & cp_elements(216));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(217),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_14463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => array_obj_ref_2882_root_address_inst_req_0); -- 
    plus_base_ra_14464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_root_address_inst_ack_0, ack => cp_elements(218)); -- 
    plus_base_cr_14465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(218), ack => array_obj_ref_2882_root_address_inst_req_1); -- 
    plus_base_ca_14466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_root_address_inst_ack_1, ack => cp_elements(219)); -- 
    final_reg_ack_14471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2882_final_reg_ack_0, ack => cp_elements(220)); -- 
    pipe_wreq_14476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(220), ack => simple_obj_ref_2880_inst_req_0); -- 
    pipe_wack_14477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2880_inst_ack_0, ack => cp_elements(221)); -- 
    cp_elements(222) <= cp_elements(204);
    cp_elements(223) <= cp_elements(222);
    cpelement_group_224 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(229));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(224),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ternary_2890_inst_req_0); -- 
    cpelement_group_225 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(226) & cp_elements(227));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(225),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14491_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => binary_2887_inst_req_0); -- 
    cp_elements(226) <= cp_elements(222);
    cp_elements(227) <= cp_elements(222);
    ra_14492_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2887_inst_ack_0, ack => cp_elements(228)); -- 
    cr_14493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => binary_2887_inst_req_1); -- 
    ca_14494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2887_inst_ack_1, ack => cp_elements(229)); -- 
    ack_14499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ternary_2890_inst_ack_0, ack => cp_elements(230)); -- 
    pipe_wreq_14504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => simple_obj_ref_2884_inst_req_0); -- 
    pipe_wack_14505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2884_inst_ack_0, ack => cp_elements(231)); -- 
    cpelement_group_232 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(206) & cp_elements(221) & cp_elements(231));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(232),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(233) <= cp_elements(155);
    cp_elements(234) <= false;
    cp_elements(235) <= cp_elements(234);
    cp_elements(236) <= cp_elements(155);
    rr_14519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => binary_2896_inst_req_0); -- 
    ra_14520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2896_inst_ack_0, ack => cp_elements(237)); -- 
    cr_14521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => binary_2896_inst_req_1); -- 
    ca_14522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2896_inst_ack_1, ack => cp_elements(238)); -- 
    branch_req_14523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => if_stmt_2893_branch_req_0); -- 
    cp_elements(239) <= cp_elements(238);
    cp_elements(240) <= cp_elements(239);
    if_choice_transition_14528_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2893_branch_ack_1, ack => cp_elements(241)); -- 
    phi_stmt_2857_req_14587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => phi_stmt_2857_req_1); -- 
    cp_elements(242) <= cp_elements(239);
    else_choice_transition_14532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2893_branch_ack_0, ack => cp_elements(243)); -- 
    cp_elements(244) <= cp_elements(145);
    cp_elements(245) <= false;
    cp_elements(246) <= cp_elements(245);
    cp_elements(247) <= cp_elements(145);
    cp_elements(248) <= OrReduce(cp_elements(156) & cp_elements(247));
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(148);
    cp_elements(251) <= false;
    cp_elements(252) <= cp_elements(251);
    cp_elements(253) <= cp_elements(148);
    cp_elements(254) <= OrReduce(cp_elements(181) & cp_elements(253));
    cp_elements(255) <= cp_elements(254);
    cp_elements(256) <= cp_elements(152);
    cp_elements(257) <= false;
    cp_elements(258) <= cp_elements(257);
    cp_elements(259) <= cp_elements(152);
    phi_stmt_2857_req_14577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => phi_stmt_2857_req_0); -- 
    cp_elements(260) <= OrReduce(cp_elements(241) & cp_elements(259));
    cp_elements(261) <= cp_elements(260);
    phi_stmt_2857_ack_14592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2857_ack_0, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(0);
    cp_elements(264) <= false; 
    cp_elements(265) <= OrReduce(cp_elements(357) & cp_elements(360));
    cp_elements(266) <= OrReduce(cp_elements(338) & cp_elements(347) & cp_elements(354));
    cp_elements(267) <= cp_elements(265);
    cp_elements(268) <= cp_elements(267);
    req_14614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => simple_obj_ref_2905_inst_req_0); -- 
    ack_14615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2905_inst_ack_0, ack => cp_elements(269)); -- 
    cpelement_group_270 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(269) & cp_elements(272) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(270),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_14700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2904_gather_scatter_req_0); -- 
    cp_elements(271) <= cp_elements(267);
    req_14623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => simple_obj_ref_2903_inst_req_0); -- 
    cp_elements(272) <= simple_obj_ref_2903_inst_ack_0;
    cp_elements(273) <= cp_elements(272);
    base_resize_req_14631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2904_base_resize_req_0); -- 
    base_resize_ack_14632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_base_resize_ack_0, ack => cp_elements(274)); -- 
    sum_rename_req_14636_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => ptr_deref_2904_root_address_inst_req_0); -- 
    cp_elements(275) <= ptr_deref_2904_root_address_inst_ack_0;
    cp_elements(276) <= cp_elements(275);
    rr_14644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(276), ack => ptr_deref_2904_addr_0_req_0); -- 
    ra_14645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_0_ack_0, ack => cp_elements(277)); -- 
    cr_14646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2904_addr_0_req_1); -- 
    ca_14647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_0_ack_1, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(275);
    rr_14651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2904_addr_1_req_0); -- 
    ra_14652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_1_ack_0, ack => cp_elements(280)); -- 
    cr_14653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(280), ack => ptr_deref_2904_addr_1_req_1); -- 
    ca_14654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_1_ack_1, ack => cp_elements(281)); -- 
    cp_elements(282) <= cp_elements(275);
    rr_14658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2904_addr_2_req_0); -- 
    ra_14659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_2_ack_0, ack => cp_elements(283)); -- 
    cr_14660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => ptr_deref_2904_addr_2_req_1); -- 
    ca_14661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_2_ack_1, ack => cp_elements(284)); -- 
    cp_elements(285) <= cp_elements(275);
    rr_14665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(285), ack => ptr_deref_2904_addr_3_req_0); -- 
    ra_14666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_3_ack_0, ack => cp_elements(286)); -- 
    cr_14667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2904_addr_3_req_1); -- 
    ca_14668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_3_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(275);
    rr_14672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2904_addr_4_req_0); -- 
    ra_14673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_4_ack_0, ack => cp_elements(289)); -- 
    cr_14674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(289), ack => ptr_deref_2904_addr_4_req_1); -- 
    ca_14675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_4_ack_1, ack => cp_elements(290)); -- 
    cp_elements(291) <= cp_elements(275);
    rr_14679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(291), ack => ptr_deref_2904_addr_5_req_0); -- 
    ra_14680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_5_ack_0, ack => cp_elements(292)); -- 
    cr_14681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => ptr_deref_2904_addr_5_req_1); -- 
    ca_14682_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_5_ack_1, ack => cp_elements(293)); -- 
    cp_elements(294) <= cp_elements(275);
    rr_14686_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(294), ack => ptr_deref_2904_addr_6_req_0); -- 
    ra_14687_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_6_ack_0, ack => cp_elements(295)); -- 
    cr_14688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => ptr_deref_2904_addr_6_req_1); -- 
    ca_14689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_6_ack_1, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(275);
    rr_14693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(297), ack => ptr_deref_2904_addr_7_req_0); -- 
    ra_14694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_7_ack_0, ack => cp_elements(298)); -- 
    cr_14695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => ptr_deref_2904_addr_7_req_1); -- 
    ca_14696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_7_ack_1, ack => cp_elements(299)); -- 
    cpelement_group_300 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(278) & cp_elements(281) & cp_elements(284) & cp_elements(287) & cp_elements(290) & cp_elements(293) & cp_elements(296) & cp_elements(299));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(300),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(301) <= ptr_deref_2904_gather_scatter_ack_0;
    cp_elements(302) <= cp_elements(301);
    rr_14708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(302), ack => ptr_deref_2904_store_0_req_0); -- 
    ra_14709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_0_ack_0, ack => cp_elements(303)); -- 
    cp_elements(304) <= cp_elements(301);
    rr_14713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(304), ack => ptr_deref_2904_store_1_req_0); -- 
    ra_14714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_1_ack_0, ack => cp_elements(305)); -- 
    cp_elements(306) <= cp_elements(301);
    rr_14718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(306), ack => ptr_deref_2904_store_2_req_0); -- 
    ra_14719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_2_ack_0, ack => cp_elements(307)); -- 
    cp_elements(308) <= cp_elements(301);
    rr_14723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => ptr_deref_2904_store_3_req_0); -- 
    ra_14724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_3_ack_0, ack => cp_elements(309)); -- 
    cp_elements(310) <= cp_elements(301);
    rr_14728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(310), ack => ptr_deref_2904_store_4_req_0); -- 
    ra_14729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_4_ack_0, ack => cp_elements(311)); -- 
    cp_elements(312) <= cp_elements(301);
    rr_14733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(312), ack => ptr_deref_2904_store_5_req_0); -- 
    ra_14734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_5_ack_0, ack => cp_elements(313)); -- 
    cp_elements(314) <= cp_elements(301);
    rr_14738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(314), ack => ptr_deref_2904_store_6_req_0); -- 
    ra_14739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_6_ack_0, ack => cp_elements(315)); -- 
    cp_elements(316) <= cp_elements(301);
    rr_14743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => ptr_deref_2904_store_7_req_0); -- 
    ra_14744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_7_ack_0, ack => cp_elements(317)); -- 
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(303) & cp_elements(305) & cp_elements(307) & cp_elements(309) & cp_elements(311) & cp_elements(313) & cp_elements(315) & cp_elements(317));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(319) <= cp_elements(318);
    cr_14754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => ptr_deref_2904_store_0_req_1); -- 
    ca_14755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_0_ack_1, ack => cp_elements(320)); -- 
    cp_elements(321) <= cp_elements(318);
    cr_14759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => ptr_deref_2904_store_1_req_1); -- 
    ca_14760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_1_ack_1, ack => cp_elements(322)); -- 
    cp_elements(323) <= cp_elements(318);
    cr_14764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(323), ack => ptr_deref_2904_store_2_req_1); -- 
    ca_14765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_2_ack_1, ack => cp_elements(324)); -- 
    cp_elements(325) <= cp_elements(318);
    cr_14769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => ptr_deref_2904_store_3_req_1); -- 
    ca_14770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_3_ack_1, ack => cp_elements(326)); -- 
    cp_elements(327) <= cp_elements(318);
    cr_14774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(327), ack => ptr_deref_2904_store_4_req_1); -- 
    ca_14775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_4_ack_1, ack => cp_elements(328)); -- 
    cp_elements(329) <= cp_elements(318);
    cr_14779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => ptr_deref_2904_store_5_req_1); -- 
    ca_14780_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_5_ack_1, ack => cp_elements(330)); -- 
    cp_elements(331) <= cp_elements(318);
    cr_14784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => ptr_deref_2904_store_6_req_1); -- 
    ca_14785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_6_ack_1, ack => cp_elements(332)); -- 
    cp_elements(333) <= cp_elements(318);
    cr_14789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => ptr_deref_2904_store_7_req_1); -- 
    ca_14790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_store_7_ack_1, ack => cp_elements(334)); -- 
    cpelement_group_335 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(320) & cp_elements(322) & cp_elements(324) & cp_elements(326) & cp_elements(328) & cp_elements(330) & cp_elements(332) & cp_elements(334));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(335),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(336) <= cp_elements(335);
    cp_elements(337) <= false;
    cp_elements(338) <= cp_elements(337);
    cp_elements(339) <= cp_elements(335);
    req_14807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => simple_obj_ref_2908_inst_req_0); -- 
    ack_14808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2908_inst_ack_0, ack => cp_elements(340)); -- 
    rr_14809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => binary_2910_inst_req_0); -- 
    ra_14810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2910_inst_ack_0, ack => cp_elements(341)); -- 
    cr_14811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => binary_2910_inst_req_1); -- 
    ca_14812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2910_inst_ack_1, ack => cp_elements(342)); -- 
    branch_req_14813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(342), ack => if_stmt_2907_branch_req_0); -- 
    cp_elements(343) <= cp_elements(342);
    cp_elements(344) <= cp_elements(343);
    if_choice_transition_14818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2907_branch_ack_1, ack => cp_elements(345)); -- 
    cp_elements(346) <= cp_elements(343);
    else_choice_transition_14822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2907_branch_ack_0, ack => cp_elements(347)); -- 
    cp_elements(348) <= cp_elements(345);
    cpelement_group_349 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(350) & cp_elements(352));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(349),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(349), ack => type_cast_2913_inst_req_0); -- 
    cp_elements(350) <= cp_elements(348);
    cp_elements(351) <= cp_elements(348);
    req_14836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(351), ack => simple_obj_ref_2912_inst_req_0); -- 
    ack_14837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2912_inst_ack_0, ack => cp_elements(352)); -- 
    ack_14842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_0, ack => cp_elements(353)); -- 
    pipe_wreq_14847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => simple_obj_ref_2911_inst_req_0); -- 
    pipe_wack_14848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2911_inst_ack_0, ack => cp_elements(354)); -- 
    cp_elements(355) <= cp_elements(263);
    cp_elements(356) <= false;
    cp_elements(357) <= cp_elements(356);
    cp_elements(358) <= cp_elements(263);
    cp_elements(359) <= OrReduce(cp_elements(266) & cp_elements(358));
    cp_elements(360) <= cp_elements(359);
    cpelement_group_361 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(102) & cp_elements(146) & cp_elements(264));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(361),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_2857 : std_logic_vector(7 downto 0);
    signal NI_2874 : std_logic_vector(7 downto 0);
    signal a_2736 : std_logic_vector(63 downto 0);
    signal array_obj_ref_2792_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2792_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2792_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2882_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2882_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2882_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2882_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2882_wire : std_logic_vector(31 downto 0);
    signal binary_2742_wire : std_logic_vector(63 downto 0);
    signal binary_2744_wire : std_logic_vector(15 downto 0);
    signal binary_2747_wire : std_logic_vector(63 downto 0);
    signal binary_2751_wire : std_logic_vector(63 downto 0);
    signal binary_2753_wire : std_logic_vector(15 downto 0);
    signal binary_2754_wire : std_logic_vector(31 downto 0);
    signal binary_2757_wire : std_logic_vector(63 downto 0);
    signal binary_2761_wire : std_logic_vector(63 downto 0);
    signal binary_2763_wire : std_logic_vector(15 downto 0);
    signal binary_2766_wire : std_logic_vector(63 downto 0);
    signal binary_2770_wire : std_logic_vector(63 downto 0);
    signal binary_2772_wire : std_logic_vector(15 downto 0);
    signal binary_2773_wire : std_logic_vector(31 downto 0);
    signal binary_2774_wire : std_logic_vector(63 downto 0);
    signal binary_2842_wire : std_logic_vector(0 downto 0);
    signal binary_2887_wire : std_logic_vector(0 downto 0);
    signal binary_2896_wire : std_logic_vector(0 downto 0);
    signal binary_2910_wire : std_logic_vector(0 downto 0);
    signal buf64_ptr_2789 : std_logic_vector(31 downto 0);
    signal buf64_ptr_2822 : std_logic_vector(31 downto 0);
    signal buf8_ptr_2785 : std_logic_vector(31 downto 0);
    signal buf8_ptr_2819 : std_logic_vector(31 downto 0);
    signal buf_2781 : std_logic_vector(31 downto 0);
    signal expr_2741_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2746_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2750_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2756_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2760_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2765_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2769_wire_constant : std_logic_vector(63 downto 0);
    signal expr_2841_wire_constant : std_logic_vector(7 downto 0);
    signal expr_2850_wire_constant : std_logic_vector(0 downto 0);
    signal expr_2872_wire_constant : std_logic_vector(7 downto 0);
    signal expr_2886_wire_constant : std_logic_vector(7 downto 0);
    signal expr_2888_wire_constant : std_logic_vector(0 downto 0);
    signal expr_2889_wire_constant : std_logic_vector(0 downto 0);
    signal expr_2895_wire_constant : std_logic_vector(7 downto 0);
    signal expr_2909_wire_constant : std_logic_vector(0 downto 0);
    signal hdr_in_ctrl_2837 : std_logic_vector(7 downto 0);
    signal hdr_in_data_2834 : std_logic_vector(63 downto 0);
    signal pkt64_ptr_2828 : std_logic_vector(31 downto 0);
    signal pkt8_ptr_2793 : std_logic_vector(31 downto 0);
    signal pkt8_ptr_2825 : std_logic_vector(31 downto 0);
    signal pkt_in_ctrl_2869 : std_logic_vector(7 downto 0);
    signal pkt_in_data_2866 : std_logic_vector(63 downto 0);
    signal ptr_deref_2904_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_4 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_5 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_6 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_7 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2904_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_7 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_7 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2881_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2881_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2903_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_2905_wire : std_logic_vector(63 downto 0);
    signal simple_obj_ref_2908_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_2912_wire : std_logic_vector(31 downto 0);
    signal ternary_2890_wire : std_logic_vector(0 downto 0);
    signal type_cast_2739_wire : std_logic_vector(7 downto 0);
    signal type_cast_2743_wire : std_logic_vector(7 downto 0);
    signal type_cast_2748_wire : std_logic_vector(7 downto 0);
    signal type_cast_2752_wire : std_logic_vector(7 downto 0);
    signal type_cast_2758_wire : std_logic_vector(7 downto 0);
    signal type_cast_2762_wire : std_logic_vector(7 downto 0);
    signal type_cast_2767_wire : std_logic_vector(7 downto 0);
    signal type_cast_2771_wire : std_logic_vector(7 downto 0);
    signal type_cast_2809_wire : std_logic_vector(31 downto 0);
    signal type_cast_2860_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2913_wire : std_logic_vector(31 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxbuf64_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxbuf64_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxbuf8_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxbuf8_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxpkt64_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxpkt64_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxpkt8_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxpkt8_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxwrite_data
    signal xxreceive_packet_pipelinexxwrite_data_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxwrite_data
    signal xxreceive_packet_pipelinexxwrite_data_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxwrite_data_last_word_flag
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxwrite_data_last_word_flag
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxwrite_data_wptr
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxwrite_data_wptr
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_2792_final_offset <= "0000000010110100";
    array_obj_ref_2882_offset_scale_factor_0 <= "0000000000001000";
    expr_2741_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    expr_2746_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    expr_2750_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    expr_2756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    expr_2760_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    expr_2765_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    expr_2769_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    expr_2841_wire_constant <= "11111111";
    expr_2850_wire_constant <= "0";
    expr_2872_wire_constant <= "00000001";
    expr_2886_wire_constant <= "00000000";
    expr_2888_wire_constant <= "0";
    expr_2889_wire_constant <= "1";
    expr_2895_wire_constant <= "00000000";
    expr_2909_wire_constant <= "0";
    ptr_deref_2904_word_offset_0 <= "0000000000000000";
    ptr_deref_2904_word_offset_1 <= "0000000000000001";
    ptr_deref_2904_word_offset_2 <= "0000000000000010";
    ptr_deref_2904_word_offset_3 <= "0000000000000011";
    ptr_deref_2904_word_offset_4 <= "0000000000000100";
    ptr_deref_2904_word_offset_5 <= "0000000000000101";
    ptr_deref_2904_word_offset_6 <= "0000000000000110";
    ptr_deref_2904_word_offset_7 <= "0000000000000111";
    type_cast_2860_wire_constant <= "00000000";
    phi_stmt_2857: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2860_wire_constant & NI_2874;
      req <= phi_stmt_2857_req_0 & phi_stmt_2857_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2857_ack_0,
          idata => idata,
          odata => I_2857,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2857
    ternary_2890_inst: SelectBase generic map(data_width => 1) -- 
      port map( x => expr_2888_wire_constant, y => expr_2889_wire_constant, sel => binary_2887_wire, z => ternary_2890_wire, req => ternary_2890_inst_req_0, ack => ternary_2890_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2792_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => buf8_ptr_2785, dout => array_obj_ref_2792_resized_base_address, req => array_obj_ref_2792_base_resize_req_0, ack => array_obj_ref_2792_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2792_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2792_root_address, dout => pkt8_ptr_2793, req => array_obj_ref_2792_final_reg_req_0, ack => array_obj_ref_2792_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2882_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => pkt64_ptr_2828, dout => array_obj_ref_2882_resized_base_address, req => array_obj_ref_2882_base_resize_req_0, ack => array_obj_ref_2882_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2882_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2882_root_address, dout => array_obj_ref_2882_wire, req => array_obj_ref_2882_final_reg_req_0, ack => array_obj_ref_2882_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2882_index_0_resize: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 16, flow_through => true ) 
      port map( din => I_2857, dout => simple_obj_ref_2881_resized, req => array_obj_ref_2882_index_0_resize_req_0, ack => array_obj_ref_2882_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2882_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_2881_scaled, dout => array_obj_ref_2882_final_offset, req => array_obj_ref_2882_offset_inst_req_0, ack => array_obj_ref_2882_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2904_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_2903_wire, dout => ptr_deref_2904_resized_base_address, req => ptr_deref_2904_base_resize_req_0, ack => ptr_deref_2904_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2739_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => a_2736, dout => type_cast_2739_wire, req => type_cast_2739_inst_req_0, ack => type_cast_2739_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2743_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2742_wire, dout => type_cast_2743_wire, req => type_cast_2743_inst_req_0, ack => type_cast_2743_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2748_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2747_wire, dout => type_cast_2748_wire, req => type_cast_2748_inst_req_0, ack => type_cast_2748_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2752_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2751_wire, dout => type_cast_2752_wire, req => type_cast_2752_inst_req_0, ack => type_cast_2752_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2758_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2757_wire, dout => type_cast_2758_wire, req => type_cast_2758_inst_req_0, ack => type_cast_2758_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2762_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2761_wire, dout => type_cast_2762_wire, req => type_cast_2762_inst_req_0, ack => type_cast_2762_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2767_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2766_wire, dout => type_cast_2767_wire, req => type_cast_2767_inst_req_0, ack => type_cast_2767_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2771_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_2770_wire, dout => type_cast_2771_wire, req => type_cast_2771_inst_req_0, ack => type_cast_2771_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2784_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_2781, dout => buf8_ptr_2785, req => type_cast_2784_inst_req_0, ack => type_cast_2784_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2788_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_2781, dout => buf64_ptr_2789, req => type_cast_2788_inst_req_0, ack => type_cast_2788_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2809_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt8_ptr_2793, dout => type_cast_2809_wire, req => type_cast_2809_inst_req_0, ack => type_cast_2809_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2913_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => simple_obj_ref_2912_wire, dout => type_cast_2913_wire, req => type_cast_2913_inst_req_0, ack => type_cast_2913_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2904_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(63 downto 0); --
    begin -- 
      ptr_deref_2904_gather_scatter_ack_0 <= ptr_deref_2904_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_2905_wire;
      ptr_deref_2904_data_7 <= aggregated_sig(63 downto 56);
      ptr_deref_2904_data_6 <= aggregated_sig(55 downto 48);
      ptr_deref_2904_data_5 <= aggregated_sig(47 downto 40);
      ptr_deref_2904_data_4 <= aggregated_sig(39 downto 32);
      ptr_deref_2904_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_2904_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_2904_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2904_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2904_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2904_root_address_inst_ack_0 <= ptr_deref_2904_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2904_resized_base_address;
      ptr_deref_2904_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_2839_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_2842_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2839_branch_req_0,
          ack0 => if_stmt_2839_branch_ack_0,
          ack1 => if_stmt_2839_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2893_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_2896_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2893_branch_req_0,
          ack0 => if_stmt_2893_branch_ack_0,
          ack1 => if_stmt_2893_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2907_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_2910_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2907_branch_req_0,
          ack0 => if_stmt_2907_branch_ack_0,
          ack1 => if_stmt_2907_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_2792_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2792_resized_base_address;
      array_obj_ref_2792_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000010110100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2792_root_address_inst_req_0,
          ackL => array_obj_ref_2792_root_address_inst_ack_0,
          reqR => array_obj_ref_2792_root_address_inst_req_1,
          ackR => array_obj_ref_2792_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2882_index_0_scale 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2881_resized;
      simple_obj_ref_2881_scaled <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2882_index_0_scale_req_0,
          ackL => array_obj_ref_2882_index_0_scale_ack_0,
          reqR => array_obj_ref_2882_index_0_scale_req_1,
          ackR => array_obj_ref_2882_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_2882_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2882_final_offset & array_obj_ref_2882_resized_base_address;
      array_obj_ref_2882_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2882_root_address_inst_req_0,
          ackL => array_obj_ref_2882_root_address_inst_ack_0,
          reqR => array_obj_ref_2882_root_address_inst_req_1,
          ackR => array_obj_ref_2882_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2742_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2742_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2742_inst_req_0,
          ackL => binary_2742_inst_ack_0,
          reqR => binary_2742_inst_req_1,
          ackR => binary_2742_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2744_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2739_wire & type_cast_2743_wire;
      binary_2744_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2744_inst_req_0,
          ackL => binary_2744_inst_ack_0,
          reqR => binary_2744_inst_req_1,
          ackR => binary_2744_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2747_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2747_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2747_inst_req_0,
          ackL => binary_2747_inst_ack_0,
          reqR => binary_2747_inst_req_1,
          ackR => binary_2747_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2751_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2751_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2751_inst_req_0,
          ackL => binary_2751_inst_ack_0,
          reqR => binary_2751_inst_req_1,
          ackR => binary_2751_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2753_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2748_wire & type_cast_2752_wire;
      binary_2753_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2753_inst_req_0,
          ackL => binary_2753_inst_ack_0,
          reqR => binary_2753_inst_req_1,
          ackR => binary_2753_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2754_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_2744_wire & binary_2753_wire;
      binary_2754_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2754_inst_req_0,
          ackL => binary_2754_inst_ack_0,
          reqR => binary_2754_inst_req_1,
          ackR => binary_2754_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2757_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2757_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2757_inst_req_0,
          ackL => binary_2757_inst_ack_0,
          reqR => binary_2757_inst_req_1,
          ackR => binary_2757_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2761_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2761_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2761_inst_req_0,
          ackL => binary_2761_inst_ack_0,
          reqR => binary_2761_inst_req_1,
          ackR => binary_2761_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_2763_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2758_wire & type_cast_2762_wire;
      binary_2763_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2763_inst_req_0,
          ackL => binary_2763_inst_ack_0,
          reqR => binary_2763_inst_req_1,
          ackR => binary_2763_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_2766_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2766_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2766_inst_req_0,
          ackL => binary_2766_inst_ack_0,
          reqR => binary_2766_inst_req_1,
          ackR => binary_2766_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_2770_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_2736;
      binary_2770_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2770_inst_req_0,
          ackL => binary_2770_inst_ack_0,
          reqR => binary_2770_inst_req_1,
          ackR => binary_2770_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_2772_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2767_wire & type_cast_2771_wire;
      binary_2772_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2772_inst_req_0,
          ackL => binary_2772_inst_ack_0,
          reqR => binary_2772_inst_req_1,
          ackR => binary_2772_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_2773_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_2763_wire & binary_2772_wire;
      binary_2773_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2773_inst_req_0,
          ackL => binary_2773_inst_ack_0,
          reqR => binary_2773_inst_req_1,
          ackR => binary_2773_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_2774_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_2754_wire & binary_2773_wire;
      binary_2774_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2774_inst_req_0,
          ackL => binary_2774_inst_ack_0,
          reqR => binary_2774_inst_req_1,
          ackR => binary_2774_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_2842_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= hdr_in_ctrl_2837;
      binary_2842_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2842_inst_req_0,
          ackL => binary_2842_inst_ack_0,
          reqR => binary_2842_inst_req_1,
          ackR => binary_2842_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_2873_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_2857;
      NI_2874 <= data_out(7 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2873_inst_req_0,
          ackL => binary_2873_inst_ack_0,
          reqR => binary_2873_inst_req_1,
          ackR => binary_2873_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_2887_inst binary_2896_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= pkt_in_ctrl_2869 & pkt_in_ctrl_2869;
      binary_2887_wire <= data_out(1 downto 1);
      binary_2896_wire <= data_out(0 downto 0);
      reqL(1) <= binary_2887_inst_req_0;
      reqL(0) <= binary_2896_inst_req_0;
      binary_2887_inst_ack_0 <= ackL(1);
      binary_2896_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_2887_inst_req_1;
      reqR(0) <= binary_2896_inst_req_1;
      binary_2887_inst_ack_1 <= ackR(1);
      binary_2896_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_2910_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2908_wire;
      binary_2910_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2910_inst_req_0,
          ackL => binary_2910_inst_ack_0,
          reqR => binary_2910_inst_req_1,
          ackR => binary_2910_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2904_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_0_req_0,
          ackL => ptr_deref_2904_addr_0_ack_0,
          reqR => ptr_deref_2904_addr_0_req_1,
          ackR => ptr_deref_2904_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2904_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_1_req_0,
          ackL => ptr_deref_2904_addr_1_ack_0,
          reqR => ptr_deref_2904_addr_1_req_1,
          ackR => ptr_deref_2904_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2904_addr_2 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_2_req_0,
          ackL => ptr_deref_2904_addr_2_ack_0,
          reqR => ptr_deref_2904_addr_2_req_1,
          ackR => ptr_deref_2904_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2904_addr_3 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_3_req_0,
          ackL => ptr_deref_2904_addr_3_ack_0,
          reqR => ptr_deref_2904_addr_3_req_1,
          ackR => ptr_deref_2904_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2904_addr_4 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_4 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_4_req_0,
          ackL => ptr_deref_2904_addr_4_ack_0,
          reqR => ptr_deref_2904_addr_4_req_1,
          ackR => ptr_deref_2904_addr_4_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2904_addr_5 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_5 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000101",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_5_req_0,
          ackL => ptr_deref_2904_addr_5_ack_0,
          reqR => ptr_deref_2904_addr_5_req_1,
          ackR => ptr_deref_2904_addr_5_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2904_addr_6 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_6 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_6_req_0,
          ackL => ptr_deref_2904_addr_6_ack_0,
          reqR => ptr_deref_2904_addr_6_req_1,
          ackR => ptr_deref_2904_addr_6_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2904_addr_7 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_7 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_7_req_0,
          ackL => ptr_deref_2904_addr_7_ack_0,
          reqR => ptr_deref_2904_addr_7_req_1,
          ackR => ptr_deref_2904_addr_7_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2904_store_4_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_4 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_4) &  " data ptr_deref_2904_data_4 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_4) severity note; --
        end if;
        if ptr_deref_2904_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_3) &  " data ptr_deref_2904_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_3) severity note; --
        end if;
        if ptr_deref_2904_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_2) &  " data ptr_deref_2904_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_2) severity note; --
        end if;
        if ptr_deref_2904_store_5_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_5 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_5) &  " data ptr_deref_2904_data_5 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_5) severity note; --
        end if;
        if ptr_deref_2904_store_6_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_6 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_6) &  " data ptr_deref_2904_data_6 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_6) severity note; --
        end if;
        if ptr_deref_2904_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_0) &  " data ptr_deref_2904_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_0) severity note; --
        end if;
        if ptr_deref_2904_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_1) &  " data ptr_deref_2904_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_1) severity note; --
        end if;
        if ptr_deref_2904_store_7_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2904_word_address_7 ="  &  convert_slv_to_hex_string(ptr_deref_2904_word_address_7) &  " data ptr_deref_2904_data_7 ="  &  convert_slv_to_hex_string(ptr_deref_2904_data_7) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2904_store_4 ptr_deref_2904_store_3 ptr_deref_2904_store_2 ptr_deref_2904_store_5 ptr_deref_2904_store_6 ptr_deref_2904_store_0 ptr_deref_2904_store_1 ptr_deref_2904_store_7 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(127 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= ptr_deref_2904_store_4_req_0;
      reqL(6) <= ptr_deref_2904_store_3_req_0;
      reqL(5) <= ptr_deref_2904_store_2_req_0;
      reqL(4) <= ptr_deref_2904_store_5_req_0;
      reqL(3) <= ptr_deref_2904_store_6_req_0;
      reqL(2) <= ptr_deref_2904_store_0_req_0;
      reqL(1) <= ptr_deref_2904_store_1_req_0;
      reqL(0) <= ptr_deref_2904_store_7_req_0;
      ptr_deref_2904_store_4_ack_0 <= ackL(7);
      ptr_deref_2904_store_3_ack_0 <= ackL(6);
      ptr_deref_2904_store_2_ack_0 <= ackL(5);
      ptr_deref_2904_store_5_ack_0 <= ackL(4);
      ptr_deref_2904_store_6_ack_0 <= ackL(3);
      ptr_deref_2904_store_0_ack_0 <= ackL(2);
      ptr_deref_2904_store_1_ack_0 <= ackL(1);
      ptr_deref_2904_store_7_ack_0 <= ackL(0);
      reqR(7) <= ptr_deref_2904_store_4_req_1;
      reqR(6) <= ptr_deref_2904_store_3_req_1;
      reqR(5) <= ptr_deref_2904_store_2_req_1;
      reqR(4) <= ptr_deref_2904_store_5_req_1;
      reqR(3) <= ptr_deref_2904_store_6_req_1;
      reqR(2) <= ptr_deref_2904_store_0_req_1;
      reqR(1) <= ptr_deref_2904_store_1_req_1;
      reqR(0) <= ptr_deref_2904_store_7_req_1;
      ptr_deref_2904_store_4_ack_1 <= ackR(7);
      ptr_deref_2904_store_3_ack_1 <= ackR(6);
      ptr_deref_2904_store_2_ack_1 <= ackR(5);
      ptr_deref_2904_store_5_ack_1 <= ackR(4);
      ptr_deref_2904_store_6_ack_1 <= ackR(3);
      ptr_deref_2904_store_0_ack_1 <= ackR(2);
      ptr_deref_2904_store_1_ack_1 <= ackR(1);
      ptr_deref_2904_store_7_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2904_word_address_4 & ptr_deref_2904_word_address_3 & ptr_deref_2904_word_address_2 & ptr_deref_2904_word_address_5 & ptr_deref_2904_word_address_6 & ptr_deref_2904_word_address_0 & ptr_deref_2904_word_address_1 & ptr_deref_2904_word_address_7;
      data_in <= ptr_deref_2904_data_4 & ptr_deref_2904_data_3 & ptr_deref_2904_data_2 & ptr_deref_2904_data_5 & ptr_deref_2904_data_6 & ptr_deref_2904_data_0 & ptr_deref_2904_data_1 & ptr_deref_2904_data_7;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 8,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    xxreceive_packet_pipelinexxbuf64_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxbuf8_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxpkt64_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxpkt8_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxwrite_data_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxwrite_data_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxwrite_data_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxwrite_data_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxwrite_data_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxwrite_data_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxwrite_data_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxwrite_data_last_word_flag_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxwrite_data_wptr_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : simple_obj_ref_2735_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2735_inst_ack_0 then -- 
            assert false report " ReadPipe in_data to wire a_2736 value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2735_inst_req_0;
      simple_obj_ref_2735_inst_ack_0 <= ack(0);
      a_2736 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_2818_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2818_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxbuf8_ptr_pipe to wire buf8_ptr_2819 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2818_inst_req_0;
      simple_obj_ref_2818_inst_ack_0 <= ack(0);
      buf8_ptr_2819 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_2821_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2821_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxbuf64_ptr_pipe to wire buf64_ptr_2822 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2821_inst_req_0;
      simple_obj_ref_2821_inst_ack_0 <= ack(0);
      buf64_ptr_2822 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_2824_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2824_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxpkt8_ptr_pipe to wire pkt8_ptr_2825 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2824_inst_req_0;
      simple_obj_ref_2824_inst_ack_0 <= ack(0);
      pkt8_ptr_2825 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_2827_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2827_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxpkt64_ptr_pipe to wire pkt64_ptr_2828 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2827_inst_req_0;
      simple_obj_ref_2827_inst_ack_0 <= ack(0);
      pkt64_ptr_2828 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : simple_obj_ref_2865_inst simple_obj_ref_2833_inst 
    InportGroup5: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2865_inst_ack_0 then -- 
            assert false report " ReadPipe swapped_in_data to wire pkt_in_data_2866 value="  &  convert_slv_to_hex_string(data_out(127 downto 64))  severity note; --
          end if;
          if simple_obj_ref_2833_inst_ack_0 then -- 
            assert false report " ReadPipe swapped_in_data to wire hdr_in_data_2834 value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(1) <= simple_obj_ref_2865_inst_req_0;
      req(0) <= simple_obj_ref_2833_inst_req_0;
      simple_obj_ref_2865_inst_ack_0 <= ack(1);
      simple_obj_ref_2833_inst_ack_0 <= ack(0);
      pkt_in_data_2866 <= data_out(127 downto 64);
      hdr_in_data_2834 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 2,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => swapped_in_data_pipe_read_req(0),
          oack => swapped_in_data_pipe_read_ack(0),
          odata => swapped_in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : simple_obj_ref_2868_inst simple_obj_ref_2836_inst 
    InportGroup6: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2868_inst_ack_0 then -- 
            assert false report " ReadPipe in_ctrl to wire pkt_in_ctrl_2869 value="  &  convert_slv_to_hex_string(data_out(15 downto 8))  severity note; --
          end if;
          if simple_obj_ref_2836_inst_ack_0 then -- 
            assert false report " ReadPipe in_ctrl to wire hdr_in_ctrl_2837 value="  &  convert_slv_to_hex_string(data_out(7 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(1) <= simple_obj_ref_2868_inst_req_0;
      req(0) <= simple_obj_ref_2836_inst_req_0;
      simple_obj_ref_2868_inst_ack_0 <= ack(1);
      simple_obj_ref_2836_inst_ack_0 <= ack(0);
      pkt_in_ctrl_2869 <= data_out(15 downto 8);
      hdr_in_ctrl_2837 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 2,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_ctrl_pipe_read_req(0),
          oack => in_ctrl_pipe_read_ack(0),
          odata => in_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : simple_obj_ref_2903_inst 
    InportGroup7: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2903_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxwrite_data_wptr to wire simple_obj_ref_2903_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2903_inst_req_0;
      simple_obj_ref_2903_inst_ack_0 <= ack(0);
      simple_obj_ref_2903_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : simple_obj_ref_2905_inst 
    InportGroup8: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2905_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxwrite_data to wire simple_obj_ref_2905_wire value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2905_inst_req_0;
      simple_obj_ref_2905_inst_ack_0 <= ack(0);
      simple_obj_ref_2905_wire <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxwrite_data_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : simple_obj_ref_2908_inst 
    InportGroup9: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2908_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxwrite_data_last_word_flag to wire simple_obj_ref_2908_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2908_inst_req_0;
      simple_obj_ref_2908_inst_ack_0 <= ack(0);
      simple_obj_ref_2908_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : simple_obj_ref_2912_inst 
    InportGroup10: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2912_inst_ack_0 then -- 
            assert false report " ReadPipe receive_packet_buf_queue to wire simple_obj_ref_2912_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2912_inst_req_0;
      simple_obj_ref_2912_inst_ack_0 <= ack(0);
      simple_obj_ref_2912_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => receive_packet_buf_queue_pipe_read_req(0),
          oack => receive_packet_buf_queue_pipe_read_ack(0),
          odata => receive_packet_buf_queue_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2737_inst_ack_0 then -- 
          assert false report " WritePipe swapped_in_data from wire binary_2774_wire value="  &  convert_slv_to_hex_string(binary_2774_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2737_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2737_inst_req_0;
      simple_obj_ref_2737_inst_ack_0 <= ack(0);
      data_in <= binary_2774_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => swapped_in_data_pipe_write_req(0),
          oack => swapped_in_data_pipe_write_ack(0),
          odata => swapped_in_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2794_inst_ack_0 then -- 
          assert false report " WritePipe receive_packet_buf_queue from wire buf_2781 value="  &  convert_slv_to_hex_string(buf_2781) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2794_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2794_inst_req_0;
      simple_obj_ref_2794_inst_ack_0 <= ack(0);
      data_in <= buf_2781;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => receive_packet_buf_queue_pipe_write_req(0),
          oack => receive_packet_buf_queue_pipe_write_ack(0),
          odata => receive_packet_buf_queue_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2798_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxbuf8_ptr_pipe from wire buf8_ptr_2785 value="  &  convert_slv_to_hex_string(buf8_ptr_2785) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (2) : simple_obj_ref_2798_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2798_inst_req_0;
      simple_obj_ref_2798_inst_ack_0 <= ack(0);
      data_in <= buf8_ptr_2785;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2801_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxbuf64_ptr_pipe from wire buf64_ptr_2789 value="  &  convert_slv_to_hex_string(buf64_ptr_2789) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (3) : simple_obj_ref_2801_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2801_inst_req_0;
      simple_obj_ref_2801_inst_ack_0 <= ack(0);
      data_in <= buf64_ptr_2789;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2804_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxpkt8_ptr_pipe from wire pkt8_ptr_2793 value="  &  convert_slv_to_hex_string(pkt8_ptr_2793) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (4) : simple_obj_ref_2804_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2804_inst_req_0;
      simple_obj_ref_2804_inst_ack_0 <= ack(0);
      data_in <= pkt8_ptr_2793;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2807_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxpkt64_ptr_pipe from wire type_cast_2809_wire value="  &  convert_slv_to_hex_string(type_cast_2809_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (5) : simple_obj_ref_2807_inst 
    OutportGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2807_inst_req_0;
      simple_obj_ref_2807_inst_ack_0 <= ack(0);
      data_in <= type_cast_2809_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2846_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data from wire hdr_in_data_2834 value="  &  convert_slv_to_hex_string(hdr_in_data_2834) severity note; --
        end if;
        if simple_obj_ref_2877_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data from wire pkt_in_data_2866 value="  &  convert_slv_to_hex_string(pkt_in_data_2866) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (6) : simple_obj_ref_2846_inst simple_obj_ref_2877_inst 
    OutportGroup6: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_2846_inst_req_0;
      req(0) <= simple_obj_ref_2877_inst_req_0;
      simple_obj_ref_2846_inst_ack_0 <= ack(1);
      simple_obj_ref_2877_inst_ack_0 <= ack(0);
      data_in <= hdr_in_data_2834 & pkt_in_data_2866;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxwrite_data_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2849_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_last_word_flag from wire expr_2850_wire_constant value="  &  convert_slv_to_hex_string(expr_2850_wire_constant) severity note; --
        end if;
        if simple_obj_ref_2884_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_last_word_flag from wire ternary_2890_wire value="  &  convert_slv_to_hex_string(ternary_2890_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (7) : simple_obj_ref_2849_inst simple_obj_ref_2884_inst 
    OutportGroup7: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_2849_inst_req_0;
      req(0) <= simple_obj_ref_2884_inst_req_0;
      simple_obj_ref_2849_inst_ack_0 <= ack(1);
      simple_obj_ref_2884_inst_ack_0 <= ack(0);
      data_in <= expr_2850_wire_constant & ternary_2890_wire;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2852_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_wptr from wire buf64_ptr_2822 value="  &  convert_slv_to_hex_string(buf64_ptr_2822) severity note; --
        end if;
        if simple_obj_ref_2880_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_wptr from wire array_obj_ref_2882_wire value="  &  convert_slv_to_hex_string(array_obj_ref_2882_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (8) : simple_obj_ref_2852_inst simple_obj_ref_2880_inst 
    OutportGroup8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_2852_inst_req_0;
      req(0) <= simple_obj_ref_2880_inst_req_0;
      simple_obj_ref_2852_inst_ack_0 <= ack(1);
      simple_obj_ref_2880_inst_ack_0 <= ack(0);
      data_in <= buf64_ptr_2822 & array_obj_ref_2882_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2911_inst_ack_0 then -- 
          assert false report " WritePipe receive_packet_pipe from wire type_cast_2913_wire value="  &  convert_slv_to_hex_string(type_cast_2913_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (9) : simple_obj_ref_2911_inst 
    OutportGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2911_inst_req_0;
      simple_obj_ref_2911_inst_ack_0 <= ack(0);
      data_in <= type_cast_2913_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => receive_packet_pipe_pipe_write_req(0),
          oack => receive_packet_pipe_pipe_write_ack(0),
          odata => receive_packet_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 9
    -- shared call operator group (0) : call_stmt_2781_call 
    CallGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_2781_call_req_0;
      call_stmt_2781_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_2781_call_req_1;
      call_stmt_2781_call_ack_1 <= ackR(0);
      buf_2781 <= data_out(31 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => ahir_packet_get_call_reqs(0),
          ackR => ahir_packet_get_call_acks(0),
          tagR => ahir_packet_get_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 32, owidth => 32, twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_packet_get_return_acks(0), -- cross-over
          ackL => ahir_packet_get_return_reqs(0), -- cross-over
          dataL => ahir_packet_get_return_data(31 downto 0),
          tagL => ahir_packet_get_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity send_packet_pipeline is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    send_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
    send_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    send_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_packet_free_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_free_call_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_free_call_data : out  std_logic_vector(31 downto 0);
    ahir_packet_free_call_tag  :  out  std_logic_vector(2 downto 0);
    ahir_packet_free_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_packet_free_return_acks : in   std_logic_vector(0 downto 0);
    ahir_packet_free_return_tag :  in   std_logic_vector(2 downto 0);
    analyze_packet_call_reqs : out  std_logic_vector(0 downto 0);
    analyze_packet_call_acks : in   std_logic_vector(0 downto 0);
    analyze_packet_call_data : out  std_logic_vector(31 downto 0);
    analyze_packet_call_tag  :  out  std_logic_vector(0 downto 0);
    analyze_packet_return_reqs : out  std_logic_vector(0 downto 0);
    analyze_packet_return_acks : in   std_logic_vector(0 downto 0);
    analyze_packet_return_data : in   std_logic_vector(63 downto 0);
    analyze_packet_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity send_packet_pipeline;
architecture Default of send_packet_pipeline is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal send_packet_pipeline_CP_14864_start: Boolean;
  -- links between control-path and data-path
  signal binary_3094_inst_ack_0 : boolean;
  signal binary_3091_inst_ack_1 : boolean;
  signal binary_3101_inst_req_0 : boolean;
  signal binary_3108_inst_req_1 : boolean;
  signal simple_obj_ref_3123_inst_ack_0 : boolean;
  signal binary_3089_inst_ack_0 : boolean;
  signal binary_3089_inst_req_0 : boolean;
  signal binary_3100_inst_ack_0 : boolean;
  signal binary_3108_inst_ack_0 : boolean;
  signal binary_3094_inst_req_1 : boolean;
  signal binary_3120_inst_req_0 : boolean;
  signal binary_3089_inst_ack_1 : boolean;
  signal simple_obj_ref_3124_inst_req_0 : boolean;
  signal binary_3108_inst_req_0 : boolean;
  signal binary_3100_inst_req_1 : boolean;
  signal simple_obj_ref_3084_inst_req_0 : boolean;
  signal binary_3108_inst_ack_1 : boolean;
  signal binary_3110_inst_ack_1 : boolean;
  signal binary_3130_inst_ack_1 : boolean;
  signal binary_3100_inst_ack_1 : boolean;
  signal binary_3101_inst_ack_1 : boolean;
  signal simple_obj_ref_3124_inst_ack_0 : boolean;
  signal binary_3120_inst_ack_0 : boolean;
  signal binary_3089_inst_req_1 : boolean;
  signal type_cast_3086_inst_req_0 : boolean;
  signal binary_3101_inst_ack_0 : boolean;
  signal type_cast_3090_inst_req_0 : boolean;
  signal binary_3101_inst_req_1 : boolean;
  signal simple_obj_ref_3123_inst_req_0 : boolean;
  signal binary_3120_inst_req_1 : boolean;
  signal binary_3094_inst_ack_1 : boolean;
  signal binary_3121_inst_req_1 : boolean;
  signal type_cast_3086_inst_ack_0 : boolean;
  signal binary_3120_inst_ack_1 : boolean;
  signal type_cast_3105_inst_ack_0 : boolean;
  signal binary_3121_inst_ack_0 : boolean;
  signal if_stmt_3127_branch_req_0 : boolean;
  signal binary_3121_inst_ack_1 : boolean;
  signal type_cast_3090_inst_ack_0 : boolean;
  signal binary_3091_inst_ack_0 : boolean;
  signal simple_obj_ref_3084_inst_ack_0 : boolean;
  signal binary_3091_inst_req_0 : boolean;
  signal binary_3121_inst_req_0 : boolean;
  signal type_cast_3105_inst_req_0 : boolean;
  signal binary_3119_inst_ack_1 : boolean;
  signal binary_3119_inst_req_1 : boolean;
  signal binary_3119_inst_ack_0 : boolean;
  signal binary_3100_inst_req_0 : boolean;
  signal type_cast_3099_inst_ack_0 : boolean;
  signal binary_3119_inst_req_0 : boolean;
  signal binary_3130_inst_req_1 : boolean;
  signal binary_3094_inst_req_0 : boolean;
  signal type_cast_3118_inst_req_0 : boolean;
  signal phi_stmt_3002_ack_0 : boolean;
  signal binary_3117_inst_ack_1 : boolean;
  signal phi_stmt_3002_req_0 : boolean;
  signal binary_3117_inst_req_1 : boolean;
  signal binary_3117_inst_ack_0 : boolean;
  signal type_cast_3099_inst_req_0 : boolean;
  signal phi_stmt_3002_req_1 : boolean;
  signal binary_3117_inst_req_0 : boolean;
  signal binary_3113_inst_req_1 : boolean;
  signal type_cast_3095_inst_ack_0 : boolean;
  signal binary_3104_inst_ack_1 : boolean;
  signal type_cast_3118_inst_ack_0 : boolean;
  signal binary_3113_inst_ack_1 : boolean;
  signal type_cast_3114_inst_ack_0 : boolean;
  signal type_cast_3114_inst_req_0 : boolean;
  signal binary_3104_inst_req_0 : boolean;
  signal type_cast_3109_inst_req_0 : boolean;
  signal binary_3104_inst_ack_0 : boolean;
  signal binary_3091_inst_req_1 : boolean;
  signal type_cast_3109_inst_ack_0 : boolean;
  signal binary_3104_inst_req_1 : boolean;
  signal type_cast_3095_inst_req_0 : boolean;
  signal simple_obj_ref_2935_inst_req_0 : boolean;
  signal simple_obj_ref_2935_inst_ack_0 : boolean;
  signal type_cast_2938_inst_req_0 : boolean;
  signal type_cast_2938_inst_ack_0 : boolean;
  signal call_stmt_2942_call_req_0 : boolean;
  signal call_stmt_2942_call_ack_0 : boolean;
  signal call_stmt_2942_call_req_1 : boolean;
  signal call_stmt_2942_call_ack_1 : boolean;
  signal type_cast_2946_inst_req_0 : boolean;
  signal type_cast_2946_inst_ack_0 : boolean;
  signal simple_obj_ref_2944_inst_req_0 : boolean;
  signal simple_obj_ref_2944_inst_ack_0 : boolean;
  signal type_cast_2950_inst_req_0 : boolean;
  signal type_cast_2950_inst_ack_0 : boolean;
  signal simple_obj_ref_2948_inst_req_0 : boolean;
  signal simple_obj_ref_2948_inst_ack_0 : boolean;
  signal simple_obj_ref_2952_inst_req_0 : boolean;
  signal simple_obj_ref_2952_inst_ack_0 : boolean;
  signal simple_obj_ref_2955_inst_req_0 : boolean;
  signal simple_obj_ref_2955_inst_ack_0 : boolean;
  signal type_cast_2960_inst_req_0 : boolean;
  signal type_cast_2960_inst_ack_0 : boolean;
  signal simple_obj_ref_2958_inst_req_0 : boolean;
  signal simple_obj_ref_2958_inst_ack_0 : boolean;
  signal simple_obj_ref_2969_inst_req_0 : boolean;
  signal simple_obj_ref_2969_inst_ack_0 : boolean;
  signal simple_obj_ref_2972_inst_req_0 : boolean;
  signal simple_obj_ref_2972_inst_ack_0 : boolean;
  signal simple_obj_ref_2975_inst_req_0 : boolean;
  signal simple_obj_ref_2975_inst_ack_0 : boolean;
  signal simple_obj_ref_2978_inst_req_0 : boolean;
  signal simple_obj_ref_2978_inst_ack_0 : boolean;
  signal binary_2984_inst_req_0 : boolean;
  signal binary_2984_inst_ack_0 : boolean;
  signal binary_2984_inst_req_1 : boolean;
  signal binary_2984_inst_ack_1 : boolean;
  signal if_stmt_2981_branch_req_0 : boolean;
  signal if_stmt_2981_branch_ack_1 : boolean;
  signal if_stmt_2981_branch_ack_0 : boolean;
  signal simple_obj_ref_2986_inst_req_0 : boolean;
  signal simple_obj_ref_2986_inst_ack_0 : boolean;
  signal simple_obj_ref_2989_inst_req_0 : boolean;
  signal simple_obj_ref_2989_inst_ack_0 : boolean;
  signal simple_obj_ref_2992_inst_req_0 : boolean;
  signal simple_obj_ref_2992_inst_ack_0 : boolean;
  signal binary_2998_inst_req_0 : boolean;
  signal binary_2998_inst_ack_0 : boolean;
  signal binary_2998_inst_req_1 : boolean;
  signal binary_2998_inst_ack_1 : boolean;
  signal simple_obj_ref_3009_inst_req_0 : boolean;
  signal simple_obj_ref_3009_inst_ack_0 : boolean;
  signal array_obj_ref_3014_index_0_resize_req_0 : boolean;
  signal array_obj_ref_3014_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_3014_index_0_scale_req_0 : boolean;
  signal array_obj_ref_3014_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_3014_index_0_scale_req_1 : boolean;
  signal array_obj_ref_3014_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_3014_offset_inst_req_0 : boolean;
  signal array_obj_ref_3014_offset_inst_ack_0 : boolean;
  signal array_obj_ref_3014_base_resize_req_0 : boolean;
  signal array_obj_ref_3014_base_resize_ack_0 : boolean;
  signal array_obj_ref_3014_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3014_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3014_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3014_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3014_final_reg_req_0 : boolean;
  signal array_obj_ref_3014_final_reg_ack_0 : boolean;
  signal simple_obj_ref_3012_inst_req_0 : boolean;
  signal simple_obj_ref_3012_inst_ack_0 : boolean;
  signal simple_obj_ref_3016_inst_req_0 : boolean;
  signal simple_obj_ref_3016_inst_ack_0 : boolean;
  signal binary_3022_inst_req_0 : boolean;
  signal binary_3022_inst_ack_0 : boolean;
  signal binary_3022_inst_req_1 : boolean;
  signal binary_3022_inst_ack_1 : boolean;
  signal binary_3028_inst_req_0 : boolean;
  signal binary_3028_inst_ack_0 : boolean;
  signal binary_3028_inst_req_1 : boolean;
  signal binary_3028_inst_ack_1 : boolean;
  signal if_stmt_3025_branch_req_0 : boolean;
  signal if_stmt_3025_branch_ack_1 : boolean;
  signal if_stmt_3025_branch_ack_0 : boolean;
  signal array_obj_ref_3033_index_0_resize_req_0 : boolean;
  signal array_obj_ref_3033_index_0_resize_ack_0 : boolean;
  signal binary_3110_inst_req_1 : boolean;
  signal binary_3110_inst_ack_0 : boolean;
  signal array_obj_ref_3033_index_0_scale_req_0 : boolean;
  signal array_obj_ref_3033_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_3033_index_0_scale_req_1 : boolean;
  signal array_obj_ref_3033_index_0_scale_ack_1 : boolean;
  signal binary_3110_inst_req_0 : boolean;
  signal array_obj_ref_3033_offset_inst_req_0 : boolean;
  signal array_obj_ref_3033_offset_inst_ack_0 : boolean;
  signal array_obj_ref_3033_base_resize_req_0 : boolean;
  signal array_obj_ref_3033_base_resize_ack_0 : boolean;
  signal array_obj_ref_3033_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3033_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3033_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3033_root_address_inst_ack_1 : boolean;
  signal binary_3130_inst_ack_0 : boolean;
  signal binary_3130_inst_req_0 : boolean;
  signal simple_obj_ref_3128_inst_ack_0 : boolean;
  signal simple_obj_ref_3128_inst_req_0 : boolean;
  signal array_obj_ref_3033_final_reg_req_0 : boolean;
  signal array_obj_ref_3033_final_reg_ack_0 : boolean;
  signal binary_3042_inst_req_0 : boolean;
  signal binary_3042_inst_ack_0 : boolean;
  signal binary_3042_inst_req_1 : boolean;
  signal binary_3042_inst_ack_1 : boolean;
  signal binary_3043_inst_req_0 : boolean;
  signal binary_3043_inst_ack_0 : boolean;
  signal binary_3043_inst_req_1 : boolean;
  signal binary_3043_inst_ack_1 : boolean;
  signal binary_3045_inst_req_0 : boolean;
  signal binary_3045_inst_ack_0 : boolean;
  signal binary_3045_inst_req_1 : boolean;
  signal binary_3045_inst_ack_1 : boolean;
  signal type_cast_3046_inst_req_0 : boolean;
  signal type_cast_3046_inst_ack_0 : boolean;
  signal binary_3047_inst_req_0 : boolean;
  signal binary_3047_inst_ack_0 : boolean;
  signal binary_3047_inst_req_1 : boolean;
  signal binary_3047_inst_ack_1 : boolean;
  signal simple_obj_ref_3036_inst_req_0 : boolean;
  signal simple_obj_ref_3036_inst_ack_0 : boolean;
  signal simple_obj_ref_3049_inst_req_0 : boolean;
  signal simple_obj_ref_3049_inst_ack_0 : boolean;
  signal simple_obj_ref_3052_inst_req_0 : boolean;
  signal simple_obj_ref_3052_inst_ack_0 : boolean;
  signal simple_obj_ref_3062_inst_req_0 : boolean;
  signal simple_obj_ref_3062_inst_ack_0 : boolean;
  signal ptr_deref_3067_base_resize_req_0 : boolean;
  signal ptr_deref_3067_base_resize_ack_0 : boolean;
  signal ptr_deref_3067_root_address_inst_req_0 : boolean;
  signal ptr_deref_3067_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3067_addr_0_req_0 : boolean;
  signal ptr_deref_3067_addr_0_ack_0 : boolean;
  signal ptr_deref_3067_addr_0_req_1 : boolean;
  signal ptr_deref_3067_addr_0_ack_1 : boolean;
  signal ptr_deref_3067_addr_1_req_0 : boolean;
  signal ptr_deref_3067_addr_1_ack_0 : boolean;
  signal ptr_deref_3067_addr_1_req_1 : boolean;
  signal ptr_deref_3067_addr_1_ack_1 : boolean;
  signal ptr_deref_3067_addr_2_req_0 : boolean;
  signal ptr_deref_3067_addr_2_ack_0 : boolean;
  signal ptr_deref_3067_addr_2_req_1 : boolean;
  signal ptr_deref_3067_addr_2_ack_1 : boolean;
  signal ptr_deref_3067_addr_3_req_0 : boolean;
  signal ptr_deref_3067_addr_3_ack_0 : boolean;
  signal ptr_deref_3067_addr_3_req_1 : boolean;
  signal ptr_deref_3067_addr_3_ack_1 : boolean;
  signal ptr_deref_3067_addr_4_req_0 : boolean;
  signal ptr_deref_3067_addr_4_ack_0 : boolean;
  signal ptr_deref_3067_addr_4_req_1 : boolean;
  signal ptr_deref_3067_addr_4_ack_1 : boolean;
  signal ptr_deref_3067_addr_5_req_0 : boolean;
  signal ptr_deref_3067_addr_5_ack_0 : boolean;
  signal ptr_deref_3067_addr_5_req_1 : boolean;
  signal ptr_deref_3067_addr_5_ack_1 : boolean;
  signal ptr_deref_3067_addr_6_req_0 : boolean;
  signal call_stmt_3132_call_ack_1 : boolean;
  signal ptr_deref_3067_addr_6_ack_0 : boolean;
  signal binary_3113_inst_ack_0 : boolean;
  signal ptr_deref_3067_addr_6_req_1 : boolean;
  signal ptr_deref_3067_addr_6_ack_1 : boolean;
  signal ptr_deref_3067_addr_7_req_0 : boolean;
  signal call_stmt_3132_call_req_1 : boolean;
  signal ptr_deref_3067_addr_7_ack_0 : boolean;
  signal binary_3113_inst_req_0 : boolean;
  signal ptr_deref_3067_addr_7_req_1 : boolean;
  signal ptr_deref_3067_addr_7_ack_1 : boolean;
  signal ptr_deref_3067_load_0_req_0 : boolean;
  signal ptr_deref_3067_load_0_ack_0 : boolean;
  signal ptr_deref_3067_load_1_req_0 : boolean;
  signal ptr_deref_3067_load_1_ack_0 : boolean;
  signal ptr_deref_3067_load_2_req_0 : boolean;
  signal ptr_deref_3067_load_2_ack_0 : boolean;
  signal ptr_deref_3067_load_3_req_0 : boolean;
  signal call_stmt_3132_call_ack_0 : boolean;
  signal ptr_deref_3067_load_3_ack_0 : boolean;
  signal ptr_deref_3067_load_4_req_0 : boolean;
  signal call_stmt_3132_call_req_0 : boolean;
  signal ptr_deref_3067_load_4_ack_0 : boolean;
  signal ptr_deref_3067_load_5_req_0 : boolean;
  signal ptr_deref_3067_load_5_ack_0 : boolean;
  signal ptr_deref_3067_load_6_req_0 : boolean;
  signal ptr_deref_3067_load_6_ack_0 : boolean;
  signal ptr_deref_3067_load_7_req_0 : boolean;
  signal ptr_deref_3067_load_7_ack_0 : boolean;
  signal ptr_deref_3067_load_0_req_1 : boolean;
  signal ptr_deref_3067_load_0_ack_1 : boolean;
  signal ptr_deref_3067_load_1_req_1 : boolean;
  signal ptr_deref_3067_load_1_ack_1 : boolean;
  signal ptr_deref_3067_load_2_req_1 : boolean;
  signal simple_obj_ref_3131_inst_ack_0 : boolean;
  signal ptr_deref_3067_load_2_ack_1 : boolean;
  signal ptr_deref_3067_load_3_req_1 : boolean;
  signal simple_obj_ref_3131_inst_req_0 : boolean;
  signal ptr_deref_3067_load_3_ack_1 : boolean;
  signal ptr_deref_3067_load_4_req_1 : boolean;
  signal ptr_deref_3067_load_4_ack_1 : boolean;
  signal ptr_deref_3067_load_5_req_1 : boolean;
  signal ptr_deref_3067_load_5_ack_1 : boolean;
  signal ptr_deref_3067_load_6_req_1 : boolean;
  signal ptr_deref_3067_load_6_ack_1 : boolean;
  signal ptr_deref_3067_load_7_req_1 : boolean;
  signal ptr_deref_3067_load_7_ack_1 : boolean;
  signal ptr_deref_3067_gather_scatter_req_0 : boolean;
  signal ptr_deref_3067_gather_scatter_ack_0 : boolean;
  signal binary_3098_inst_ack_1 : boolean;
  signal simple_obj_ref_3065_inst_req_0 : boolean;
  signal simple_obj_ref_3065_inst_ack_0 : boolean;
  signal simple_obj_ref_3070_inst_req_0 : boolean;
  signal if_stmt_3127_branch_ack_0 : boolean;
  signal simple_obj_ref_3070_inst_ack_0 : boolean;
  signal binary_3098_inst_req_1 : boolean;
  signal simple_obj_ref_3069_inst_req_0 : boolean;
  signal simple_obj_ref_3069_inst_ack_0 : boolean;
  signal simple_obj_ref_3073_inst_req_0 : boolean;
  signal simple_obj_ref_3073_inst_ack_0 : boolean;
  signal binary_3098_inst_ack_0 : boolean;
  signal simple_obj_ref_3072_inst_req_0 : boolean;
  signal simple_obj_ref_3072_inst_ack_0 : boolean;
  signal if_stmt_3127_branch_ack_1 : boolean;
  signal binary_3098_inst_req_0 : boolean;
  signal simple_obj_ref_3081_inst_req_0 : boolean;
  signal simple_obj_ref_3081_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  send_packet_pipeline_CP_14864: Block -- control-path 
    signal cp_elements: BooleanArray(388 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(388);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(388), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    cp_elements(2) <= false; 
    cp_elements(3) <= OrReduce(cp_elements(39) & cp_elements(42));
    req_14893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2935_inst_req_0); -- 
    cp_elements(4) <= cp_elements(36);
    ack_14894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2935_inst_ack_0, ack => cp_elements(5)); -- 
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(8) & cp_elements(9));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => type_cast_2938_inst_req_0); -- 
    cp_elements(8) <= cp_elements(6);
    cp_elements(9) <= cp_elements(6);
    ack_14905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2938_inst_ack_0, ack => cp_elements(10)); -- 
    crr_14911_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => call_stmt_2942_call_req_0); -- 
    cra_14912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2942_call_ack_0, ack => cp_elements(11)); -- 
    ccr_14916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => call_stmt_2942_call_req_1); -- 
    cca_14917_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2942_call_ack_1, ack => cp_elements(12)); -- 
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= cp_elements(13);
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => type_cast_2946_inst_req_0); -- 
    cp_elements(16) <= cp_elements(14);
    cp_elements(17) <= cp_elements(14);
    ack_14935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2946_inst_ack_0, ack => cp_elements(18)); -- 
    pipe_wreq_14940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => simple_obj_ref_2944_inst_req_0); -- 
    pipe_wack_14941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2944_inst_ack_0, ack => cp_elements(19)); -- 
    cp_elements(20) <= cp_elements(13);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14953_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => type_cast_2950_inst_req_0); -- 
    cp_elements(22) <= cp_elements(20);
    cp_elements(23) <= cp_elements(20);
    ack_14954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2950_inst_ack_0, ack => cp_elements(24)); -- 
    pipe_wreq_14959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => simple_obj_ref_2948_inst_req_0); -- 
    pipe_wack_14960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2948_inst_ack_0, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(13);
    pipe_wreq_14971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => simple_obj_ref_2952_inst_req_0); -- 
    pipe_wack_14972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2952_inst_ack_0, ack => cp_elements(27)); -- 
    cp_elements(28) <= cp_elements(13);
    pipe_wreq_14983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => simple_obj_ref_2955_inst_req_0); -- 
    pipe_wack_14984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2955_inst_ack_0, ack => cp_elements(29)); -- 
    cp_elements(30) <= cp_elements(13);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(33));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => type_cast_2960_inst_req_0); -- 
    cp_elements(32) <= cp_elements(30);
    cp_elements(33) <= cp_elements(30);
    ack_14997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2960_inst_ack_0, ack => cp_elements(34)); -- 
    pipe_wreq_15002_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => simple_obj_ref_2958_inst_req_0); -- 
    pipe_wack_15003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2958_inst_ack_0, ack => cp_elements(35)); -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(25) & cp_elements(27) & cp_elements(29) & cp_elements(35));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(37) <= cp_elements(1);
    cp_elements(38) <= false;
    cp_elements(39) <= cp_elements(38);
    cp_elements(40) <= cp_elements(1);
    cp_elements(41) <= OrReduce(cp_elements(4) & cp_elements(40));
    cp_elements(42) <= cp_elements(41);
    cp_elements(43) <= cp_elements(0);
    cp_elements(44) <= false; 
    cp_elements(45) <= OrReduce(cp_elements(177) & cp_elements(180));
    cp_elements(46) <= cp_elements(57);
    cp_elements(47) <= OrReduce(cp_elements(60) & cp_elements(68) & cp_elements(73));
    cp_elements(48) <= cp_elements(45);
    cp_elements(49) <= cp_elements(48);
    req_15043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => simple_obj_ref_2969_inst_req_0); -- 
    ack_15044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2969_inst_ack_0, ack => cp_elements(50)); -- 
    cp_elements(51) <= cp_elements(48);
    req_15054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => simple_obj_ref_2972_inst_req_0); -- 
    ack_15055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2972_inst_ack_0, ack => cp_elements(52)); -- 
    cp_elements(53) <= cp_elements(48);
    req_15065_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => simple_obj_ref_2975_inst_req_0); -- 
    ack_15066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2975_inst_ack_0, ack => cp_elements(54)); -- 
    cp_elements(55) <= cp_elements(48);
    req_15076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => simple_obj_ref_2978_inst_req_0); -- 
    ack_15077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2978_inst_ack_0, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(52) & cp_elements(54) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(58) <= cp_elements(46);
    cp_elements(59) <= false;
    cp_elements(60) <= cp_elements(59);
    cp_elements(61) <= cp_elements(46);
    rr_15091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => binary_2984_inst_req_0); -- 
    ra_15092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2984_inst_ack_0, ack => cp_elements(62)); -- 
    cr_15093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => binary_2984_inst_req_1); -- 
    ca_15094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2984_inst_ack_1, ack => cp_elements(63)); -- 
    branch_req_15095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => if_stmt_2981_branch_req_0); -- 
    cp_elements(64) <= cp_elements(63);
    cp_elements(65) <= cp_elements(64);
    if_choice_transition_15100_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2981_branch_ack_1, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(64);
    else_choice_transition_15104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2981_branch_ack_0, ack => cp_elements(68)); -- 
    cp_elements(69) <= cp_elements(87);
    cp_elements(70) <= OrReduce(cp_elements(170) & cp_elements(174));
    cp_elements(71) <= cp_elements(114);
    cp_elements(72) <= OrReduce(cp_elements(117) & cp_elements(125));
    cp_elements(73) <= cp_elements(167);
    cp_elements(74) <= cp_elements(66);
    cp_elements(75) <= cp_elements(74);
    pipe_wreq_15129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => simple_obj_ref_2986_inst_req_0); -- 
    pipe_wack_15130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2986_inst_ack_0, ack => cp_elements(76)); -- 
    cp_elements(77) <= cp_elements(74);
    pipe_wreq_15141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => simple_obj_ref_2989_inst_req_0); -- 
    pipe_wack_15142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2989_inst_ack_0, ack => cp_elements(78)); -- 
    cp_elements(79) <= cp_elements(74);
    pipe_wreq_15152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => simple_obj_ref_2992_inst_req_0); -- 
    pipe_wack_15153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2992_inst_ack_0, ack => cp_elements(80)); -- 
    cp_elements(81) <= cp_elements(74);
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => binary_2998_inst_req_0); -- 
    cp_elements(83) <= cp_elements(81);
    cp_elements(84) <= cp_elements(81);
    ra_15166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2998_inst_ack_0, ack => cp_elements(85)); -- 
    cr_15167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => binary_2998_inst_req_1); -- 
    ca_15168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2998_inst_ack_1, ack => cp_elements(86)); -- 
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(78) & cp_elements(80) & cp_elements(86));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(88) <= cp_elements(70);
    cp_elements(89) <= cp_elements(88);
    pipe_wreq_15181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => simple_obj_ref_3009_inst_req_0); -- 
    pipe_wack_15182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3009_inst_ack_0, ack => cp_elements(90)); -- 
    cp_elements(91) <= cp_elements(88);
    cp_elements(92) <= cp_elements(91);
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(92) & cp_elements(103));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_15231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => array_obj_ref_3014_final_reg_req_0); -- 
    cp_elements(94) <= cp_elements(91);
    base_resize_req_15218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => array_obj_ref_3014_base_resize_req_0); -- 
    cp_elements(95) <= cp_elements(91);
    index_resize_req_15200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_3014_index_0_resize_req_0); -- 
    index_resize_ack_15201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_index_0_resize_ack_0, ack => cp_elements(96)); -- 
    scale_rr_15205_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => array_obj_ref_3014_index_0_scale_req_0); -- 
    scale_ra_15206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_index_0_scale_ack_0, ack => cp_elements(97)); -- 
    scale_cr_15207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => array_obj_ref_3014_index_0_scale_req_1); -- 
    scale_ca_15208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_index_0_scale_ack_1, ack => cp_elements(98)); -- 
    final_index_req_15212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_3014_offset_inst_req_0); -- 
    final_index_ack_15213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_offset_inst_ack_0, ack => cp_elements(99)); -- 
    base_resize_ack_15219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_base_resize_ack_0, ack => cp_elements(100)); -- 
    cpelement_group_101 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(99) & cp_elements(100));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(101),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_15224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => array_obj_ref_3014_root_address_inst_req_0); -- 
    plus_base_ra_15225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_root_address_inst_ack_0, ack => cp_elements(102)); -- 
    plus_base_cr_15226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => array_obj_ref_3014_root_address_inst_req_1); -- 
    plus_base_ca_15227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_root_address_inst_ack_1, ack => cp_elements(103)); -- 
    final_reg_ack_15232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3014_final_reg_ack_0, ack => cp_elements(104)); -- 
    pipe_wreq_15237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => simple_obj_ref_3012_inst_req_0); -- 
    pipe_wack_15238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3012_inst_ack_0, ack => cp_elements(105)); -- 
    cp_elements(106) <= cp_elements(88);
    pipe_wreq_15248_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => simple_obj_ref_3016_inst_req_0); -- 
    pipe_wack_15249_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3016_inst_ack_0, ack => cp_elements(107)); -- 
    cp_elements(108) <= cp_elements(88);
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(111));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => binary_3022_inst_req_0); -- 
    cp_elements(110) <= cp_elements(108);
    cp_elements(111) <= cp_elements(108);
    ra_15262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3022_inst_ack_0, ack => cp_elements(112)); -- 
    cr_15263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => binary_3022_inst_req_1); -- 
    ca_15264_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3022_inst_ack_1, ack => cp_elements(113)); -- 
    cpelement_group_114 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(90) & cp_elements(105) & cp_elements(107) & cp_elements(113));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(114),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(115) <= cp_elements(71);
    cp_elements(116) <= false;
    cp_elements(117) <= cp_elements(116);
    cp_elements(118) <= cp_elements(71);
    rr_15278_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => binary_3028_inst_req_0); -- 
    ra_15279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3028_inst_ack_0, ack => cp_elements(119)); -- 
    cr_15280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => binary_3028_inst_req_1); -- 
    ca_15281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3028_inst_ack_1, ack => cp_elements(120)); -- 
    branch_req_15282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => if_stmt_3025_branch_req_0); -- 
    cp_elements(121) <= cp_elements(120);
    cp_elements(122) <= cp_elements(121);
    if_choice_transition_15287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3025_branch_ack_1, ack => cp_elements(123)); -- 
    phi_stmt_3002_req_15447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => phi_stmt_3002_req_1); -- 
    cp_elements(124) <= cp_elements(121);
    else_choice_transition_15291_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3025_branch_ack_0, ack => cp_elements(125)); -- 
    cp_elements(126) <= cp_elements(72);
    cp_elements(127) <= cp_elements(126);
    cpelement_group_128 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(138));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(128),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_15341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => array_obj_ref_3033_final_reg_req_0); -- 
    cp_elements(129) <= cp_elements(126);
    base_resize_req_15328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => array_obj_ref_3033_base_resize_req_0); -- 
    cp_elements(130) <= cp_elements(126);
    index_resize_req_15310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => array_obj_ref_3033_index_0_resize_req_0); -- 
    index_resize_ack_15311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_index_0_resize_ack_0, ack => cp_elements(131)); -- 
    scale_rr_15315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => array_obj_ref_3033_index_0_scale_req_0); -- 
    scale_ra_15316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_index_0_scale_ack_0, ack => cp_elements(132)); -- 
    scale_cr_15317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => array_obj_ref_3033_index_0_scale_req_1); -- 
    scale_ca_15318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_index_0_scale_ack_1, ack => cp_elements(133)); -- 
    final_index_req_15322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => array_obj_ref_3033_offset_inst_req_0); -- 
    final_index_ack_15323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_offset_inst_ack_0, ack => cp_elements(134)); -- 
    base_resize_ack_15329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_base_resize_ack_0, ack => cp_elements(135)); -- 
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(135));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_15334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => array_obj_ref_3033_root_address_inst_req_0); -- 
    plus_base_ra_15335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_root_address_inst_ack_0, ack => cp_elements(137)); -- 
    plus_base_cr_15336_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(137), ack => array_obj_ref_3033_root_address_inst_req_1); -- 
    plus_base_ca_15337_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_root_address_inst_ack_1, ack => cp_elements(138)); -- 
    final_reg_ack_15342_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3033_final_reg_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(139);
    cp_elements(141) <= cp_elements(140);
    cpelement_group_142 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(159));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(142),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => binary_3047_inst_req_0); -- 
    cp_elements(143) <= cp_elements(141);
    cpelement_group_144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(145) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => type_cast_3046_inst_req_0); -- 
    cp_elements(145) <= cp_elements(141);
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(147) & cp_elements(156));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(146), ack => binary_3045_inst_req_0); -- 
    cp_elements(147) <= cp_elements(141);
    cpelement_group_148 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(148),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => binary_3043_inst_req_0); -- 
    cp_elements(149) <= cp_elements(141);
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(151) & cp_elements(152));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(150), ack => binary_3042_inst_req_0); -- 
    cp_elements(151) <= cp_elements(141);
    cp_elements(152) <= cp_elements(141);
    ra_15366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3042_inst_ack_0, ack => cp_elements(153)); -- 
    cr_15367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => binary_3042_inst_req_1); -- 
    ca_15368_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3042_inst_ack_1, ack => cp_elements(154)); -- 
    ra_15373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3043_inst_ack_0, ack => cp_elements(155)); -- 
    cr_15374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => binary_3043_inst_req_1); -- 
    ca_15375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3043_inst_ack_1, ack => cp_elements(156)); -- 
    ra_15380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3045_inst_ack_0, ack => cp_elements(157)); -- 
    cr_15381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => binary_3045_inst_req_1); -- 
    ca_15382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3045_inst_ack_1, ack => cp_elements(158)); -- 
    ack_15387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3046_inst_ack_0, ack => cp_elements(159)); -- 
    ra_15392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3047_inst_ack_0, ack => cp_elements(160)); -- 
    cr_15393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_3047_inst_req_1); -- 
    ca_15394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3047_inst_ack_1, ack => cp_elements(161)); -- 
    pipe_wreq_15399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => simple_obj_ref_3036_inst_req_0); -- 
    pipe_wack_15400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3036_inst_ack_0, ack => cp_elements(162)); -- 
    cp_elements(163) <= cp_elements(140);
    pipe_wreq_15411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => simple_obj_ref_3049_inst_req_0); -- 
    pipe_wack_15412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3049_inst_ack_0, ack => cp_elements(164)); -- 
    cp_elements(165) <= cp_elements(140);
    pipe_wreq_15422_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => simple_obj_ref_3052_inst_req_0); -- 
    pipe_wack_15423_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3052_inst_ack_0, ack => cp_elements(166)); -- 
    cpelement_group_167 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(162) & cp_elements(164) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(167),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(168) <= cp_elements(69);
    cp_elements(169) <= false;
    cp_elements(170) <= cp_elements(169);
    cp_elements(171) <= cp_elements(69);
    phi_stmt_3002_req_15437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => phi_stmt_3002_req_0); -- 
    cp_elements(172) <= OrReduce(cp_elements(123) & cp_elements(171));
    cp_elements(173) <= cp_elements(172);
    phi_stmt_3002_ack_15452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3002_ack_0, ack => cp_elements(174)); -- 
    cp_elements(175) <= cp_elements(43);
    cp_elements(176) <= false;
    cp_elements(177) <= cp_elements(176);
    cp_elements(178) <= cp_elements(43);
    cp_elements(179) <= OrReduce(cp_elements(47) & cp_elements(178));
    cp_elements(180) <= cp_elements(179);
    cp_elements(181) <= cp_elements(0);
    cp_elements(182) <= false; 
    cp_elements(183) <= OrReduce(cp_elements(262) & cp_elements(265));
    req_15489_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => simple_obj_ref_3062_inst_req_0); -- 
    cp_elements(184) <= cp_elements(259);
    ack_15490_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3062_inst_ack_0, ack => cp_elements(185)); -- 
    cp_elements(186) <= cp_elements(185);
    cp_elements(187) <= cp_elements(186);
    cpelement_group_188 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(187) & cp_elements(216));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(188),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(189) <= cp_elements(187);
    base_resize_req_15509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => ptr_deref_3067_base_resize_req_0); -- 
    base_resize_ack_15510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_base_resize_ack_0, ack => cp_elements(190)); -- 
    sum_rename_req_15514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_3067_root_address_inst_req_0); -- 
    cp_elements(191) <= ptr_deref_3067_root_address_inst_ack_0;
    cp_elements(192) <= cp_elements(191);
    rr_15522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => ptr_deref_3067_addr_0_req_0); -- 
    ra_15523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_0_ack_0, ack => cp_elements(193)); -- 
    cr_15524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => ptr_deref_3067_addr_0_req_1); -- 
    ca_15525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_0_ack_1, ack => cp_elements(194)); -- 
    cp_elements(195) <= cp_elements(191);
    rr_15529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => ptr_deref_3067_addr_1_req_0); -- 
    ra_15530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_1_ack_0, ack => cp_elements(196)); -- 
    cr_15531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => ptr_deref_3067_addr_1_req_1); -- 
    ca_15532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_1_ack_1, ack => cp_elements(197)); -- 
    cp_elements(198) <= cp_elements(191);
    rr_15536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => ptr_deref_3067_addr_2_req_0); -- 
    ra_15537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_2_ack_0, ack => cp_elements(199)); -- 
    cr_15538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => ptr_deref_3067_addr_2_req_1); -- 
    ca_15539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_2_ack_1, ack => cp_elements(200)); -- 
    cp_elements(201) <= cp_elements(191);
    rr_15543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => ptr_deref_3067_addr_3_req_0); -- 
    ra_15544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_3_ack_0, ack => cp_elements(202)); -- 
    cr_15545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(202), ack => ptr_deref_3067_addr_3_req_1); -- 
    ca_15546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_3_ack_1, ack => cp_elements(203)); -- 
    cp_elements(204) <= cp_elements(191);
    rr_15550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_3067_addr_4_req_0); -- 
    ra_15551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_4_ack_0, ack => cp_elements(205)); -- 
    cr_15552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => ptr_deref_3067_addr_4_req_1); -- 
    ca_15553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_4_ack_1, ack => cp_elements(206)); -- 
    cp_elements(207) <= cp_elements(191);
    rr_15557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_3067_addr_5_req_0); -- 
    ra_15558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_5_ack_0, ack => cp_elements(208)); -- 
    cr_15559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => ptr_deref_3067_addr_5_req_1); -- 
    ca_15560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_5_ack_1, ack => cp_elements(209)); -- 
    cp_elements(210) <= cp_elements(191);
    rr_15564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_3067_addr_6_req_0); -- 
    ra_15565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_6_ack_0, ack => cp_elements(211)); -- 
    cr_15566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => ptr_deref_3067_addr_6_req_1); -- 
    ca_15567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_6_ack_1, ack => cp_elements(212)); -- 
    cp_elements(213) <= cp_elements(191);
    rr_15571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_3067_addr_7_req_0); -- 
    ra_15572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_7_ack_0, ack => cp_elements(214)); -- 
    cr_15573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => ptr_deref_3067_addr_7_req_1); -- 
    ca_15574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_addr_7_ack_1, ack => cp_elements(215)); -- 
    cpelement_group_216 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(194) & cp_elements(197) & cp_elements(200) & cp_elements(203) & cp_elements(206) & cp_elements(209) & cp_elements(212) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(216),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(217) <= cp_elements(188);
    rr_15584_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_3067_load_0_req_0); -- 
    ra_15585_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(188);
    rr_15589_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_3067_load_1_req_0); -- 
    ra_15590_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_1_ack_0, ack => cp_elements(220)); -- 
    cp_elements(221) <= cp_elements(188);
    rr_15594_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => ptr_deref_3067_load_2_req_0); -- 
    ra_15595_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_2_ack_0, ack => cp_elements(222)); -- 
    cp_elements(223) <= cp_elements(188);
    rr_15599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => ptr_deref_3067_load_3_req_0); -- 
    ra_15600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_3_ack_0, ack => cp_elements(224)); -- 
    cp_elements(225) <= cp_elements(188);
    rr_15604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => ptr_deref_3067_load_4_req_0); -- 
    ra_15605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_4_ack_0, ack => cp_elements(226)); -- 
    cp_elements(227) <= cp_elements(188);
    rr_15609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => ptr_deref_3067_load_5_req_0); -- 
    ra_15610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_5_ack_0, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(188);
    rr_15614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => ptr_deref_3067_load_6_req_0); -- 
    ra_15615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_6_ack_0, ack => cp_elements(230)); -- 
    cp_elements(231) <= cp_elements(188);
    rr_15619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_3067_load_7_req_0); -- 
    ra_15620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_7_ack_0, ack => cp_elements(232)); -- 
    cpelement_group_233 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220) & cp_elements(222) & cp_elements(224) & cp_elements(226) & cp_elements(228) & cp_elements(230) & cp_elements(232));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(233),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(234) <= cp_elements(233);
    cr_15630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_3067_load_0_req_1); -- 
    ca_15631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_0_ack_1, ack => cp_elements(235)); -- 
    cp_elements(236) <= cp_elements(233);
    cr_15635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_3067_load_1_req_1); -- 
    ca_15636_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_1_ack_1, ack => cp_elements(237)); -- 
    cp_elements(238) <= cp_elements(233);
    cr_15640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => ptr_deref_3067_load_2_req_1); -- 
    ca_15641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_2_ack_1, ack => cp_elements(239)); -- 
    cp_elements(240) <= cp_elements(233);
    cr_15645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_3067_load_3_req_1); -- 
    ca_15646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_3_ack_1, ack => cp_elements(241)); -- 
    cp_elements(242) <= cp_elements(233);
    cr_15650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => ptr_deref_3067_load_4_req_1); -- 
    ca_15651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_4_ack_1, ack => cp_elements(243)); -- 
    cp_elements(244) <= cp_elements(233);
    cr_15655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_3067_load_5_req_1); -- 
    ca_15656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_5_ack_1, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(233);
    cr_15660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_3067_load_6_req_1); -- 
    ca_15661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_6_ack_1, ack => cp_elements(247)); -- 
    cp_elements(248) <= cp_elements(233);
    cr_15665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => ptr_deref_3067_load_7_req_1); -- 
    ca_15666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_load_7_ack_1, ack => cp_elements(249)); -- 
    cpelement_group_250 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(235) & cp_elements(237) & cp_elements(239) & cp_elements(241) & cp_elements(243) & cp_elements(245) & cp_elements(247) & cp_elements(249));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(250),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_15667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_3067_gather_scatter_req_0); -- 
    merge_ack_15668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3067_gather_scatter_ack_0, ack => cp_elements(251)); -- 
    pipe_wreq_15673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => simple_obj_ref_3065_inst_req_0); -- 
    pipe_wack_15674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3065_inst_ack_0, ack => cp_elements(252)); -- 
    cp_elements(253) <= cp_elements(186);
    req_15684_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(253), ack => simple_obj_ref_3070_inst_req_0); -- 
    ack_15685_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3070_inst_ack_0, ack => cp_elements(254)); -- 
    pipe_wreq_15690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(254), ack => simple_obj_ref_3069_inst_req_0); -- 
    pipe_wack_15691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3069_inst_ack_0, ack => cp_elements(255)); -- 
    cp_elements(256) <= cp_elements(186);
    req_15701_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => simple_obj_ref_3073_inst_req_0); -- 
    ack_15702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3073_inst_ack_0, ack => cp_elements(257)); -- 
    pipe_wreq_15707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => simple_obj_ref_3072_inst_req_0); -- 
    pipe_wack_15708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3072_inst_ack_0, ack => cp_elements(258)); -- 
    cpelement_group_259 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(252) & cp_elements(255) & cp_elements(258));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(260) <= cp_elements(181);
    cp_elements(261) <= false;
    cp_elements(262) <= cp_elements(261);
    cp_elements(263) <= cp_elements(181);
    cp_elements(264) <= OrReduce(cp_elements(184) & cp_elements(263));
    cp_elements(265) <= cp_elements(264);
    cp_elements(266) <= cp_elements(0);
    cp_elements(267) <= false; 
    cp_elements(268) <= OrReduce(cp_elements(384) & cp_elements(387));
    req_15747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => simple_obj_ref_3081_inst_req_0); -- 
    cp_elements(269) <= cp_elements(366);
    cp_elements(270) <= OrReduce(cp_elements(369) & cp_elements(378) & cp_elements(381));
    ack_15748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3081_inst_ack_0, ack => cp_elements(271)); -- 
    cp_elements(272) <= cp_elements(271);
    cp_elements(273) <= cp_elements(272);
    cpelement_group_274 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(275) & cp_elements(315) & cp_elements(359));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(274),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => binary_3121_inst_req_0); -- 
    cp_elements(275) <= cp_elements(273);
    cpelement_group_276 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(277) & cp_elements(293) & cp_elements(313));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(276),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(276), ack => binary_3101_inst_req_0); -- 
    cp_elements(277) <= cp_elements(273);
    cpelement_group_278 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(279) & cp_elements(283) & cp_elements(291));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(278),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(278), ack => binary_3091_inst_req_0); -- 
    cp_elements(279) <= cp_elements(273);
    cpelement_group_280 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(281) & cp_elements(282));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(280),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(280), ack => type_cast_3086_inst_req_0); -- 
    cp_elements(281) <= cp_elements(273);
    cp_elements(282) <= cp_elements(273);
    ack_15770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3086_inst_ack_0, ack => cp_elements(283)); -- 
    cpelement_group_284 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(285) & cp_elements(290));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(284),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => type_cast_3090_inst_req_0); -- 
    cp_elements(285) <= cp_elements(273);
    cpelement_group_286 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(287) & cp_elements(288));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(286),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => binary_3089_inst_req_0); -- 
    cp_elements(287) <= cp_elements(273);
    cp_elements(288) <= cp_elements(273);
    ra_15780_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3089_inst_ack_0, ack => cp_elements(289)); -- 
    cr_15781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(289), ack => binary_3089_inst_req_1); -- 
    ca_15782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3089_inst_ack_1, ack => cp_elements(290)); -- 
    ack_15787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3090_inst_ack_0, ack => cp_elements(291)); -- 
    ra_15792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3091_inst_ack_0, ack => cp_elements(292)); -- 
    cr_15793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => binary_3091_inst_req_1); -- 
    ca_15794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3091_inst_ack_1, ack => cp_elements(293)); -- 
    cpelement_group_294 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(295) & cp_elements(303) & cp_elements(311));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(294),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(294), ack => binary_3100_inst_req_0); -- 
    cp_elements(295) <= cp_elements(273);
    cpelement_group_296 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(297) & cp_elements(302));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(296),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(296), ack => type_cast_3095_inst_req_0); -- 
    cp_elements(297) <= cp_elements(273);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => binary_3094_inst_req_0); -- 
    cp_elements(299) <= cp_elements(273);
    cp_elements(300) <= cp_elements(273);
    ra_15806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3094_inst_ack_0, ack => cp_elements(301)); -- 
    cr_15807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => binary_3094_inst_req_1); -- 
    ca_15808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3094_inst_ack_1, ack => cp_elements(302)); -- 
    ack_15813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3095_inst_ack_0, ack => cp_elements(303)); -- 
    cpelement_group_304 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(305) & cp_elements(310));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(304),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(304), ack => type_cast_3099_inst_req_0); -- 
    cp_elements(305) <= cp_elements(273);
    cpelement_group_306 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(307) & cp_elements(308));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(306),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(306), ack => binary_3098_inst_req_0); -- 
    cp_elements(307) <= cp_elements(273);
    cp_elements(308) <= cp_elements(273);
    ra_15823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3098_inst_ack_0, ack => cp_elements(309)); -- 
    cr_15824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(309), ack => binary_3098_inst_req_1); -- 
    ca_15825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3098_inst_ack_1, ack => cp_elements(310)); -- 
    ack_15830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3099_inst_ack_0, ack => cp_elements(311)); -- 
    ra_15835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3100_inst_ack_0, ack => cp_elements(312)); -- 
    cr_15836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(312), ack => binary_3100_inst_req_1); -- 
    ca_15837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3100_inst_ack_1, ack => cp_elements(313)); -- 
    ra_15842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3101_inst_ack_0, ack => cp_elements(314)); -- 
    cr_15843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(314), ack => binary_3101_inst_req_1); -- 
    ca_15844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3101_inst_ack_1, ack => cp_elements(315)); -- 
    cpelement_group_316 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(317) & cp_elements(337) & cp_elements(357));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(316),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => binary_3120_inst_req_0); -- 
    cp_elements(317) <= cp_elements(273);
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(319) & cp_elements(327) & cp_elements(335));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => binary_3110_inst_req_0); -- 
    cp_elements(319) <= cp_elements(273);
    cpelement_group_320 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(321) & cp_elements(326));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(320),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(320), ack => type_cast_3105_inst_req_0); -- 
    cp_elements(321) <= cp_elements(273);
    cpelement_group_322 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(323) & cp_elements(324));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(322),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(322), ack => binary_3104_inst_req_0); -- 
    cp_elements(323) <= cp_elements(273);
    cp_elements(324) <= cp_elements(273);
    ra_15858_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3104_inst_ack_0, ack => cp_elements(325)); -- 
    cr_15859_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => binary_3104_inst_req_1); -- 
    ca_15860_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3104_inst_ack_1, ack => cp_elements(326)); -- 
    ack_15865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3105_inst_ack_0, ack => cp_elements(327)); -- 
    cpelement_group_328 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(329) & cp_elements(334));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => type_cast_3109_inst_req_0); -- 
    cp_elements(329) <= cp_elements(273);
    cpelement_group_330 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(331) & cp_elements(332));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(330),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => binary_3108_inst_req_0); -- 
    cp_elements(331) <= cp_elements(273);
    cp_elements(332) <= cp_elements(273);
    ra_15875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3108_inst_ack_0, ack => cp_elements(333)); -- 
    cr_15876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => binary_3108_inst_req_1); -- 
    ca_15877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3108_inst_ack_1, ack => cp_elements(334)); -- 
    ack_15882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3109_inst_ack_0, ack => cp_elements(335)); -- 
    ra_15887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3110_inst_ack_0, ack => cp_elements(336)); -- 
    cr_15888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => binary_3110_inst_req_1); -- 
    ca_15889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3110_inst_ack_1, ack => cp_elements(337)); -- 
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(339) & cp_elements(347) & cp_elements(355));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => binary_3119_inst_req_0); -- 
    cp_elements(339) <= cp_elements(273);
    cpelement_group_340 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(341) & cp_elements(346));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(340),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => type_cast_3114_inst_req_0); -- 
    cp_elements(341) <= cp_elements(273);
    cpelement_group_342 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(343) & cp_elements(344));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(342),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15900_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(342), ack => binary_3113_inst_req_0); -- 
    cp_elements(343) <= cp_elements(273);
    cp_elements(344) <= cp_elements(273);
    ra_15901_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3113_inst_ack_0, ack => cp_elements(345)); -- 
    cr_15902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => binary_3113_inst_req_1); -- 
    ca_15903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3113_inst_ack_1, ack => cp_elements(346)); -- 
    ack_15908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3114_inst_ack_0, ack => cp_elements(347)); -- 
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(349) & cp_elements(354));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => type_cast_3118_inst_req_0); -- 
    cp_elements(349) <= cp_elements(273);
    cpelement_group_350 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(351) & cp_elements(352));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(350),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => binary_3117_inst_req_0); -- 
    cp_elements(351) <= cp_elements(273);
    cp_elements(352) <= cp_elements(273);
    ra_15918_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3117_inst_ack_0, ack => cp_elements(353)); -- 
    cr_15919_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => binary_3117_inst_req_1); -- 
    ca_15920_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3117_inst_ack_1, ack => cp_elements(354)); -- 
    ack_15925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3118_inst_ack_0, ack => cp_elements(355)); -- 
    ra_15930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3119_inst_ack_0, ack => cp_elements(356)); -- 
    cr_15931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => binary_3119_inst_req_1); -- 
    ca_15932_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3119_inst_ack_1, ack => cp_elements(357)); -- 
    ra_15937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3120_inst_ack_0, ack => cp_elements(358)); -- 
    cr_15938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(358), ack => binary_3120_inst_req_1); -- 
    ca_15939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3120_inst_ack_1, ack => cp_elements(359)); -- 
    ra_15944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3121_inst_ack_0, ack => cp_elements(360)); -- 
    cr_15945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => binary_3121_inst_req_1); -- 
    ca_15946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3121_inst_ack_1, ack => cp_elements(361)); -- 
    pipe_wreq_15951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(361), ack => simple_obj_ref_3084_inst_req_0); -- 
    pipe_wack_15952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3084_inst_ack_0, ack => cp_elements(362)); -- 
    cp_elements(363) <= cp_elements(272);
    req_15962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(363), ack => simple_obj_ref_3124_inst_req_0); -- 
    ack_15963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3124_inst_ack_0, ack => cp_elements(364)); -- 
    pipe_wreq_15968_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(364), ack => simple_obj_ref_3123_inst_req_0); -- 
    pipe_wack_15969_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3123_inst_ack_0, ack => cp_elements(365)); -- 
    cpelement_group_366 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(362) & cp_elements(365));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(366),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(367) <= cp_elements(269);
    cp_elements(368) <= false;
    cp_elements(369) <= cp_elements(368);
    cp_elements(370) <= cp_elements(269);
    req_15986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(370), ack => simple_obj_ref_3128_inst_req_0); -- 
    ack_15987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3128_inst_ack_0, ack => cp_elements(371)); -- 
    rr_15988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => binary_3130_inst_req_0); -- 
    ra_15989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3130_inst_ack_0, ack => cp_elements(372)); -- 
    cr_15990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(372), ack => binary_3130_inst_req_1); -- 
    ca_15991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3130_inst_ack_1, ack => cp_elements(373)); -- 
    branch_req_15992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(373), ack => if_stmt_3127_branch_req_0); -- 
    cp_elements(374) <= cp_elements(373);
    cp_elements(375) <= cp_elements(374);
    if_choice_transition_15997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3127_branch_ack_1, ack => cp_elements(376)); -- 
    req_16011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(376), ack => simple_obj_ref_3131_inst_req_0); -- 
    cp_elements(377) <= cp_elements(374);
    else_choice_transition_16001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3127_branch_ack_0, ack => cp_elements(378)); -- 
    ack_16012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3131_inst_ack_0, ack => cp_elements(379)); -- 
    crr_16018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(379), ack => call_stmt_3132_call_req_0); -- 
    cra_16019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3132_call_ack_0, ack => cp_elements(380)); -- 
    ccr_16023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => call_stmt_3132_call_req_1); -- 
    cca_16024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3132_call_ack_1, ack => cp_elements(381)); -- 
    cp_elements(382) <= cp_elements(266);
    cp_elements(383) <= false;
    cp_elements(384) <= cp_elements(383);
    cp_elements(385) <= cp_elements(266);
    cp_elements(386) <= OrReduce(cp_elements(270) & cp_elements(385));
    cp_elements(387) <= cp_elements(386);
    cpelement_group_388 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(44) & cp_elements(182) & cp_elements(267));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(388),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_3002 : std_logic_vector(15 downto 0);
    signal LI_2999 : std_logic_vector(15 downto 0);
    signal NI_3023 : std_logic_vector(15 downto 0);
    signal a_3082 : std_logic_vector(63 downto 0);
    signal array_obj_ref_3014_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3014_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_3014_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3014_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3014_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_3033_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3033_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_3033_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3033_root_address : std_logic_vector(15 downto 0);
    signal binary_2984_wire : std_logic_vector(0 downto 0);
    signal binary_3028_wire : std_logic_vector(0 downto 0);
    signal binary_3042_wire : std_logic_vector(15 downto 0);
    signal binary_3043_wire : std_logic_vector(15 downto 0);
    signal binary_3045_wire : std_logic_vector(15 downto 0);
    signal binary_3047_wire : std_logic_vector(7 downto 0);
    signal binary_3089_wire : std_logic_vector(63 downto 0);
    signal binary_3091_wire : std_logic_vector(15 downto 0);
    signal binary_3094_wire : std_logic_vector(63 downto 0);
    signal binary_3098_wire : std_logic_vector(63 downto 0);
    signal binary_3100_wire : std_logic_vector(15 downto 0);
    signal binary_3101_wire : std_logic_vector(31 downto 0);
    signal binary_3104_wire : std_logic_vector(63 downto 0);
    signal binary_3108_wire : std_logic_vector(63 downto 0);
    signal binary_3110_wire : std_logic_vector(15 downto 0);
    signal binary_3113_wire : std_logic_vector(63 downto 0);
    signal binary_3117_wire : std_logic_vector(63 downto 0);
    signal binary_3119_wire : std_logic_vector(15 downto 0);
    signal binary_3120_wire : std_logic_vector(31 downto 0);
    signal binary_3121_wire : std_logic_vector(63 downto 0);
    signal binary_3130_wire : std_logic_vector(0 downto 0);
    signal blen_2942 : std_logic_vector(15 downto 0);
    signal blen_2973 : std_logic_vector(15 downto 0);
    signal buf64_2976 : std_logic_vector(31 downto 0);
    signal buf_2942 : std_logic_vector(31 downto 0);
    signal expr_2983_wire_constant : std_logic_vector(15 downto 0);
    signal expr_2987_wire_constant : std_logic_vector(7 downto 0);
    signal expr_2993_wire_constant : std_logic_vector(0 downto 0);
    signal expr_2997_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3010_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3017_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3021_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3039_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3041_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3044_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3053_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3088_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3093_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3097_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3103_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3107_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3112_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3116_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3129_wire_constant : std_logic_vector(0 downto 0);
    signal last_word_ptr_3034 : std_logic_vector(31 downto 0);
    signal pkt64_2979 : std_logic_vector(31 downto 0);
    signal pkt_2936 : std_logic_vector(31 downto 0);
    signal ptr_3063 : std_logic_vector(31 downto 0);
    signal ptr_deref_3067_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_4 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_5 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_6 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_data_7 : std_logic_vector(7 downto 0);
    signal ptr_deref_3067_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3067_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_address_7 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_3067_word_offset_7 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3013_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3013_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3032_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3032_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3070_wire : std_logic_vector(7 downto 0);
    signal simple_obj_ref_3073_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3124_wire : std_logic_vector(7 downto 0);
    signal simple_obj_ref_3128_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3131_wire : std_logic_vector(31 downto 0);
    signal type_cast_2938_wire : std_logic_vector(31 downto 0);
    signal type_cast_2946_wire : std_logic_vector(31 downto 0);
    signal type_cast_2950_wire : std_logic_vector(31 downto 0);
    signal type_cast_2960_wire : std_logic_vector(31 downto 0);
    signal type_cast_3005_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3038_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3046_wire : std_logic_vector(7 downto 0);
    signal type_cast_3086_wire : std_logic_vector(7 downto 0);
    signal type_cast_3090_wire : std_logic_vector(7 downto 0);
    signal type_cast_3095_wire : std_logic_vector(7 downto 0);
    signal type_cast_3099_wire : std_logic_vector(7 downto 0);
    signal type_cast_3105_wire : std_logic_vector(7 downto 0);
    signal type_cast_3109_wire : std_logic_vector(7 downto 0);
    signal type_cast_3114_wire : std_logic_vector(7 downto 0);
    signal type_cast_3118_wire : std_logic_vector(7 downto 0);
    signal wlen_2942 : std_logic_vector(15 downto 0);
    signal wlen_2970 : std_logic_vector(15 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxblen_pipe
    signal xxsend_packet_pipelinexxblen_pipe_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxblen_pipe
    signal xxsend_packet_pipelinexxblen_pipe_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxbuf64_pipe
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxbuf64_pipe
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxpkt64_pipe
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxpkt64_pipe
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxread_ctrl_in
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxread_ctrl_in
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxread_last_word_in
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxread_last_word_in
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxread_pointer
    signal xxsend_packet_pipelinexxread_pointer_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxread_pointer
    signal xxsend_packet_pipelinexxread_pointer_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxswap_ctrl_in
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxswap_ctrl_in
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxswap_data_in
    signal xxsend_packet_pipelinexxswap_data_in_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxswap_data_in
    signal xxsend_packet_pipelinexxswap_data_in_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxswap_last_word_in
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxswap_last_word_in
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxwlen_pipe
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxwlen_pipe
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_3014_offset_scale_factor_0 <= "0000000000001000";
    array_obj_ref_3033_offset_scale_factor_0 <= "0000000000001000";
    expr_2983_wire_constant <= "0000000000000000";
    expr_2987_wire_constant <= "11111111";
    expr_2993_wire_constant <= "0";
    expr_2997_wire_constant <= "0000000000000001";
    expr_3010_wire_constant <= "00000000";
    expr_3017_wire_constant <= "0";
    expr_3021_wire_constant <= "0000000000000001";
    expr_3039_wire_constant <= "0000000000001000";
    expr_3041_wire_constant <= "0000000000000111";
    expr_3044_wire_constant <= "0000000000000111";
    expr_3053_wire_constant <= "1";
    expr_3088_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    expr_3093_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    expr_3097_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    expr_3103_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    expr_3107_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    expr_3112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    expr_3116_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    expr_3129_wire_constant <= "0";
    ptr_deref_3067_word_offset_0 <= "0000000000000000";
    ptr_deref_3067_word_offset_1 <= "0000000000000001";
    ptr_deref_3067_word_offset_2 <= "0000000000000010";
    ptr_deref_3067_word_offset_3 <= "0000000000000011";
    ptr_deref_3067_word_offset_4 <= "0000000000000100";
    ptr_deref_3067_word_offset_5 <= "0000000000000101";
    ptr_deref_3067_word_offset_6 <= "0000000000000110";
    ptr_deref_3067_word_offset_7 <= "0000000000000111";
    type_cast_3005_wire_constant <= "0000000000000000";
    type_cast_3038_wire_constant <= "00000001";
    phi_stmt_3002: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3005_wire_constant & NI_3023;
      req <= phi_stmt_3002_req_0 & phi_stmt_3002_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3002_ack_0,
          idata => idata,
          odata => I_3002,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3002
    array_obj_ref_3014_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => pkt64_2979, dout => array_obj_ref_3014_resized_base_address, req => array_obj_ref_3014_base_resize_req_0, ack => array_obj_ref_3014_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3014_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3014_root_address, dout => array_obj_ref_3014_wire, req => array_obj_ref_3014_final_reg_req_0, ack => array_obj_ref_3014_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3014_index_0_resize: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => I_3002, dout => simple_obj_ref_3013_resized, req => array_obj_ref_3014_index_0_resize_req_0, ack => array_obj_ref_3014_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3014_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3013_scaled, dout => array_obj_ref_3014_final_offset, req => array_obj_ref_3014_offset_inst_req_0, ack => array_obj_ref_3014_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3033_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => pkt64_2979, dout => array_obj_ref_3033_resized_base_address, req => array_obj_ref_3033_base_resize_req_0, ack => array_obj_ref_3033_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3033_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3033_root_address, dout => last_word_ptr_3034, req => array_obj_ref_3033_final_reg_req_0, ack => array_obj_ref_3033_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3033_index_0_resize: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => LI_2999, dout => simple_obj_ref_3032_resized, req => array_obj_ref_3033_index_0_resize_req_0, ack => array_obj_ref_3033_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3033_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3032_scaled, dout => array_obj_ref_3033_final_offset, req => array_obj_ref_3033_offset_inst_req_0, ack => array_obj_ref_3033_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3067_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => ptr_3063, dout => ptr_deref_3067_resized_base_address, req => ptr_deref_3067_base_resize_req_0, ack => ptr_deref_3067_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2938_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt_2936, dout => type_cast_2938_wire, req => type_cast_2938_inst_req_0, ack => type_cast_2938_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2946_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => buf_2942, dout => type_cast_2946_wire, req => type_cast_2946_inst_req_0, ack => type_cast_2946_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2950_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt_2936, dout => type_cast_2950_wire, req => type_cast_2950_inst_req_0, ack => type_cast_2950_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2960_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt_2936, dout => type_cast_2960_wire, req => type_cast_2960_inst_req_0, ack => type_cast_2960_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3046_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3045_wire, dout => type_cast_3046_wire, req => type_cast_3046_inst_req_0, ack => type_cast_3046_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3086_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => a_3082, dout => type_cast_3086_wire, req => type_cast_3086_inst_req_0, ack => type_cast_3086_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3090_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3089_wire, dout => type_cast_3090_wire, req => type_cast_3090_inst_req_0, ack => type_cast_3090_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3095_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3094_wire, dout => type_cast_3095_wire, req => type_cast_3095_inst_req_0, ack => type_cast_3095_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3099_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3098_wire, dout => type_cast_3099_wire, req => type_cast_3099_inst_req_0, ack => type_cast_3099_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3105_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3104_wire, dout => type_cast_3105_wire, req => type_cast_3105_inst_req_0, ack => type_cast_3105_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3109_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3108_wire, dout => type_cast_3109_wire, req => type_cast_3109_inst_req_0, ack => type_cast_3109_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3114_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3113_wire, dout => type_cast_3114_wire, req => type_cast_3114_inst_req_0, ack => type_cast_3114_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3118_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3117_wire, dout => type_cast_3118_wire, req => type_cast_3118_inst_req_0, ack => type_cast_3118_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3067_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(63 downto 0); --
    begin -- 
      ptr_deref_3067_gather_scatter_ack_0 <= ptr_deref_3067_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3067_data_7 & ptr_deref_3067_data_6 & ptr_deref_3067_data_5 & ptr_deref_3067_data_4 & ptr_deref_3067_data_3 & ptr_deref_3067_data_2 & ptr_deref_3067_data_1 & ptr_deref_3067_data_0;
      ptr_deref_3067_wire <= aggregated_sig(63 downto 0);
      --
    end Block;
    ptr_deref_3067_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3067_root_address_inst_ack_0 <= ptr_deref_3067_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3067_resized_base_address;
      ptr_deref_3067_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_2981_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_2984_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2981_branch_req_0,
          ack0 => if_stmt_2981_branch_ack_0,
          ack1 => if_stmt_2981_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3025_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3028_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3025_branch_req_0,
          ack0 => if_stmt_3025_branch_ack_0,
          ack1 => if_stmt_3025_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3127_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3130_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3127_branch_req_0,
          ack0 => if_stmt_3127_branch_ack_0,
          ack1 => if_stmt_3127_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_3014_index_0_scale array_obj_ref_3033_index_0_scale 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3013_resized & simple_obj_ref_3032_resized;
      simple_obj_ref_3013_scaled <= data_out(31 downto 16);
      simple_obj_ref_3032_scaled <= data_out(15 downto 0);
      reqL(1) <= array_obj_ref_3014_index_0_scale_req_0;
      reqL(0) <= array_obj_ref_3033_index_0_scale_req_0;
      array_obj_ref_3014_index_0_scale_ack_0 <= ackL(1);
      array_obj_ref_3033_index_0_scale_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_3014_index_0_scale_req_1;
      reqR(0) <= array_obj_ref_3033_index_0_scale_req_1;
      array_obj_ref_3014_index_0_scale_ack_1 <= ackR(1);
      array_obj_ref_3033_index_0_scale_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_3014_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3014_final_offset & array_obj_ref_3014_resized_base_address;
      array_obj_ref_3014_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3014_root_address_inst_req_0,
          ackL => array_obj_ref_3014_root_address_inst_ack_0,
          reqR => array_obj_ref_3014_root_address_inst_req_1,
          ackR => array_obj_ref_3014_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_3033_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3033_final_offset & array_obj_ref_3033_resized_base_address;
      array_obj_ref_3033_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3033_root_address_inst_req_0,
          ackL => array_obj_ref_3033_root_address_inst_ack_0,
          reqR => array_obj_ref_3033_root_address_inst_req_1,
          ackR => array_obj_ref_3033_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2984_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= wlen_2970;
      binary_2984_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2984_inst_req_0,
          ackL => binary_2984_inst_ack_0,
          reqR => binary_2984_inst_req_1,
          ackR => binary_2984_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2998_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= wlen_2970;
      LI_2999 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2998_inst_req_0,
          ackL => binary_2998_inst_ack_0,
          reqR => binary_2998_inst_req_1,
          ackR => binary_2998_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_3022_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_3002;
      NI_3023 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3022_inst_req_0,
          ackL => binary_3022_inst_ack_0,
          reqR => binary_3022_inst_req_1,
          ackR => binary_3022_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_3028_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= NI_3023 & LI_2999;
      binary_3028_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3028_inst_req_0,
          ackL => binary_3028_inst_ack_0,
          reqR => binary_3028_inst_req_1,
          ackR => binary_3028_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_3042_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= blen_2973;
      binary_3042_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3042_inst_req_0,
          ackL => binary_3042_inst_ack_0,
          reqR => binary_3042_inst_req_1,
          ackR => binary_3042_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_3043_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= expr_3039_wire_constant & binary_3042_wire;
      binary_3043_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3043_inst_req_0,
          ackL => binary_3043_inst_ack_0,
          reqR => binary_3043_inst_req_1,
          ackR => binary_3043_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_3045_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3043_wire;
      binary_3045_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3045_inst_req_0,
          ackL => binary_3045_inst_ack_0,
          reqR => binary_3045_inst_req_1,
          ackR => binary_3045_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_3047_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3038_wire_constant & type_cast_3046_wire;
      binary_3047_wire <= data_out(7 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3047_inst_req_0,
          ackL => binary_3047_inst_ack_0,
          reqR => binary_3047_inst_req_1,
          ackR => binary_3047_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_3089_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3089_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3089_inst_req_0,
          ackL => binary_3089_inst_ack_0,
          reqR => binary_3089_inst_req_1,
          ackR => binary_3089_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_3091_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3086_wire & type_cast_3090_wire;
      binary_3091_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3091_inst_req_0,
          ackL => binary_3091_inst_ack_0,
          reqR => binary_3091_inst_req_1,
          ackR => binary_3091_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_3094_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3094_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3094_inst_req_0,
          ackL => binary_3094_inst_ack_0,
          reqR => binary_3094_inst_req_1,
          ackR => binary_3094_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_3098_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3098_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3098_inst_req_0,
          ackL => binary_3098_inst_ack_0,
          reqR => binary_3098_inst_req_1,
          ackR => binary_3098_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_3100_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3095_wire & type_cast_3099_wire;
      binary_3100_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3100_inst_req_0,
          ackL => binary_3100_inst_ack_0,
          reqR => binary_3100_inst_req_1,
          ackR => binary_3100_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_3101_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3091_wire & binary_3100_wire;
      binary_3101_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3101_inst_req_0,
          ackL => binary_3101_inst_ack_0,
          reqR => binary_3101_inst_req_1,
          ackR => binary_3101_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_3104_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3104_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3104_inst_req_0,
          ackL => binary_3104_inst_ack_0,
          reqR => binary_3104_inst_req_1,
          ackR => binary_3104_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_3108_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3108_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3108_inst_req_0,
          ackL => binary_3108_inst_ack_0,
          reqR => binary_3108_inst_req_1,
          ackR => binary_3108_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_3110_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3105_wire & type_cast_3109_wire;
      binary_3110_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3110_inst_req_0,
          ackL => binary_3110_inst_ack_0,
          reqR => binary_3110_inst_req_1,
          ackR => binary_3110_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_3113_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3113_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3113_inst_req_0,
          ackL => binary_3113_inst_ack_0,
          reqR => binary_3113_inst_req_1,
          ackR => binary_3113_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_3117_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3082;
      binary_3117_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3117_inst_req_0,
          ackL => binary_3117_inst_ack_0,
          reqR => binary_3117_inst_req_1,
          ackR => binary_3117_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_3119_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3114_wire & type_cast_3118_wire;
      binary_3119_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3119_inst_req_0,
          ackL => binary_3119_inst_ack_0,
          reqR => binary_3119_inst_req_1,
          ackR => binary_3119_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_3120_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3110_wire & binary_3119_wire;
      binary_3120_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3120_inst_req_0,
          ackL => binary_3120_inst_ack_0,
          reqR => binary_3120_inst_req_1,
          ackR => binary_3120_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_3121_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3101_wire & binary_3120_wire;
      binary_3121_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3121_inst_req_0,
          ackL => binary_3121_inst_ack_0,
          reqR => binary_3121_inst_req_1,
          ackR => binary_3121_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_3130_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3128_wire;
      binary_3130_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3130_inst_req_0,
          ackL => binary_3130_inst_ack_0,
          reqR => binary_3130_inst_req_1,
          ackR => binary_3130_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_3067_addr_0 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_0_req_0,
          ackL => ptr_deref_3067_addr_0_ack_0,
          reqR => ptr_deref_3067_addr_0_req_1,
          ackR => ptr_deref_3067_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_3067_addr_1 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_1_req_0,
          ackL => ptr_deref_3067_addr_1_ack_0,
          reqR => ptr_deref_3067_addr_1_req_1,
          ackR => ptr_deref_3067_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_3067_addr_2 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_2_req_0,
          ackL => ptr_deref_3067_addr_2_ack_0,
          reqR => ptr_deref_3067_addr_2_req_1,
          ackR => ptr_deref_3067_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : ptr_deref_3067_addr_3 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_3_req_0,
          ackL => ptr_deref_3067_addr_3_ack_0,
          reqR => ptr_deref_3067_addr_3_req_1,
          ackR => ptr_deref_3067_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : ptr_deref_3067_addr_4 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_4 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_4_req_0,
          ackL => ptr_deref_3067_addr_4_ack_0,
          reqR => ptr_deref_3067_addr_4_req_1,
          ackR => ptr_deref_3067_addr_4_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : ptr_deref_3067_addr_5 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_5 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000101",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_5_req_0,
          ackL => ptr_deref_3067_addr_5_ack_0,
          reqR => ptr_deref_3067_addr_5_req_1,
          ackR => ptr_deref_3067_addr_5_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : ptr_deref_3067_addr_6 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_6 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_6_req_0,
          ackL => ptr_deref_3067_addr_6_ack_0,
          reqR => ptr_deref_3067_addr_6_req_1,
          ackR => ptr_deref_3067_addr_6_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : ptr_deref_3067_addr_7 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3067_root_address;
      ptr_deref_3067_word_address_7 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3067_addr_7_req_0,
          ackL => ptr_deref_3067_addr_7_ack_0,
          reqR => ptr_deref_3067_addr_7_req_1,
          ackR => ptr_deref_3067_addr_7_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared load operator group (0) : ptr_deref_3067_load_1 ptr_deref_3067_load_5 ptr_deref_3067_load_3 ptr_deref_3067_load_2 ptr_deref_3067_load_6 ptr_deref_3067_load_7 ptr_deref_3067_load_0 ptr_deref_3067_load_4 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3067_load_1_req_0,
        ptr_deref_3067_load_1_ack_0,
        ptr_deref_3067_load_1_req_1,
        ptr_deref_3067_load_1_ack_1,
        "ptr_deref_3067_load_1",
        "memory_space_5" ,
        ptr_deref_3067_data_1,
        ptr_deref_3067_word_address_1,
        "ptr_deref_3067_data_1",
        "ptr_deref_3067_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_5_req_0,
        ptr_deref_3067_load_5_ack_0,
        ptr_deref_3067_load_5_req_1,
        ptr_deref_3067_load_5_ack_1,
        "ptr_deref_3067_load_5",
        "memory_space_5" ,
        ptr_deref_3067_data_5,
        ptr_deref_3067_word_address_5,
        "ptr_deref_3067_data_5",
        "ptr_deref_3067_word_address_5" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_3_req_0,
        ptr_deref_3067_load_3_ack_0,
        ptr_deref_3067_load_3_req_1,
        ptr_deref_3067_load_3_ack_1,
        "ptr_deref_3067_load_3",
        "memory_space_5" ,
        ptr_deref_3067_data_3,
        ptr_deref_3067_word_address_3,
        "ptr_deref_3067_data_3",
        "ptr_deref_3067_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_2_req_0,
        ptr_deref_3067_load_2_ack_0,
        ptr_deref_3067_load_2_req_1,
        ptr_deref_3067_load_2_ack_1,
        "ptr_deref_3067_load_2",
        "memory_space_5" ,
        ptr_deref_3067_data_2,
        ptr_deref_3067_word_address_2,
        "ptr_deref_3067_data_2",
        "ptr_deref_3067_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_6_req_0,
        ptr_deref_3067_load_6_ack_0,
        ptr_deref_3067_load_6_req_1,
        ptr_deref_3067_load_6_ack_1,
        "ptr_deref_3067_load_6",
        "memory_space_5" ,
        ptr_deref_3067_data_6,
        ptr_deref_3067_word_address_6,
        "ptr_deref_3067_data_6",
        "ptr_deref_3067_word_address_6" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_7_req_0,
        ptr_deref_3067_load_7_ack_0,
        ptr_deref_3067_load_7_req_1,
        ptr_deref_3067_load_7_ack_1,
        "ptr_deref_3067_load_7",
        "memory_space_5" ,
        ptr_deref_3067_data_7,
        ptr_deref_3067_word_address_7,
        "ptr_deref_3067_data_7",
        "ptr_deref_3067_word_address_7" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_0_req_0,
        ptr_deref_3067_load_0_ack_0,
        ptr_deref_3067_load_0_req_1,
        ptr_deref_3067_load_0_ack_1,
        "ptr_deref_3067_load_0",
        "memory_space_5" ,
        ptr_deref_3067_data_0,
        ptr_deref_3067_word_address_0,
        "ptr_deref_3067_data_0",
        "ptr_deref_3067_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3067_load_4_req_0,
        ptr_deref_3067_load_4_ack_0,
        ptr_deref_3067_load_4_req_1,
        ptr_deref_3067_load_4_ack_1,
        "ptr_deref_3067_load_4",
        "memory_space_5" ,
        ptr_deref_3067_data_4,
        ptr_deref_3067_word_address_4,
        "ptr_deref_3067_data_4",
        "ptr_deref_3067_word_address_4" -- 
      );
      reqL(7) <= ptr_deref_3067_load_1_req_0;
      reqL(6) <= ptr_deref_3067_load_5_req_0;
      reqL(5) <= ptr_deref_3067_load_3_req_0;
      reqL(4) <= ptr_deref_3067_load_2_req_0;
      reqL(3) <= ptr_deref_3067_load_6_req_0;
      reqL(2) <= ptr_deref_3067_load_7_req_0;
      reqL(1) <= ptr_deref_3067_load_0_req_0;
      reqL(0) <= ptr_deref_3067_load_4_req_0;
      ptr_deref_3067_load_1_ack_0 <= ackL(7);
      ptr_deref_3067_load_5_ack_0 <= ackL(6);
      ptr_deref_3067_load_3_ack_0 <= ackL(5);
      ptr_deref_3067_load_2_ack_0 <= ackL(4);
      ptr_deref_3067_load_6_ack_0 <= ackL(3);
      ptr_deref_3067_load_7_ack_0 <= ackL(2);
      ptr_deref_3067_load_0_ack_0 <= ackL(1);
      ptr_deref_3067_load_4_ack_0 <= ackL(0);
      reqR(7) <= ptr_deref_3067_load_1_req_1;
      reqR(6) <= ptr_deref_3067_load_5_req_1;
      reqR(5) <= ptr_deref_3067_load_3_req_1;
      reqR(4) <= ptr_deref_3067_load_2_req_1;
      reqR(3) <= ptr_deref_3067_load_6_req_1;
      reqR(2) <= ptr_deref_3067_load_7_req_1;
      reqR(1) <= ptr_deref_3067_load_0_req_1;
      reqR(0) <= ptr_deref_3067_load_4_req_1;
      ptr_deref_3067_load_1_ack_1 <= ackR(7);
      ptr_deref_3067_load_5_ack_1 <= ackR(6);
      ptr_deref_3067_load_3_ack_1 <= ackR(5);
      ptr_deref_3067_load_2_ack_1 <= ackR(4);
      ptr_deref_3067_load_6_ack_1 <= ackR(3);
      ptr_deref_3067_load_7_ack_1 <= ackR(2);
      ptr_deref_3067_load_0_ack_1 <= ackR(1);
      ptr_deref_3067_load_4_ack_1 <= ackR(0);
      data_in <= ptr_deref_3067_word_address_1 & ptr_deref_3067_word_address_5 & ptr_deref_3067_word_address_3 & ptr_deref_3067_word_address_2 & ptr_deref_3067_word_address_6 & ptr_deref_3067_word_address_7 & ptr_deref_3067_word_address_0 & ptr_deref_3067_word_address_4;
      ptr_deref_3067_data_1 <= data_out(63 downto 56);
      ptr_deref_3067_data_5 <= data_out(55 downto 48);
      ptr_deref_3067_data_3 <= data_out(47 downto 40);
      ptr_deref_3067_data_2 <= data_out(39 downto 32);
      ptr_deref_3067_data_6 <= data_out(31 downto 24);
      ptr_deref_3067_data_7 <= data_out(23 downto 16);
      ptr_deref_3067_data_0 <= data_out(15 downto 8);
      ptr_deref_3067_data_4 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 8,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 8,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    xxsend_packet_pipelinexxblen_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxblen_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxblen_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxblen_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxblen_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxblen_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxblen_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxbuf64_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxpkt64_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxread_ctrl_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxread_last_word_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxread_last_word_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxread_last_word_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxread_last_word_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxread_last_word_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxread_last_word_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxread_last_word_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxread_pointer_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxread_pointer_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxread_pointer_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxread_pointer_pipe_read_data,
        write_req => xxsend_packet_pipelinexxread_pointer_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxread_pointer_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxread_pointer_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxswap_ctrl_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxswap_data_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxswap_data_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxswap_data_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxswap_data_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxswap_data_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxswap_data_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxswap_data_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxswap_last_word_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxwlen_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxwlen_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxwlen_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxwlen_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxwlen_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxwlen_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxwlen_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : simple_obj_ref_2935_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2935_inst_ack_0 then -- 
            assert false report " ReadPipe send_packet_pipe to wire pkt_2936 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2935_inst_req_0;
      simple_obj_ref_2935_inst_ack_0 <= ack(0);
      pkt_2936 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => send_packet_pipe_pipe_read_req(0),
          oack => send_packet_pipe_pipe_read_ack(0),
          odata => send_packet_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_2969_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2969_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxwlen_pipe to wire wlen_2970 value="  &  convert_slv_to_hex_string(data_out(15 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2969_inst_req_0;
      simple_obj_ref_2969_inst_ack_0 <= ack(0);
      wlen_2970 <= data_out(15 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxwlen_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxwlen_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxwlen_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_2972_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2972_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxblen_pipe to wire blen_2973 value="  &  convert_slv_to_hex_string(data_out(15 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2972_inst_req_0;
      simple_obj_ref_2972_inst_ack_0 <= ack(0);
      blen_2973 <= data_out(15 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxblen_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxblen_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxblen_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_2975_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2975_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxbuf64_pipe to wire buf64_2976 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2975_inst_req_0;
      simple_obj_ref_2975_inst_ack_0 <= ack(0);
      buf64_2976 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_2978_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2978_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxpkt64_pipe to wire pkt64_2979 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2978_inst_req_0;
      simple_obj_ref_2978_inst_ack_0 <= ack(0);
      pkt64_2979 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : simple_obj_ref_3062_inst 
    InportGroup5: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3062_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxread_pointer to wire ptr_3063 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3062_inst_req_0;
      simple_obj_ref_3062_inst_ack_0 <= ack(0);
      ptr_3063 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxread_pointer_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxread_pointer_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxread_pointer_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : simple_obj_ref_3070_inst 
    InportGroup6: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3070_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxread_ctrl_in to wire simple_obj_ref_3070_wire value="  &  convert_slv_to_hex_string(data_out(7 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3070_inst_req_0;
      simple_obj_ref_3070_inst_ack_0 <= ack(0);
      simple_obj_ref_3070_wire <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : simple_obj_ref_3073_inst 
    InportGroup7: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3073_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxread_last_word_in to wire simple_obj_ref_3073_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3073_inst_req_0;
      simple_obj_ref_3073_inst_ack_0 <= ack(0);
      simple_obj_ref_3073_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxread_last_word_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxread_last_word_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxread_last_word_in_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : simple_obj_ref_3081_inst 
    InportGroup8: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3081_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxswap_data_in to wire a_3082 value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3081_inst_req_0;
      simple_obj_ref_3081_inst_ack_0 <= ack(0);
      a_3082 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxswap_data_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxswap_data_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxswap_data_in_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : simple_obj_ref_3124_inst 
    InportGroup9: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3124_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxswap_ctrl_in to wire simple_obj_ref_3124_wire value="  &  convert_slv_to_hex_string(data_out(7 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3124_inst_req_0;
      simple_obj_ref_3124_inst_ack_0 <= ack(0);
      simple_obj_ref_3124_wire <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : simple_obj_ref_3128_inst 
    InportGroup10: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3128_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxswap_last_word_in to wire simple_obj_ref_3128_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3128_inst_req_0;
      simple_obj_ref_3128_inst_ack_0 <= ack(0);
      simple_obj_ref_3128_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : simple_obj_ref_3131_inst 
    InportGroup11: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3131_inst_ack_0 then -- 
            assert false report " ReadPipe send_packet_buf_queue to wire simple_obj_ref_3131_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3131_inst_req_0;
      simple_obj_ref_3131_inst_ack_0 <= ack(0);
      simple_obj_ref_3131_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => send_packet_buf_queue_pipe_read_req(0),
          oack => send_packet_buf_queue_pipe_read_ack(0),
          odata => send_packet_buf_queue_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2944_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxbuf64_pipe from wire type_cast_2946_wire value="  &  convert_slv_to_hex_string(type_cast_2946_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2944_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2944_inst_req_0;
      simple_obj_ref_2944_inst_ack_0 <= ack(0);
      data_in <= type_cast_2946_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2948_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxpkt64_pipe from wire type_cast_2950_wire value="  &  convert_slv_to_hex_string(type_cast_2950_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2948_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2948_inst_req_0;
      simple_obj_ref_2948_inst_ack_0 <= ack(0);
      data_in <= type_cast_2950_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2952_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxwlen_pipe from wire wlen_2942 value="  &  convert_slv_to_hex_string(wlen_2942) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (2) : simple_obj_ref_2952_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2952_inst_req_0;
      simple_obj_ref_2952_inst_ack_0 <= ack(0);
      data_in <= wlen_2942;
      outport: OutputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxwlen_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxwlen_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxwlen_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2955_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxblen_pipe from wire blen_2942 value="  &  convert_slv_to_hex_string(blen_2942) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (3) : simple_obj_ref_2955_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2955_inst_req_0;
      simple_obj_ref_2955_inst_ack_0 <= ack(0);
      data_in <= blen_2942;
      outport: OutputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxblen_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxblen_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxblen_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2958_inst_ack_0 then -- 
          assert false report " WritePipe send_packet_buf_queue from wire type_cast_2960_wire value="  &  convert_slv_to_hex_string(type_cast_2960_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (4) : simple_obj_ref_2958_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2958_inst_req_0;
      simple_obj_ref_2958_inst_ack_0 <= ack(0);
      data_in <= type_cast_2960_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => send_packet_buf_queue_pipe_write_req(0),
          oack => send_packet_buf_queue_pipe_write_ack(0),
          odata => send_packet_buf_queue_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3036_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_ctrl_in from wire binary_3047_wire value="  &  convert_slv_to_hex_string(binary_3047_wire) severity note; --
        end if;
        if simple_obj_ref_2986_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_ctrl_in from wire expr_2987_wire_constant value="  &  convert_slv_to_hex_string(expr_2987_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3009_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_ctrl_in from wire expr_3010_wire_constant value="  &  convert_slv_to_hex_string(expr_3010_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (5) : simple_obj_ref_3036_inst simple_obj_ref_2986_inst simple_obj_ref_3009_inst 
    OutportGroup5: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_3036_inst_req_0;
      req(1) <= simple_obj_ref_2986_inst_req_0;
      req(0) <= simple_obj_ref_3009_inst_req_0;
      simple_obj_ref_3036_inst_ack_0 <= ack(2);
      simple_obj_ref_2986_inst_ack_0 <= ack(1);
      simple_obj_ref_3009_inst_ack_0 <= ack(0);
      data_in <= binary_3047_wire & expr_2987_wire_constant & expr_3010_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 3,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3012_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_pointer from wire array_obj_ref_3014_wire value="  &  convert_slv_to_hex_string(array_obj_ref_3014_wire) severity note; --
        end if;
        if simple_obj_ref_2989_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_pointer from wire buf64_2976 value="  &  convert_slv_to_hex_string(buf64_2976) severity note; --
        end if;
        if simple_obj_ref_3049_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_pointer from wire last_word_ptr_3034 value="  &  convert_slv_to_hex_string(last_word_ptr_3034) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (6) : simple_obj_ref_3012_inst simple_obj_ref_2989_inst simple_obj_ref_3049_inst 
    OutportGroup6: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_3012_inst_req_0;
      req(1) <= simple_obj_ref_2989_inst_req_0;
      req(0) <= simple_obj_ref_3049_inst_req_0;
      simple_obj_ref_3012_inst_ack_0 <= ack(2);
      simple_obj_ref_2989_inst_ack_0 <= ack(1);
      simple_obj_ref_3049_inst_ack_0 <= ack(0);
      data_in <= array_obj_ref_3014_wire & buf64_2976 & last_word_ptr_3034;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 3,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxread_pointer_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxread_pointer_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxread_pointer_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2992_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_last_word_in from wire expr_2993_wire_constant value="  &  convert_slv_to_hex_string(expr_2993_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3016_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_last_word_in from wire expr_3017_wire_constant value="  &  convert_slv_to_hex_string(expr_3017_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3052_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_last_word_in from wire expr_3053_wire_constant value="  &  convert_slv_to_hex_string(expr_3053_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (7) : simple_obj_ref_2992_inst simple_obj_ref_3016_inst simple_obj_ref_3052_inst 
    OutportGroup7: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_2992_inst_req_0;
      req(1) <= simple_obj_ref_3016_inst_req_0;
      req(0) <= simple_obj_ref_3052_inst_req_0;
      simple_obj_ref_2992_inst_ack_0 <= ack(2);
      simple_obj_ref_3016_inst_ack_0 <= ack(1);
      simple_obj_ref_3052_inst_ack_0 <= ack(0);
      data_in <= expr_2993_wire_constant & expr_3017_wire_constant & expr_3053_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 3,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxread_last_word_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxread_last_word_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxread_last_word_in_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3065_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxswap_data_in from wire ptr_deref_3067_wire value="  &  convert_slv_to_hex_string(ptr_deref_3067_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (8) : simple_obj_ref_3065_inst 
    OutportGroup8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3065_inst_req_0;
      simple_obj_ref_3065_inst_ack_0 <= ack(0);
      data_in <= ptr_deref_3067_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxswap_data_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxswap_data_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxswap_data_in_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3069_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxswap_ctrl_in from wire simple_obj_ref_3070_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3070_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (9) : simple_obj_ref_3069_inst 
    OutportGroup9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3069_inst_req_0;
      simple_obj_ref_3069_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3070_wire;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 9
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3072_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxswap_last_word_in from wire simple_obj_ref_3073_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3073_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (10) : simple_obj_ref_3072_inst 
    OutportGroup10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3072_inst_req_0;
      simple_obj_ref_3072_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3073_wire;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 10
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3084_inst_ack_0 then -- 
          assert false report " WritePipe out_data from wire binary_3121_wire value="  &  convert_slv_to_hex_string(binary_3121_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (11) : simple_obj_ref_3084_inst 
    OutportGroup11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3084_inst_req_0;
      simple_obj_ref_3084_inst_ack_0 <= ack(0);
      data_in <= binary_3121_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 11
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3123_inst_ack_0 then -- 
          assert false report " WritePipe out_ctrl from wire simple_obj_ref_3124_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3124_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (12) : simple_obj_ref_3123_inst 
    OutportGroup12: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3123_inst_req_0;
      simple_obj_ref_3123_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3124_wire;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_ctrl_pipe_write_req(0),
          oack => out_ctrl_pipe_write_ack(0),
          odata => out_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 12
    -- shared call operator group (0) : call_stmt_2942_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_2942_call_req_0;
      call_stmt_2942_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_2942_call_req_1;
      call_stmt_2942_call_ack_1 <= ackR(0);
      data_in <= type_cast_2938_wire;
      buf_2942 <= data_out(63 downto 32);
      wlen_2942 <= data_out(31 downto 16);
      blen_2942 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 32,
        owidth => 32,
        twidth => 1,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => analyze_packet_call_reqs(0),
          ackR => analyze_packet_call_acks(0),
          dataR => analyze_packet_call_data(31 downto 0),
          tagR => analyze_packet_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 64, owidth => 64, twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => analyze_packet_return_acks(0), -- cross-over
          ackL => analyze_packet_return_reqs(0), -- cross-over
          dataL => analyze_packet_return_data(63 downto 0),
          tagL => analyze_packet_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_3132_call 
    CallGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3132_call_req_0;
      call_stmt_3132_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3132_call_req_1;
      call_stmt_3132_call_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_3131_wire;
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 32,
        owidth => 32,
        twidth => 3,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_packet_free_call_reqs(0),
          ackR => ahir_packet_free_call_acks(0),
          dataR => ahir_packet_free_call_data(31 downto 0),
          tagR => ahir_packet_free_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 3, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => ahir_packet_free_return_acks(0), -- cross-over
          ackL => ahir_packet_free_return_reqs(0), -- cross-over
          tagL => ahir_packet_free_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_input is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    receive_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    src_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    src_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    src_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
    free_queue_init_call_reqs : out  std_logic_vector(0 downto 0);
    free_queue_init_call_acks : in   std_logic_vector(0 downto 0);
    free_queue_init_call_tag  :  out  std_logic_vector(0 downto 0);
    free_queue_init_return_reqs : out  std_logic_vector(0 downto 0);
    free_queue_init_return_acks : in   std_logic_vector(0 downto 0);
    free_queue_init_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_input;
architecture Default of wrapper_input is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_input_CP_16042_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_3153_addr_0_ack_0 : boolean;
  signal call_stmt_3145_call_req_0 : boolean;
  signal simple_obj_ref_3160_inst_req_0 : boolean;
  signal ptr_deref_3153_store_0_ack_0 : boolean;
  signal ptr_deref_3153_root_address_inst_req_0 : boolean;
  signal ptr_deref_3158_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_3160_inst_ack_0 : boolean;
  signal ptr_deref_3153_addr_0_req_0 : boolean;
  signal ptr_deref_3153_base_resize_ack_0 : boolean;
  signal ptr_deref_3158_base_resize_req_0 : boolean;
  signal ptr_deref_3158_base_resize_ack_0 : boolean;
  signal ptr_deref_3153_store_0_ack_1 : boolean;
  signal ptr_deref_3153_store_0_req_1 : boolean;
  signal ptr_deref_3153_store_0_req_0 : boolean;
  signal ptr_deref_3153_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3158_gather_scatter_req_0 : boolean;
  signal ptr_deref_3153_gather_scatter_req_0 : boolean;
  signal ptr_deref_3158_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_3150_inst_req_0 : boolean;
  signal ptr_deref_3158_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3158_addr_0_req_0 : boolean;
  signal call_stmt_3145_call_ack_0 : boolean;
  signal ptr_deref_3158_addr_0_ack_0 : boolean;
  signal simple_obj_ref_3150_inst_ack_0 : boolean;
  signal ptr_deref_3153_gather_scatter_ack_0 : boolean;
  signal call_stmt_3146_call_req_0 : boolean;
  signal ptr_deref_3158_load_0_req_0 : boolean;
  signal call_stmt_3146_call_ack_0 : boolean;
  signal ptr_deref_3158_load_0_ack_0 : boolean;
  signal call_stmt_3145_call_req_1 : boolean;
  signal call_stmt_3145_call_ack_1 : boolean;
  signal call_stmt_3146_call_req_1 : boolean;
  signal call_stmt_3146_call_ack_1 : boolean;
  signal ptr_deref_3153_base_resize_req_0 : boolean;
  signal ptr_deref_3158_load_0_req_1 : boolean;
  signal ptr_deref_3158_load_0_ack_1 : boolean;
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_input_CP_16042: Block -- control-path 
    signal cp_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    crr_16078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => call_stmt_3145_call_req_0); -- 
    cp_elements(1) <= cp_elements(29);
    pipe_wreq_16225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => simple_obj_ref_3160_inst_req_0); -- 
    cp_elements(2) <= false; 
    cra_16079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3145_call_ack_0, ack => cp_elements(3)); -- 
    ccr_16083_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => call_stmt_3145_call_req_1); -- 
    cca_16084_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3145_call_ack_1, ack => cp_elements(4)); -- 
    crr_16095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => call_stmt_3146_call_req_0); -- 
    cra_16096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3146_call_ack_0, ack => cp_elements(5)); -- 
    ccr_16100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => call_stmt_3146_call_req_1); -- 
    cca_16101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3146_call_ack_1, ack => cp_elements(6)); -- 
    ack_16114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3150_inst_ack_0, ack => cp_elements(7)); -- 
    cp_elements(8) <= cp_elements(7);
    cp_elements(9) <= cp_elements(8);
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(9) & cp_elements(11) & cp_elements(15));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_3153_gather_scatter_req_0); -- 
    cp_elements(11) <= cp_elements(8);
    cp_elements(12) <= cp_elements(11);
    base_resize_req_16131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => ptr_deref_3153_base_resize_req_0); -- 
    base_resize_ack_16132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3153_base_resize_ack_0, ack => cp_elements(13)); -- 
    sum_rename_req_16136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_3153_root_address_inst_req_0); -- 
    sum_rename_ack_16137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3153_root_address_inst_ack_0, ack => cp_elements(14)); -- 
    root_rename_req_16141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => ptr_deref_3153_addr_0_req_0); -- 
    root_rename_ack_16142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3153_addr_0_ack_0, ack => cp_elements(15)); -- 
    split_ack_16147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3153_gather_scatter_ack_0, ack => cp_elements(16)); -- 
    rr_16154_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_3153_store_0_req_0); -- 
    cp_elements(17) <= ptr_deref_3153_store_0_ack_0;
    cp_elements(18) <= cp_elements(17);
    cr_16165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_3153_store_0_req_1); -- 
    ca_16166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3153_store_0_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(17) & cp_elements(21) & cp_elements(25));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_3158_load_0_req_0); -- 
    cp_elements(21) <= cp_elements(8);
    cp_elements(22) <= cp_elements(21);
    base_resize_req_16179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => ptr_deref_3158_base_resize_req_0); -- 
    base_resize_ack_16180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3158_base_resize_ack_0, ack => cp_elements(23)); -- 
    sum_rename_req_16184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => ptr_deref_3158_root_address_inst_req_0); -- 
    sum_rename_ack_16185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3158_root_address_inst_ack_0, ack => cp_elements(24)); -- 
    root_rename_req_16189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => ptr_deref_3158_addr_0_req_0); -- 
    root_rename_ack_16190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3158_addr_0_ack_0, ack => cp_elements(25)); -- 
    ra_16201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3158_load_0_ack_0, ack => cp_elements(26)); -- 
    cr_16211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => ptr_deref_3158_load_0_req_1); -- 
    ca_16212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3158_load_0_ack_1, ack => cp_elements(27)); -- 
    merge_req_16213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => ptr_deref_3158_gather_scatter_req_0); -- 
    merge_ack_16214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3158_gather_scatter_ack_0, ack => cp_elements(28)); -- 
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(28));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_16226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3160_inst_ack_0, ack => cp_elements(30)); -- 
    cp_elements(31) <= OrReduce(cp_elements(6) & cp_elements(30));
    cp_elements(32) <= cp_elements(31);
    req_16113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => simple_obj_ref_3150_inst_req_0); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal buf1_3144 : std_logic_vector(31 downto 0);
    signal iNsTr_4_3151 : std_logic_vector(31 downto 0);
    signal iNsTr_6_3159 : std_logic_vector(31 downto 0);
    signal ptr_deref_3153_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3153_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3153_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3153_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3153_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3153_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3158_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3158_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3158_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3158_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3158_word_offset_0 : std_logic_vector(0 downto 0);
    signal xxwrapper_inputxxbodyxxbuf1_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    buf1_3144 <= "00000000000000000000000000000000";
    ptr_deref_3153_word_offset_0 <= "0";
    ptr_deref_3158_word_offset_0 <= "0";
    xxwrapper_inputxxbodyxxbuf1_alloc_base_address <= "0";
    ptr_deref_3153_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => buf1_3144, dout => ptr_deref_3153_resized_base_address, req => ptr_deref_3153_base_resize_req_0, ack => ptr_deref_3153_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3158_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => buf1_3144, dout => ptr_deref_3158_resized_base_address, req => ptr_deref_3158_base_resize_req_0, ack => ptr_deref_3158_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3153_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3153_addr_0_ack_0 <= ptr_deref_3153_addr_0_req_0;
      aggregated_sig <= ptr_deref_3153_root_address;
      ptr_deref_3153_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3153_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3153_gather_scatter_ack_0 <= ptr_deref_3153_gather_scatter_req_0;
      aggregated_sig <= iNsTr_4_3151;
      ptr_deref_3153_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3153_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3153_root_address_inst_ack_0 <= ptr_deref_3153_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3153_resized_base_address;
      ptr_deref_3153_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3158_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3158_addr_0_ack_0 <= ptr_deref_3158_addr_0_req_0;
      aggregated_sig <= ptr_deref_3158_root_address;
      ptr_deref_3158_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3158_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3158_gather_scatter_ack_0 <= ptr_deref_3158_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3158_data_0;
      iNsTr_6_3159 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3158_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3158_root_address_inst_ack_0 <= ptr_deref_3158_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3158_resized_base_address;
      ptr_deref_3158_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    -- shared load operator group (0) : ptr_deref_3158_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3158_load_0_req_0,
        ptr_deref_3158_load_0_ack_0,
        ptr_deref_3158_load_0_req_1,
        ptr_deref_3158_load_0_ack_1,
        "ptr_deref_3158_load_0",
        "memory_space_7" ,
        ptr_deref_3158_data_0,
        ptr_deref_3158_word_address_0,
        "ptr_deref_3158_data_0",
        "ptr_deref_3158_word_address_0" -- 
      );
      reqL(0) <= ptr_deref_3158_load_0_req_0;
      ptr_deref_3158_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3158_load_0_req_1;
      ptr_deref_3158_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3158_word_address_0;
      ptr_deref_3158_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(31 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3153_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_7 address ptr_deref_3153_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3153_word_address_0) &  " data ptr_deref_3153_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3153_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_3153_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_3153_store_0_req_0;
      ptr_deref_3153_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3153_store_0_req_1;
      ptr_deref_3153_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3153_word_address_0;
      data_in <= ptr_deref_3153_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(31 downto 0),
          mtag => memory_space_7_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_3150_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3150_inst_ack_0 then -- 
            assert false report " ReadPipe receive_packet_pipe to wire iNsTr_4_3151 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3150_inst_req_0;
      simple_obj_ref_3150_inst_ack_0 <= ack(0);
      iNsTr_4_3151 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => receive_packet_pipe_pipe_read_req(0),
          oack => receive_packet_pipe_pipe_read_ack(0),
          odata => receive_packet_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3160_inst_ack_0 then -- 
          assert false report " WritePipe src_in0 from wire iNsTr_6_3159 value="  &  convert_slv_to_hex_string(iNsTr_6_3159) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3160_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3160_inst_req_0;
      simple_obj_ref_3160_inst_ack_0 <= ack(0);
      data_in <= iNsTr_6_3159;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => src_in0_pipe_write_req(0),
          oack => src_in0_pipe_write_ack(0),
          odata => src_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_3145_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3145_call_req_0;
      call_stmt_3145_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3145_call_req_1;
      call_stmt_3145_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => global_storage_initializer_x_call_reqs(0),
          ackR => global_storage_initializer_x_call_acks(0),
          tagR => global_storage_initializer_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => global_storage_initializer_x_return_acks(0), -- cross-over
          ackL => global_storage_initializer_x_return_reqs(0), -- cross-over
          tagL => global_storage_initializer_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_3146_call 
    CallGroup1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3146_call_req_0;
      call_stmt_3146_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3146_call_req_1;
      call_stmt_3146_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => free_queue_init_call_reqs(0),
          ackR => free_queue_init_call_acks(0),
          tagR => free_queue_init_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => free_queue_init_return_acks(0), -- cross-over
          ackL => free_queue_init_return_reqs(0), -- cross-over
          tagL => free_queue_init_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_output is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    tofpga0_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga1_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga2_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga3_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_read_data : in   std_logic_vector(31 downto 0);
    send_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_output;
architecture Default of wrapper_output is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_output_CP_16246_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_3231_store_0_req_0 : boolean;
  signal ptr_deref_3244_root_address_inst_ack_0 : boolean;
  signal type_cast_3228_inst_ack_0 : boolean;
  signal ptr_deref_3264_addr_0_ack_0 : boolean;
  signal ptr_deref_3244_store_0_ack_1 : boolean;
  signal ptr_deref_3231_root_address_inst_req_0 : boolean;
  signal type_cast_3254_inst_ack_0 : boolean;
  signal ptr_deref_3264_load_0_ack_1 : boolean;
  signal ptr_deref_3244_root_address_inst_req_0 : boolean;
  signal ptr_deref_3244_store_0_req_1 : boolean;
  signal type_cast_3241_inst_req_0 : boolean;
  signal ptr_deref_3264_load_0_req_1 : boolean;
  signal simple_obj_ref_3250_inst_req_0 : boolean;
  signal ptr_deref_3244_addr_0_req_0 : boolean;
  signal ptr_deref_3231_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3244_store_0_req_0 : boolean;
  signal type_cast_3268_inst_req_0 : boolean;
  signal type_cast_3268_inst_ack_0 : boolean;
  signal ptr_deref_3231_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3231_base_resize_req_0 : boolean;
  signal type_cast_3254_inst_req_0 : boolean;
  signal ptr_deref_3231_base_resize_ack_0 : boolean;
  signal type_cast_3241_inst_ack_0 : boolean;
  signal ptr_deref_3244_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3257_addr_0_req_0 : boolean;
  signal ptr_deref_3257_addr_0_ack_0 : boolean;
  signal ptr_deref_3231_store_0_ack_0 : boolean;
  signal ptr_deref_3244_addr_0_ack_0 : boolean;
  signal ptr_deref_3231_addr_0_req_0 : boolean;
  signal simple_obj_ref_3250_inst_ack_0 : boolean;
  signal simple_obj_ref_3237_inst_req_0 : boolean;
  signal ptr_deref_3231_addr_0_ack_0 : boolean;
  signal ptr_deref_3257_base_resize_req_0 : boolean;
  signal ptr_deref_3264_load_0_req_0 : boolean;
  signal ptr_deref_3257_base_resize_ack_0 : boolean;
  signal ptr_deref_3257_store_0_req_1 : boolean;
  signal ptr_deref_3257_store_0_ack_1 : boolean;
  signal simple_obj_ref_3237_inst_ack_0 : boolean;
  signal ptr_deref_3264_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3257_root_address_inst_req_0 : boolean;
  signal ptr_deref_3264_gather_scatter_req_0 : boolean;
  signal ptr_deref_3231_gather_scatter_req_0 : boolean;
  signal ptr_deref_3244_store_0_ack_0 : boolean;
  signal ptr_deref_3264_root_address_inst_req_0 : boolean;
  signal ptr_deref_3264_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3231_store_0_req_1 : boolean;
  signal ptr_deref_3264_addr_0_req_0 : boolean;
  signal simple_obj_ref_3270_inst_req_0 : boolean;
  signal simple_obj_ref_3270_inst_ack_0 : boolean;
  signal type_cast_3228_inst_req_0 : boolean;
  signal ptr_deref_3231_store_0_ack_1 : boolean;
  signal ptr_deref_3257_store_0_req_0 : boolean;
  signal ptr_deref_3257_store_0_ack_0 : boolean;
  signal ptr_deref_3244_base_resize_req_0 : boolean;
  signal ptr_deref_3244_base_resize_ack_0 : boolean;
  signal ptr_deref_3257_gather_scatter_req_0 : boolean;
  signal ptr_deref_3257_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3244_gather_scatter_req_0 : boolean;
  signal ptr_deref_3264_base_resize_req_0 : boolean;
  signal ptr_deref_3264_base_resize_ack_0 : boolean;
  signal ptr_deref_3264_load_0_ack_0 : boolean;
  signal ptr_deref_3257_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_3183_inst_req_0 : boolean;
  signal simple_obj_ref_3183_inst_ack_0 : boolean;
  signal ptr_deref_3186_base_resize_req_0 : boolean;
  signal ptr_deref_3186_base_resize_ack_0 : boolean;
  signal ptr_deref_3186_root_address_inst_req_0 : boolean;
  signal ptr_deref_3186_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3186_addr_0_req_0 : boolean;
  signal ptr_deref_3186_addr_0_ack_0 : boolean;
  signal ptr_deref_3186_gather_scatter_req_0 : boolean;
  signal ptr_deref_3186_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3186_store_0_req_0 : boolean;
  signal ptr_deref_3186_store_0_ack_0 : boolean;
  signal ptr_deref_3186_store_0_req_1 : boolean;
  signal ptr_deref_3186_store_0_ack_1 : boolean;
  signal ptr_deref_3191_base_resize_req_0 : boolean;
  signal ptr_deref_3191_base_resize_ack_0 : boolean;
  signal ptr_deref_3191_root_address_inst_req_0 : boolean;
  signal ptr_deref_3191_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3191_addr_0_req_0 : boolean;
  signal ptr_deref_3191_addr_0_ack_0 : boolean;
  signal ptr_deref_3191_load_0_req_0 : boolean;
  signal ptr_deref_3191_load_0_ack_0 : boolean;
  signal ptr_deref_3191_load_0_req_1 : boolean;
  signal ptr_deref_3191_load_0_ack_1 : boolean;
  signal ptr_deref_3191_gather_scatter_req_0 : boolean;
  signal ptr_deref_3191_gather_scatter_ack_0 : boolean;
  signal switch_stmt_3193_branch_default_req_0 : boolean;
  signal switch_stmt_3193_select_expr_0_req_0 : boolean;
  signal switch_stmt_3193_select_expr_0_ack_0 : boolean;
  signal switch_stmt_3193_select_expr_0_req_1 : boolean;
  signal switch_stmt_3193_select_expr_0_ack_1 : boolean;
  signal switch_stmt_3193_branch_0_req_0 : boolean;
  signal switch_stmt_3193_select_expr_1_req_0 : boolean;
  signal switch_stmt_3193_select_expr_1_ack_0 : boolean;
  signal switch_stmt_3193_select_expr_1_req_1 : boolean;
  signal switch_stmt_3193_select_expr_1_ack_1 : boolean;
  signal switch_stmt_3193_branch_1_req_0 : boolean;
  signal switch_stmt_3193_select_expr_2_req_0 : boolean;
  signal switch_stmt_3193_select_expr_2_ack_0 : boolean;
  signal switch_stmt_3193_select_expr_2_req_1 : boolean;
  signal switch_stmt_3193_select_expr_2_ack_1 : boolean;
  signal switch_stmt_3193_branch_2_req_0 : boolean;
  signal switch_stmt_3193_select_expr_3_req_0 : boolean;
  signal switch_stmt_3193_select_expr_3_ack_0 : boolean;
  signal switch_stmt_3193_select_expr_3_req_1 : boolean;
  signal switch_stmt_3193_select_expr_3_ack_1 : boolean;
  signal switch_stmt_3193_branch_3_req_0 : boolean;
  signal switch_stmt_3193_branch_0_ack_1 : boolean;
  signal switch_stmt_3193_branch_1_ack_1 : boolean;
  signal switch_stmt_3193_branch_2_ack_1 : boolean;
  signal switch_stmt_3193_branch_3_ack_1 : boolean;
  signal switch_stmt_3193_branch_default_ack_0 : boolean;
  signal simple_obj_ref_3211_inst_req_0 : boolean;
  signal simple_obj_ref_3211_inst_ack_0 : boolean;
  signal type_cast_3215_inst_req_0 : boolean;
  signal type_cast_3215_inst_ack_0 : boolean;
  signal ptr_deref_3218_base_resize_req_0 : boolean;
  signal ptr_deref_3218_base_resize_ack_0 : boolean;
  signal ptr_deref_3218_root_address_inst_req_0 : boolean;
  signal ptr_deref_3218_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3218_addr_0_req_0 : boolean;
  signal ptr_deref_3218_addr_0_ack_0 : boolean;
  signal ptr_deref_3218_gather_scatter_req_0 : boolean;
  signal ptr_deref_3218_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3218_store_0_req_0 : boolean;
  signal ptr_deref_3218_store_0_ack_0 : boolean;
  signal ptr_deref_3218_store_0_req_1 : boolean;
  signal ptr_deref_3218_store_0_ack_1 : boolean;
  signal simple_obj_ref_3224_inst_req_0 : boolean;
  signal simple_obj_ref_3224_inst_ack_0 : boolean;
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_9_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_9_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_output_CP_16246: Block -- control-path 
    signal cp_elements: BooleanArray(135 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(3);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(3), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(26);
    cp_elements(2) <= OrReduce(cp_elements(47) & cp_elements(133));
    req_16486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => simple_obj_ref_3211_inst_req_0); -- 
    cp_elements(3) <= false; 
    ack_16310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3183_inst_ack_0, ack => cp_elements(4)); -- 
    cp_elements(5) <= cp_elements(4);
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8) & cp_elements(12));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_3186_gather_scatter_req_0); -- 
    cp_elements(8) <= cp_elements(5);
    cp_elements(9) <= cp_elements(8);
    base_resize_req_16327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => ptr_deref_3186_base_resize_req_0); -- 
    base_resize_ack_16328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_base_resize_ack_0, ack => cp_elements(10)); -- 
    sum_rename_req_16332_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_3186_root_address_inst_req_0); -- 
    sum_rename_ack_16333_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_root_address_inst_ack_0, ack => cp_elements(11)); -- 
    root_rename_req_16337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => ptr_deref_3186_addr_0_req_0); -- 
    root_rename_ack_16338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_addr_0_ack_0, ack => cp_elements(12)); -- 
    split_ack_16343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_gather_scatter_ack_0, ack => cp_elements(13)); -- 
    rr_16350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_3186_store_0_req_0); -- 
    cp_elements(14) <= ptr_deref_3186_store_0_ack_0;
    cp_elements(15) <= cp_elements(14);
    cr_16361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => ptr_deref_3186_store_0_req_1); -- 
    ca_16362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_store_0_ack_1, ack => cp_elements(16)); -- 
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(18) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_3191_load_0_req_0); -- 
    cp_elements(18) <= cp_elements(5);
    cp_elements(19) <= cp_elements(18);
    base_resize_req_16375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => ptr_deref_3191_base_resize_req_0); -- 
    base_resize_ack_16376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3191_base_resize_ack_0, ack => cp_elements(20)); -- 
    sum_rename_req_16380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_3191_root_address_inst_req_0); -- 
    sum_rename_ack_16381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3191_root_address_inst_ack_0, ack => cp_elements(21)); -- 
    root_rename_req_16385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => ptr_deref_3191_addr_0_req_0); -- 
    root_rename_ack_16386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3191_addr_0_ack_0, ack => cp_elements(22)); -- 
    ra_16397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3191_load_0_ack_0, ack => cp_elements(23)); -- 
    cr_16407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => ptr_deref_3191_load_0_req_1); -- 
    ca_16408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3191_load_0_ack_1, ack => cp_elements(24)); -- 
    merge_req_16409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => ptr_deref_3191_gather_scatter_req_0); -- 
    merge_ack_16410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3191_gather_scatter_ack_0, ack => cp_elements(25)); -- 
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(25));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(27) <= cp_elements(1);
    cp_elements(28) <= false;
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= cp_elements(1);
    cp_elements(31) <= cp_elements(30);
    cp_elements(32) <= cp_elements(31);
    rr_16422_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => switch_stmt_3193_select_expr_0_req_0); -- 
    ra_16423_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_0_ack_0, ack => cp_elements(33)); -- 
    cr_16424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => switch_stmt_3193_select_expr_0_req_1); -- 
    ca_16425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_0_ack_1, ack => cp_elements(34)); -- 
    cmp_16426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => switch_stmt_3193_branch_0_req_0); -- 
    cp_elements(35) <= cp_elements(31);
    rr_16430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => switch_stmt_3193_select_expr_1_req_0); -- 
    ra_16431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_1_ack_0, ack => cp_elements(36)); -- 
    cr_16432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => switch_stmt_3193_select_expr_1_req_1); -- 
    ca_16433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_1_ack_1, ack => cp_elements(37)); -- 
    cmp_16434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => switch_stmt_3193_branch_1_req_0); -- 
    cp_elements(38) <= cp_elements(31);
    rr_16438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => switch_stmt_3193_select_expr_2_req_0); -- 
    ra_16439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_2_ack_0, ack => cp_elements(39)); -- 
    cr_16440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => switch_stmt_3193_select_expr_2_req_1); -- 
    ca_16441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_2_ack_1, ack => cp_elements(40)); -- 
    cmp_16442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => switch_stmt_3193_branch_2_req_0); -- 
    cp_elements(41) <= cp_elements(31);
    rr_16446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => switch_stmt_3193_select_expr_3_req_0); -- 
    ra_16447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_3_ack_0, ack => cp_elements(42)); -- 
    cr_16448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => switch_stmt_3193_select_expr_3_req_1); -- 
    ca_16449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_select_expr_3_ack_1, ack => cp_elements(43)); -- 
    cmp_16450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => switch_stmt_3193_branch_3_req_0); -- 
    cpelement_group_44 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(34) & cp_elements(37) & cp_elements(40) & cp_elements(43));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(44),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    Xexit_16418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => switch_stmt_3193_branch_default_req_0); -- 
    cp_elements(45) <= cp_elements(44);
    cp_elements(46) <= cp_elements(45);
    ack1_16455_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_branch_0_ack_1, ack => cp_elements(47)); -- 
    cp_elements(48) <= cp_elements(45);
    ack1_16460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_branch_1_ack_1, ack => cp_elements(49)); -- 
    req_16559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => simple_obj_ref_3224_inst_req_0); -- 
    cp_elements(50) <= cp_elements(45);
    ack1_16465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_branch_2_ack_1, ack => cp_elements(51)); -- 
    req_16632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => simple_obj_ref_3237_inst_req_0); -- 
    cp_elements(52) <= cp_elements(45);
    ack1_16470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_branch_3_ack_1, ack => cp_elements(53)); -- 
    req_16705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => simple_obj_ref_3250_inst_req_0); -- 
    cp_elements(54) <= cp_elements(45);
    ack0_16475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3193_branch_default_ack_0, ack => cp_elements(55)); -- 
    ack_16487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3211_inst_ack_0, ack => cp_elements(56)); -- 
    cp_elements(57) <= cp_elements(56);
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(59) & cp_elements(60));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => type_cast_3215_inst_req_0); -- 
    cp_elements(59) <= cp_elements(57);
    cp_elements(60) <= cp_elements(57);
    ack_16500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3215_inst_ack_0, ack => cp_elements(61)); -- 
    cpelement_group_62 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(63) & cp_elements(67));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(62),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_3218_gather_scatter_req_0); -- 
    cp_elements(63) <= cp_elements(57);
    cp_elements(64) <= cp_elements(63);
    base_resize_req_16514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => ptr_deref_3218_base_resize_req_0); -- 
    base_resize_ack_16515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3218_base_resize_ack_0, ack => cp_elements(65)); -- 
    sum_rename_req_16519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_3218_root_address_inst_req_0); -- 
    sum_rename_ack_16520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3218_root_address_inst_ack_0, ack => cp_elements(66)); -- 
    root_rename_req_16524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => ptr_deref_3218_addr_0_req_0); -- 
    root_rename_ack_16525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3218_addr_0_ack_0, ack => cp_elements(67)); -- 
    split_ack_16530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3218_gather_scatter_ack_0, ack => cp_elements(68)); -- 
    rr_16537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_3218_store_0_req_0); -- 
    ra_16538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3218_store_0_ack_0, ack => cp_elements(69)); -- 
    cr_16548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_3218_store_0_req_1); -- 
    ca_16549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3218_store_0_ack_1, ack => cp_elements(70)); -- 
    ack_16560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3224_inst_ack_0, ack => cp_elements(71)); -- 
    cp_elements(72) <= cp_elements(71);
    cpelement_group_73 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(74) & cp_elements(75));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(73),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => type_cast_3228_inst_req_0); -- 
    cp_elements(74) <= cp_elements(72);
    cp_elements(75) <= cp_elements(72);
    ack_16573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3228_inst_ack_0, ack => cp_elements(76)); -- 
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(78) & cp_elements(82));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_3231_gather_scatter_req_0); -- 
    cp_elements(78) <= cp_elements(72);
    cp_elements(79) <= cp_elements(78);
    base_resize_req_16587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_3231_base_resize_req_0); -- 
    base_resize_ack_16588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3231_base_resize_ack_0, ack => cp_elements(80)); -- 
    sum_rename_req_16592_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_3231_root_address_inst_req_0); -- 
    sum_rename_ack_16593_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3231_root_address_inst_ack_0, ack => cp_elements(81)); -- 
    root_rename_req_16597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_3231_addr_0_req_0); -- 
    root_rename_ack_16598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3231_addr_0_ack_0, ack => cp_elements(82)); -- 
    split_ack_16603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3231_gather_scatter_ack_0, ack => cp_elements(83)); -- 
    rr_16610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_3231_store_0_req_0); -- 
    ra_16611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3231_store_0_ack_0, ack => cp_elements(84)); -- 
    cr_16621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_3231_store_0_req_1); -- 
    ca_16622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3231_store_0_ack_1, ack => cp_elements(85)); -- 
    ack_16633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3237_inst_ack_0, ack => cp_elements(86)); -- 
    cp_elements(87) <= cp_elements(86);
    cpelement_group_88 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(88),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => type_cast_3241_inst_req_0); -- 
    cp_elements(89) <= cp_elements(87);
    cp_elements(90) <= cp_elements(87);
    ack_16646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3241_inst_ack_0, ack => cp_elements(91)); -- 
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(93) & cp_elements(97));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16675_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_3244_gather_scatter_req_0); -- 
    cp_elements(93) <= cp_elements(87);
    cp_elements(94) <= cp_elements(93);
    base_resize_req_16660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_3244_base_resize_req_0); -- 
    base_resize_ack_16661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3244_base_resize_ack_0, ack => cp_elements(95)); -- 
    sum_rename_req_16665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => ptr_deref_3244_root_address_inst_req_0); -- 
    sum_rename_ack_16666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3244_root_address_inst_ack_0, ack => cp_elements(96)); -- 
    root_rename_req_16670_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_3244_addr_0_req_0); -- 
    root_rename_ack_16671_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3244_addr_0_ack_0, ack => cp_elements(97)); -- 
    split_ack_16676_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3244_gather_scatter_ack_0, ack => cp_elements(98)); -- 
    rr_16683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_3244_store_0_req_0); -- 
    ra_16684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3244_store_0_ack_0, ack => cp_elements(99)); -- 
    cr_16694_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => ptr_deref_3244_store_0_req_1); -- 
    ca_16695_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3244_store_0_ack_1, ack => cp_elements(100)); -- 
    ack_16706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3250_inst_ack_0, ack => cp_elements(101)); -- 
    cp_elements(102) <= cp_elements(101);
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(104) & cp_elements(105));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => type_cast_3254_inst_req_0); -- 
    cp_elements(104) <= cp_elements(102);
    cp_elements(105) <= cp_elements(102);
    ack_16719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3254_inst_ack_0, ack => cp_elements(106)); -- 
    cpelement_group_107 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(106) & cp_elements(108) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_3257_gather_scatter_req_0); -- 
    cp_elements(108) <= cp_elements(102);
    cp_elements(109) <= cp_elements(108);
    base_resize_req_16733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_3257_base_resize_req_0); -- 
    base_resize_ack_16734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3257_base_resize_ack_0, ack => cp_elements(110)); -- 
    sum_rename_req_16738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ptr_deref_3257_root_address_inst_req_0); -- 
    sum_rename_ack_16739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3257_root_address_inst_ack_0, ack => cp_elements(111)); -- 
    root_rename_req_16743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_3257_addr_0_req_0); -- 
    root_rename_ack_16744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3257_addr_0_ack_0, ack => cp_elements(112)); -- 
    split_ack_16749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3257_gather_scatter_ack_0, ack => cp_elements(113)); -- 
    rr_16756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_3257_store_0_req_0); -- 
    ra_16757_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3257_store_0_ack_0, ack => cp_elements(114)); -- 
    cr_16767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => ptr_deref_3257_store_0_req_1); -- 
    ca_16768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3257_store_0_ack_1, ack => cp_elements(115)); -- 
    cp_elements(116) <= cp_elements(135);
    cpelement_group_117 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(122));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_3264_load_0_req_0); -- 
    cp_elements(118) <= cp_elements(116);
    cp_elements(119) <= cp_elements(118);
    base_resize_req_16784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_3264_base_resize_req_0); -- 
    base_resize_ack_16785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3264_base_resize_ack_0, ack => cp_elements(120)); -- 
    sum_rename_req_16789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => ptr_deref_3264_root_address_inst_req_0); -- 
    sum_rename_ack_16790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3264_root_address_inst_ack_0, ack => cp_elements(121)); -- 
    root_rename_req_16794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => ptr_deref_3264_addr_0_req_0); -- 
    root_rename_ack_16795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3264_addr_0_ack_0, ack => cp_elements(122)); -- 
    ra_16806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3264_load_0_ack_0, ack => cp_elements(123)); -- 
    cr_16816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_3264_load_0_req_1); -- 
    ca_16817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3264_load_0_ack_1, ack => cp_elements(124)); -- 
    merge_req_16818_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => ptr_deref_3264_gather_scatter_req_0); -- 
    merge_ack_16819_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3264_gather_scatter_ack_0, ack => cp_elements(125)); -- 
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(127));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => type_cast_3268_inst_req_0); -- 
    cp_elements(127) <= cp_elements(116);
    ack_16829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3268_inst_ack_0, ack => cp_elements(128)); -- 
    pipe_wreq_16840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => simple_obj_ref_3270_inst_req_0); -- 
    pipe_wack_16841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3270_inst_ack_0, ack => cp_elements(129)); -- 
    cp_elements(130) <= OrReduce(cp_elements(0) & cp_elements(129));
    cp_elements(131) <= cp_elements(130);
    req_16309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => simple_obj_ref_3183_inst_req_0); -- 
    cp_elements(132) <= false;
    cp_elements(133) <= cp_elements(132);
    cp_elements(134) <= OrReduce(cp_elements(55) & cp_elements(70) & cp_elements(85) & cp_elements(100) & cp_elements(115));
    cp_elements(135) <= cp_elements(134);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal expr_3195_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3195_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3198_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3198_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3201_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3201_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3204_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3204_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal iNsTr_12_3212 : std_logic_vector(31 downto 0);
    signal iNsTr_13_3216 : std_logic_vector(31 downto 0);
    signal iNsTr_17_3225 : std_logic_vector(31 downto 0);
    signal iNsTr_18_3229 : std_logic_vector(31 downto 0);
    signal iNsTr_22_3238 : std_logic_vector(31 downto 0);
    signal iNsTr_23_3242 : std_logic_vector(31 downto 0);
    signal iNsTr_27_3251 : std_logic_vector(31 downto 0);
    signal iNsTr_28_3255 : std_logic_vector(31 downto 0);
    signal iNsTr_2_3184 : std_logic_vector(31 downto 0);
    signal iNsTr_4_3192 : std_logic_vector(31 downto 0);
    signal iNsTr_6_3265 : std_logic_vector(31 downto 0);
    signal iNsTr_7_3269 : std_logic_vector(31 downto 0);
    signal pkt_3175 : std_logic_vector(31 downto 0);
    signal port_number_3179 : std_logic_vector(31 downto 0);
    signal ptr_deref_3186_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3186_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3186_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3186_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3186_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3186_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3191_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3191_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3191_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3191_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3191_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3218_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3218_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3218_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3218_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3218_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3218_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3231_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3231_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3231_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3231_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3231_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3231_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3244_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3244_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3244_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3244_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3244_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3244_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3257_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3257_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3257_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3257_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3257_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3257_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3264_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3264_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3264_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3264_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3264_word_offset_0 : std_logic_vector(0 downto 0);
    signal xxwrapper_outputxxbodyxxpkt_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxwrapper_outputxxbodyxxport_number_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    expr_3195_wire_constant <= "00000000000000000000000000000001";
    expr_3198_wire_constant <= "00000000000000000000000000000010";
    expr_3201_wire_constant <= "00000000000000000000000000000011";
    expr_3204_wire_constant <= "00000000000000000000000000000100";
    pkt_3175 <= "00000000000000000000000000000000";
    port_number_3179 <= "00000000000000000000000000000000";
    ptr_deref_3186_word_offset_0 <= "0";
    ptr_deref_3191_word_offset_0 <= "0";
    ptr_deref_3218_word_offset_0 <= "0";
    ptr_deref_3231_word_offset_0 <= "0";
    ptr_deref_3244_word_offset_0 <= "0";
    ptr_deref_3257_word_offset_0 <= "0";
    ptr_deref_3264_word_offset_0 <= "0";
    xxwrapper_outputxxbodyxxpkt_alloc_base_address <= "0";
    xxwrapper_outputxxbodyxxport_number_alloc_base_address <= "0";
    ptr_deref_3186_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => port_number_3179, dout => ptr_deref_3186_resized_base_address, req => ptr_deref_3186_base_resize_req_0, ack => ptr_deref_3186_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3191_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => port_number_3179, dout => ptr_deref_3191_resized_base_address, req => ptr_deref_3191_base_resize_req_0, ack => ptr_deref_3191_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3218_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3175, dout => ptr_deref_3218_resized_base_address, req => ptr_deref_3218_base_resize_req_0, ack => ptr_deref_3218_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3231_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3175, dout => ptr_deref_3231_resized_base_address, req => ptr_deref_3231_base_resize_req_0, ack => ptr_deref_3231_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3244_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3175, dout => ptr_deref_3244_resized_base_address, req => ptr_deref_3244_base_resize_req_0, ack => ptr_deref_3244_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3257_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3175, dout => ptr_deref_3257_resized_base_address, req => ptr_deref_3257_base_resize_req_0, ack => ptr_deref_3257_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3264_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3175, dout => ptr_deref_3264_resized_base_address, req => ptr_deref_3264_base_resize_req_0, ack => ptr_deref_3264_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_3215_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_12_3212, dout => iNsTr_13_3216, req => type_cast_3215_inst_req_0, ack => type_cast_3215_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3228_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_17_3225, dout => iNsTr_18_3229, req => type_cast_3228_inst_req_0, ack => type_cast_3228_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3241_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_22_3238, dout => iNsTr_23_3242, req => type_cast_3241_inst_req_0, ack => type_cast_3241_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3254_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_27_3251, dout => iNsTr_28_3255, req => type_cast_3254_inst_req_0, ack => type_cast_3254_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3268_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_6_3265, dout => iNsTr_7_3269, req => type_cast_3268_inst_req_0, ack => type_cast_3268_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3186_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3186_addr_0_ack_0 <= ptr_deref_3186_addr_0_req_0;
      aggregated_sig <= ptr_deref_3186_root_address;
      ptr_deref_3186_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3186_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3186_gather_scatter_ack_0 <= ptr_deref_3186_gather_scatter_req_0;
      aggregated_sig <= iNsTr_2_3184;
      ptr_deref_3186_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3186_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3186_root_address_inst_ack_0 <= ptr_deref_3186_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3186_resized_base_address;
      ptr_deref_3186_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3191_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3191_addr_0_ack_0 <= ptr_deref_3191_addr_0_req_0;
      aggregated_sig <= ptr_deref_3191_root_address;
      ptr_deref_3191_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3191_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3191_gather_scatter_ack_0 <= ptr_deref_3191_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3191_data_0;
      iNsTr_4_3192 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3191_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3191_root_address_inst_ack_0 <= ptr_deref_3191_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3191_resized_base_address;
      ptr_deref_3191_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3218_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3218_addr_0_ack_0 <= ptr_deref_3218_addr_0_req_0;
      aggregated_sig <= ptr_deref_3218_root_address;
      ptr_deref_3218_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3218_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3218_gather_scatter_ack_0 <= ptr_deref_3218_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_3216;
      ptr_deref_3218_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3218_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3218_root_address_inst_ack_0 <= ptr_deref_3218_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3218_resized_base_address;
      ptr_deref_3218_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3231_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3231_addr_0_ack_0 <= ptr_deref_3231_addr_0_req_0;
      aggregated_sig <= ptr_deref_3231_root_address;
      ptr_deref_3231_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3231_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3231_gather_scatter_ack_0 <= ptr_deref_3231_gather_scatter_req_0;
      aggregated_sig <= iNsTr_18_3229;
      ptr_deref_3231_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3231_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3231_root_address_inst_ack_0 <= ptr_deref_3231_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3231_resized_base_address;
      ptr_deref_3231_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3244_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3244_addr_0_ack_0 <= ptr_deref_3244_addr_0_req_0;
      aggregated_sig <= ptr_deref_3244_root_address;
      ptr_deref_3244_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3244_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3244_gather_scatter_ack_0 <= ptr_deref_3244_gather_scatter_req_0;
      aggregated_sig <= iNsTr_23_3242;
      ptr_deref_3244_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3244_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3244_root_address_inst_ack_0 <= ptr_deref_3244_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3244_resized_base_address;
      ptr_deref_3244_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3257_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3257_addr_0_ack_0 <= ptr_deref_3257_addr_0_req_0;
      aggregated_sig <= ptr_deref_3257_root_address;
      ptr_deref_3257_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3257_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3257_gather_scatter_ack_0 <= ptr_deref_3257_gather_scatter_req_0;
      aggregated_sig <= iNsTr_28_3255;
      ptr_deref_3257_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3257_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3257_root_address_inst_ack_0 <= ptr_deref_3257_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3257_resized_base_address;
      ptr_deref_3257_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3264_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3264_addr_0_ack_0 <= ptr_deref_3264_addr_0_req_0;
      aggregated_sig <= ptr_deref_3264_root_address;
      ptr_deref_3264_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3264_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3264_gather_scatter_ack_0 <= ptr_deref_3264_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3264_data_0;
      iNsTr_6_3265 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3264_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3264_root_address_inst_ack_0 <= ptr_deref_3264_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3264_resized_base_address;
      ptr_deref_3264_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    switch_stmt_3193_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3195_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3193_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_3193_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3193_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3198_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3193_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_3193_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3193_branch_2: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3201_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3193_branch_2_req_0,
          ack0 => open,
          ack1 => switch_stmt_3193_branch_2_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3193_branch_3: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3204_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3193_branch_3_req_0,
          ack0 => open,
          ack1 => switch_stmt_3193_branch_3_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3193_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(3 downto 0);
      begin 
      condition_sig <= expr_3195_wire_constant_cmp & expr_3198_wire_constant_cmp & expr_3201_wire_constant_cmp & expr_3204_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 4)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3193_branch_default_req_0,
          ack0 => switch_stmt_3193_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : switch_stmt_3193_select_expr_0 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3192;
      expr_3195_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3193_select_expr_0_req_0,
          ackL => switch_stmt_3193_select_expr_0_ack_0,
          reqR => switch_stmt_3193_select_expr_0_req_1,
          ackR => switch_stmt_3193_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : switch_stmt_3193_select_expr_1 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3192;
      expr_3198_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3193_select_expr_1_req_0,
          ackL => switch_stmt_3193_select_expr_1_ack_0,
          reqR => switch_stmt_3193_select_expr_1_req_1,
          ackR => switch_stmt_3193_select_expr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : switch_stmt_3193_select_expr_2 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3192;
      expr_3201_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3193_select_expr_2_req_0,
          ackL => switch_stmt_3193_select_expr_2_ack_0,
          reqR => switch_stmt_3193_select_expr_2_req_1,
          ackR => switch_stmt_3193_select_expr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : switch_stmt_3193_select_expr_3 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3192;
      expr_3204_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3193_select_expr_3_req_0,
          ackL => switch_stmt_3193_select_expr_3_ack_0,
          reqR => switch_stmt_3193_select_expr_3_req_1,
          ackR => switch_stmt_3193_select_expr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared load operator group (0) : ptr_deref_3191_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3191_load_0_req_0,
        ptr_deref_3191_load_0_ack_0,
        ptr_deref_3191_load_0_req_1,
        ptr_deref_3191_load_0_ack_1,
        "ptr_deref_3191_load_0",
        "memory_space_9" ,
        ptr_deref_3191_data_0,
        ptr_deref_3191_word_address_0,
        "ptr_deref_3191_data_0",
        "ptr_deref_3191_word_address_0" -- 
      );
      reqL(0) <= ptr_deref_3191_load_0_req_0;
      ptr_deref_3191_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3191_load_0_req_1;
      ptr_deref_3191_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3191_word_address_0;
      ptr_deref_3191_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_9_lr_req(0),
          mack => memory_space_9_lr_ack(0),
          maddr => memory_space_9_lr_addr(0 downto 0),
          mtag => memory_space_9_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_9_lc_req(0),
          mack => memory_space_9_lc_ack(0),
          mdata => memory_space_9_lc_data(31 downto 0),
          mtag => memory_space_9_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_3264_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3264_load_0_req_0,
        ptr_deref_3264_load_0_ack_0,
        ptr_deref_3264_load_0_req_1,
        ptr_deref_3264_load_0_ack_1,
        "ptr_deref_3264_load_0",
        "memory_space_8" ,
        ptr_deref_3264_data_0,
        ptr_deref_3264_word_address_0,
        "ptr_deref_3264_data_0",
        "ptr_deref_3264_word_address_0" -- 
      );
      reqL(0) <= ptr_deref_3264_load_0_req_0;
      ptr_deref_3264_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3264_load_0_req_1;
      ptr_deref_3264_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3264_word_address_0;
      ptr_deref_3264_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(31 downto 0),
          mtag => memory_space_8_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3186_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_9 address ptr_deref_3186_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3186_word_address_0) &  " data ptr_deref_3186_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3186_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_3186_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_3186_store_0_req_0;
      ptr_deref_3186_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3186_store_0_req_1;
      ptr_deref_3186_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3186_word_address_0;
      data_in <= ptr_deref_3186_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(0 downto 0),
          mdata => memory_space_9_sr_data(31 downto 0),
          mtag => memory_space_9_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3218_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3218_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3218_word_address_0) &  " data ptr_deref_3218_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3218_data_0) severity note; --
        end if;
        if ptr_deref_3231_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3231_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3231_word_address_0) &  " data ptr_deref_3231_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3231_data_0) severity note; --
        end if;
        if ptr_deref_3244_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3244_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3244_word_address_0) &  " data ptr_deref_3244_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3244_data_0) severity note; --
        end if;
        if ptr_deref_3257_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3257_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3257_word_address_0) &  " data ptr_deref_3257_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3257_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (1) : ptr_deref_3218_store_0 ptr_deref_3231_store_0 ptr_deref_3244_store_0 ptr_deref_3257_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      -- 
    begin -- 
      reqL(3) <= ptr_deref_3218_store_0_req_0;
      reqL(2) <= ptr_deref_3231_store_0_req_0;
      reqL(1) <= ptr_deref_3244_store_0_req_0;
      reqL(0) <= ptr_deref_3257_store_0_req_0;
      ptr_deref_3218_store_0_ack_0 <= ackL(3);
      ptr_deref_3231_store_0_ack_0 <= ackL(2);
      ptr_deref_3244_store_0_ack_0 <= ackL(1);
      ptr_deref_3257_store_0_ack_0 <= ackL(0);
      reqR(3) <= ptr_deref_3218_store_0_req_1;
      reqR(2) <= ptr_deref_3231_store_0_req_1;
      reqR(1) <= ptr_deref_3244_store_0_req_1;
      reqR(0) <= ptr_deref_3257_store_0_req_1;
      ptr_deref_3218_store_0_ack_1 <= ackR(3);
      ptr_deref_3231_store_0_ack_1 <= ackR(2);
      ptr_deref_3244_store_0_ack_1 <= ackR(1);
      ptr_deref_3257_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3218_word_address_0 & ptr_deref_3231_word_address_0 & ptr_deref_3244_word_address_0 & ptr_deref_3257_word_address_0;
      data_in <= ptr_deref_3218_data_0 & ptr_deref_3231_data_0 & ptr_deref_3244_data_0 & ptr_deref_3257_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(31 downto 0),
          mtag => memory_space_8_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 4,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : simple_obj_ref_3183_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3183_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga_port_number to wire iNsTr_2_3184 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3183_inst_req_0;
      simple_obj_ref_3183_inst_ack_0 <= ack(0);
      iNsTr_2_3184 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga_port_number_pipe_read_req(0),
          oack => tofpga_port_number_pipe_read_ack(0),
          odata => tofpga_port_number_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_3211_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3211_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga0_out0 to wire iNsTr_12_3212 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3211_inst_req_0;
      simple_obj_ref_3211_inst_ack_0 <= ack(0);
      iNsTr_12_3212 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga0_out0_pipe_read_req(0),
          oack => tofpga0_out0_pipe_read_ack(0),
          odata => tofpga0_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_3224_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3224_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga1_out0 to wire iNsTr_17_3225 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3224_inst_req_0;
      simple_obj_ref_3224_inst_ack_0 <= ack(0);
      iNsTr_17_3225 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga1_out0_pipe_read_req(0),
          oack => tofpga1_out0_pipe_read_ack(0),
          odata => tofpga1_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_3237_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3237_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga2_out0 to wire iNsTr_22_3238 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3237_inst_req_0;
      simple_obj_ref_3237_inst_ack_0 <= ack(0);
      iNsTr_22_3238 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga2_out0_pipe_read_req(0),
          oack => tofpga2_out0_pipe_read_ack(0),
          odata => tofpga2_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_3250_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3250_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga3_out0 to wire iNsTr_27_3251 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3250_inst_req_0;
      simple_obj_ref_3250_inst_ack_0 <= ack(0);
      iNsTr_27_3251 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga3_out0_pipe_read_req(0),
          oack => tofpga3_out0_pipe_read_ack(0),
          odata => tofpga3_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3270_inst_ack_0 then -- 
          assert false report " WritePipe send_packet_pipe from wire iNsTr_7_3269 value="  &  convert_slv_to_hex_string(iNsTr_7_3269) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3270_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3270_inst_req_0;
      simple_obj_ref_3270_inst_ack_0 <= ack(0);
      data_in <= iNsTr_7_3269;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => send_packet_pipe_pipe_write_req(0),
          oack => send_packet_pipe_pipe_write_ack(0),
          odata => send_packet_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_9: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_9_lr_addr,
      lr_req_in => memory_space_9_lr_req,
      lr_ack_out => memory_space_9_lr_ack,
      lr_tag_in => memory_space_9_lr_tag,
      lc_req_in => memory_space_9_lc_req,
      lc_ack_out => memory_space_9_lc_ack,
      lc_data_out => memory_space_9_lc_data,
      lc_tag_out => memory_space_9_lc_tag,
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
    in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
    in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
    out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(8 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(8 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(143 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(98 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(8 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(8 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(71 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(44 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(6 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(6 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(111 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(55 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(76 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(6 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(6 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(34 downto 0);
  -- declarations related to module GV_15_initializer_in_click_bc
  component GV_15_initializer_in_click_bc is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module GV_15_initializer_in_click_bc
  signal GV_15_initializer_in_click_bc_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal GV_15_initializer_in_click_bc_tag_out   : std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_start_req : std_logic;
  signal GV_15_initializer_in_click_bc_start_ack : std_logic;
  signal GV_15_initializer_in_click_bc_fin_req   : std_logic;
  signal GV_15_initializer_in_click_bc_fin_ack : std_logic;
  -- caller side aggregated signals for module GV_15_initializer_in_click_bc
  signal GV_15_initializer_in_click_bc_call_reqs: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_call_acks: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_return_reqs: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_return_acks: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_call_tag: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module GV_16_initializer_in_click_bc
  component GV_16_initializer_in_click_bc is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module GV_16_initializer_in_click_bc
  signal GV_16_initializer_in_click_bc_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal GV_16_initializer_in_click_bc_tag_out   : std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_start_req : std_logic;
  signal GV_16_initializer_in_click_bc_start_ack : std_logic;
  signal GV_16_initializer_in_click_bc_fin_req   : std_logic;
  signal GV_16_initializer_in_click_bc_fin_ack : std_logic;
  -- caller side aggregated signals for module GV_16_initializer_in_click_bc
  signal GV_16_initializer_in_click_bc_call_reqs: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_call_acks: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_return_reqs: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_return_acks: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_call_tag: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module ahir_glue_bswap_i16
  component ahir_glue_bswap_i16 is -- 
    generic (tag_length : integer); 
    port ( -- 
      i : in  std_logic_vector(15 downto 0);
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_bswap_i16
  signal ahir_glue_bswap_i16_i :  std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_in_args    : std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_out_args   : std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal ahir_glue_bswap_i16_tag_out   : std_logic_vector(2 downto 0);
  signal ahir_glue_bswap_i16_start_req : std_logic;
  signal ahir_glue_bswap_i16_start_ack : std_logic;
  signal ahir_glue_bswap_i16_fin_req   : std_logic;
  signal ahir_glue_bswap_i16_fin_ack : std_logic;
  -- caller side aggregated signals for module ahir_glue_bswap_i16
  signal ahir_glue_bswap_i16_call_reqs: std_logic_vector(5 downto 0);
  signal ahir_glue_bswap_i16_call_acks: std_logic_vector(5 downto 0);
  signal ahir_glue_bswap_i16_return_reqs: std_logic_vector(5 downto 0);
  signal ahir_glue_bswap_i16_return_acks: std_logic_vector(5 downto 0);
  signal ahir_glue_bswap_i16_call_data: std_logic_vector(95 downto 0);
  signal ahir_glue_bswap_i16_call_tag: std_logic_vector(11 downto 0);
  signal ahir_glue_bswap_i16_return_data: std_logic_vector(95 downto 0);
  signal ahir_glue_bswap_i16_return_tag: std_logic_vector(11 downto 0);
  -- declarations related to module ahir_glue_chk
  component ahir_glue_chk is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      chk_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      chk_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      chk_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      rtt_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      rtt_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      rtt_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      ahir_packet_free_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_free_call_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_free_call_data : out  std_logic_vector(31 downto 0);
      ahir_packet_free_call_tag  :  out  std_logic_vector(2 downto 0);
      ahir_packet_free_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_free_return_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_free_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_chk
  signal ahir_glue_chk_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_chk_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_chk_start_req : std_logic;
  signal ahir_glue_chk_start_ack : std_logic;
  signal ahir_glue_chk_fin_req   : std_logic;
  signal ahir_glue_chk_fin_ack : std_logic;
  -- declarations related to module ahir_glue_rtt
  component ahir_glue_rtt is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(4 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      rtt_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      rtt_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rtt_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      to0_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to0_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to0_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      to1_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to1_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to1_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      to2_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to2_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to2_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      to3_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to3_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to3_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_packet_free_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_free_call_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_free_call_data : out  std_logic_vector(31 downto 0);
      ahir_packet_free_call_tag  :  out  std_logic_vector(2 downto 0);
      ahir_packet_free_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_free_return_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_free_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_rtt
  signal ahir_glue_rtt_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_rtt_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_rtt_start_req : std_logic;
  signal ahir_glue_rtt_start_ack : std_logic;
  signal ahir_glue_rtt_fin_req   : std_logic;
  signal ahir_glue_rtt_fin_ack : std_logic;
  -- declarations related to module ahir_glue_src
  component ahir_glue_src is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      src_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      src_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      src_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      chk_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      chk_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      chk_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_src
  signal ahir_glue_src_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_src_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_src_start_req : std_logic;
  signal ahir_glue_src_start_ack : std_logic;
  signal ahir_glue_src_fin_req   : std_logic;
  signal ahir_glue_src_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to0
  component ahir_glue_to0 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to0_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to0_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to0_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga0_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to0
  signal ahir_glue_to0_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to0_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to0_start_req : std_logic;
  signal ahir_glue_to0_start_ack : std_logic;
  signal ahir_glue_to0_fin_req   : std_logic;
  signal ahir_glue_to0_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to1
  component ahir_glue_to1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to1_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to1_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to1_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga1_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to1
  signal ahir_glue_to1_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to1_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to1_start_req : std_logic;
  signal ahir_glue_to1_start_ack : std_logic;
  signal ahir_glue_to1_fin_req   : std_logic;
  signal ahir_glue_to1_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to2
  component ahir_glue_to2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to2_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to2_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to2_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga2_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to2
  signal ahir_glue_to2_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to2_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to2_start_req : std_logic;
  signal ahir_glue_to2_start_ack : std_logic;
  signal ahir_glue_to2_fin_req   : std_logic;
  signal ahir_glue_to2_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to3
  component ahir_glue_to3 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to3_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to3_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to3_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga3_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to3
  signal ahir_glue_to3_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to3_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to3_start_req : std_logic;
  signal ahir_glue_to3_start_ack : std_logic;
  signal ahir_glue_to3_fin_req   : std_logic;
  signal ahir_glue_to3_fin_ack : std_logic;
  -- declarations related to module ahir_packet_free
  component ahir_packet_free is -- 
    generic (tag_length : integer); 
    port ( -- 
      pkt : in  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_packet_free
  signal ahir_packet_free_pkt :  std_logic_vector(31 downto 0);
  signal ahir_packet_free_in_args    : std_logic_vector(31 downto 0);
  signal ahir_packet_free_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ahir_packet_free_tag_out   : std_logic_vector(1 downto 0);
  signal ahir_packet_free_start_req : std_logic;
  signal ahir_packet_free_start_ack : std_logic;
  signal ahir_packet_free_fin_req   : std_logic;
  signal ahir_packet_free_fin_ack : std_logic;
  -- caller side aggregated signals for module ahir_packet_free
  signal ahir_packet_free_call_reqs: std_logic_vector(2 downto 0);
  signal ahir_packet_free_call_acks: std_logic_vector(2 downto 0);
  signal ahir_packet_free_return_reqs: std_logic_vector(2 downto 0);
  signal ahir_packet_free_return_acks: std_logic_vector(2 downto 0);
  signal ahir_packet_free_call_data: std_logic_vector(95 downto 0);
  signal ahir_packet_free_call_tag: std_logic_vector(8 downto 0);
  signal ahir_packet_free_return_tag: std_logic_vector(8 downto 0);
  -- declarations related to module ahir_packet_get
  component ahir_packet_get is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      free_queue_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_packet_get
  signal ahir_packet_get_buf :  std_logic_vector(31 downto 0);
  signal ahir_packet_get_out_args   : std_logic_vector(31 downto 0);
  signal ahir_packet_get_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_packet_get_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_packet_get_start_req : std_logic;
  signal ahir_packet_get_start_ack : std_logic;
  signal ahir_packet_get_fin_req   : std_logic;
  signal ahir_packet_get_fin_ack : std_logic;
  -- caller side aggregated signals for module ahir_packet_get
  signal ahir_packet_get_call_reqs: std_logic_vector(0 downto 0);
  signal ahir_packet_get_call_acks: std_logic_vector(0 downto 0);
  signal ahir_packet_get_return_reqs: std_logic_vector(0 downto 0);
  signal ahir_packet_get_return_acks: std_logic_vector(0 downto 0);
  signal ahir_packet_get_call_tag: std_logic_vector(0 downto 0);
  signal ahir_packet_get_return_data: std_logic_vector(31 downto 0);
  signal ahir_packet_get_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module analyze_packet
  component analyze_packet is -- 
    generic (tag_length : integer); 
    port ( -- 
      pkt : in  std_logic_vector(31 downto 0);
      buf : out  std_logic_vector(31 downto 0);
      wlen : out  std_logic_vector(15 downto 0);
      blen : out  std_logic_vector(15 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module analyze_packet
  signal analyze_packet_pkt :  std_logic_vector(31 downto 0);
  signal analyze_packet_buf :  std_logic_vector(31 downto 0);
  signal analyze_packet_wlen :  std_logic_vector(15 downto 0);
  signal analyze_packet_blen :  std_logic_vector(15 downto 0);
  signal analyze_packet_in_args    : std_logic_vector(31 downto 0);
  signal analyze_packet_out_args   : std_logic_vector(63 downto 0);
  signal analyze_packet_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal analyze_packet_tag_out   : std_logic_vector(0 downto 0);
  signal analyze_packet_start_req : std_logic;
  signal analyze_packet_start_ack : std_logic;
  signal analyze_packet_fin_req   : std_logic;
  signal analyze_packet_fin_ack : std_logic;
  -- caller side aggregated signals for module analyze_packet
  signal analyze_packet_call_reqs: std_logic_vector(0 downto 0);
  signal analyze_packet_call_acks: std_logic_vector(0 downto 0);
  signal analyze_packet_return_reqs: std_logic_vector(0 downto 0);
  signal analyze_packet_return_acks: std_logic_vector(0 downto 0);
  signal analyze_packet_call_data: std_logic_vector(31 downto 0);
  signal analyze_packet_call_tag: std_logic_vector(0 downto 0);
  signal analyze_packet_return_data: std_logic_vector(63 downto 0);
  signal analyze_packet_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module click_bc_storage_initializer_x
  component click_bc_storage_initializer_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      GV_15_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module click_bc_storage_initializer_x
  signal click_bc_storage_initializer_x_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal click_bc_storage_initializer_x_tag_out   : std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_start_req : std_logic;
  signal click_bc_storage_initializer_x_start_ack : std_logic;
  signal click_bc_storage_initializer_x_fin_req   : std_logic;
  signal click_bc_storage_initializer_x_fin_ack : std_logic;
  -- caller side aggregated signals for module click_bc_storage_initializer_x
  signal click_bc_storage_initializer_x_call_reqs: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_call_acks: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_return_reqs: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_return_acks: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_call_tag: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module free_queue_init
  component free_queue_init is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_init
  signal free_queue_init_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal free_queue_init_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_init_start_req : std_logic;
  signal free_queue_init_start_ack : std_logic;
  signal free_queue_init_fin_req   : std_logic;
  signal free_queue_init_fin_ack : std_logic;
  -- caller side aggregated signals for module free_queue_init
  signal free_queue_init_call_reqs: std_logic_vector(0 downto 0);
  signal free_queue_init_call_acks: std_logic_vector(0 downto 0);
  signal free_queue_init_return_reqs: std_logic_vector(0 downto 0);
  signal free_queue_init_return_acks: std_logic_vector(0 downto 0);
  signal free_queue_init_call_tag: std_logic_vector(0 downto 0);
  signal free_queue_init_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module global_storage_initializer_x
  component global_storage_initializer_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      click_bc_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module global_storage_initializer_x
  signal global_storage_initializer_x_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal global_storage_initializer_x_tag_out   : std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_start_req : std_logic;
  signal global_storage_initializer_x_start_ack : std_logic;
  signal global_storage_initializer_x_fin_req   : std_logic;
  signal global_storage_initializer_x_fin_ack : std_logic;
  -- caller side aggregated signals for module global_storage_initializer_x
  signal global_storage_initializer_x_call_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_tag: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module receive_packet_pipeline
  component receive_packet_pipeline is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      receive_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
      swapped_in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      swapped_in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      swapped_in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      receive_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
      swapped_in_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      swapped_in_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      swapped_in_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      receive_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_packet_get_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_get_call_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_get_call_tag  :  out  std_logic_vector(0 downto 0);
      ahir_packet_get_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_get_return_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_get_return_data : in   std_logic_vector(31 downto 0);
      ahir_packet_get_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module receive_packet_pipeline
  signal receive_packet_pipeline_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal receive_packet_pipeline_tag_out   : std_logic_vector(0 downto 0);
  signal receive_packet_pipeline_start_req : std_logic;
  signal receive_packet_pipeline_start_ack : std_logic;
  signal receive_packet_pipeline_fin_req   : std_logic;
  signal receive_packet_pipeline_fin_ack : std_logic;
  -- declarations related to module send_packet_pipeline
  component send_packet_pipeline is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      send_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
      send_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      send_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_packet_free_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_free_call_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_free_call_data : out  std_logic_vector(31 downto 0);
      ahir_packet_free_call_tag  :  out  std_logic_vector(2 downto 0);
      ahir_packet_free_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_packet_free_return_acks : in   std_logic_vector(0 downto 0);
      ahir_packet_free_return_tag :  in   std_logic_vector(2 downto 0);
      analyze_packet_call_reqs : out  std_logic_vector(0 downto 0);
      analyze_packet_call_acks : in   std_logic_vector(0 downto 0);
      analyze_packet_call_data : out  std_logic_vector(31 downto 0);
      analyze_packet_call_tag  :  out  std_logic_vector(0 downto 0);
      analyze_packet_return_reqs : out  std_logic_vector(0 downto 0);
      analyze_packet_return_acks : in   std_logic_vector(0 downto 0);
      analyze_packet_return_data : in   std_logic_vector(63 downto 0);
      analyze_packet_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module send_packet_pipeline
  signal send_packet_pipeline_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal send_packet_pipeline_tag_out   : std_logic_vector(0 downto 0);
  signal send_packet_pipeline_start_req : std_logic;
  signal send_packet_pipeline_start_ack : std_logic;
  signal send_packet_pipeline_fin_req   : std_logic;
  signal send_packet_pipeline_fin_ack : std_logic;
  -- declarations related to module wrapper_input
  component wrapper_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      receive_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      src_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      src_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      src_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
      free_queue_init_call_reqs : out  std_logic_vector(0 downto 0);
      free_queue_init_call_acks : in   std_logic_vector(0 downto 0);
      free_queue_init_call_tag  :  out  std_logic_vector(0 downto 0);
      free_queue_init_return_reqs : out  std_logic_vector(0 downto 0);
      free_queue_init_return_acks : in   std_logic_vector(0 downto 0);
      free_queue_init_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_input
  signal wrapper_input_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_input_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic;
  signal wrapper_input_start_ack : std_logic;
  signal wrapper_input_fin_req   : std_logic;
  signal wrapper_input_fin_ack : std_logic;
  -- declarations related to module wrapper_output
  component wrapper_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tofpga0_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga1_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga2_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga3_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_read_data : in   std_logic_vector(31 downto 0);
      send_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_output
  signal wrapper_output_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_output_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic;
  signal wrapper_output_start_ack : std_logic;
  signal wrapper_output_fin_req   : std_logic;
  signal wrapper_output_fin_ack : std_logic;
  -- aggregate signals for write to pipe chk_in0
  signal chk_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal chk_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal chk_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe chk_in0
  signal chk_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal chk_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal chk_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_pipe
  signal free_queue_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal free_queue_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal free_queue_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe free_queue_pipe
  signal free_queue_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_ctrl
  signal in_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_ctrl
  signal out_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe receive_packet_buf_queue
  signal receive_packet_buf_queue_pipe_write_data: std_logic_vector(31 downto 0);
  signal receive_packet_buf_queue_pipe_write_req: std_logic_vector(0 downto 0);
  signal receive_packet_buf_queue_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe receive_packet_buf_queue
  signal receive_packet_buf_queue_pipe_read_data: std_logic_vector(31 downto 0);
  signal receive_packet_buf_queue_pipe_read_req: std_logic_vector(0 downto 0);
  signal receive_packet_buf_queue_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe receive_packet_pipe
  signal receive_packet_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal receive_packet_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal receive_packet_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe receive_packet_pipe
  signal receive_packet_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal receive_packet_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal receive_packet_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe rtt_in0
  signal rtt_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal rtt_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal rtt_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe rtt_in0
  signal rtt_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal rtt_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal rtt_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe send_packet_buf_queue
  signal send_packet_buf_queue_pipe_write_data: std_logic_vector(31 downto 0);
  signal send_packet_buf_queue_pipe_write_req: std_logic_vector(0 downto 0);
  signal send_packet_buf_queue_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe send_packet_buf_queue
  signal send_packet_buf_queue_pipe_read_data: std_logic_vector(31 downto 0);
  signal send_packet_buf_queue_pipe_read_req: std_logic_vector(0 downto 0);
  signal send_packet_buf_queue_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe send_packet_pipe
  signal send_packet_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal send_packet_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal send_packet_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe send_packet_pipe
  signal send_packet_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal send_packet_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal send_packet_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe src_in0
  signal src_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal src_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal src_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe src_in0
  signal src_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal src_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal src_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe swapped_in_data
  signal swapped_in_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal swapped_in_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal swapped_in_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe swapped_in_data
  signal swapped_in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal swapped_in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal swapped_in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to0_in0
  signal to0_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to0_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to0_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to0_in0
  signal to0_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to0_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to0_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to1_in0
  signal to1_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to1_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to1_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to1_in0
  signal to1_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to1_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to1_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to2_in0
  signal to2_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to2_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to2_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to2_in0
  signal to2_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to2_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to2_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to3_in0
  signal to3_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to3_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to3_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to3_in0
  signal to3_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to3_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to3_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga0_out0
  signal tofpga0_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga0_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga0_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga0_out0
  signal tofpga0_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga0_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga0_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga1_out0
  signal tofpga1_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga1_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga1_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga1_out0
  signal tofpga1_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga1_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga1_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga2_out0
  signal tofpga2_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga2_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga2_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga2_out0
  signal tofpga2_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga2_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga2_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga3_out0
  signal tofpga3_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga3_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga3_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga3_out0
  signal tofpga3_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga3_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga3_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga_port_number
  signal tofpga_port_number_pipe_write_data: std_logic_vector(127 downto 0);
  signal tofpga_port_number_pipe_write_req: std_logic_vector(3 downto 0);
  signal tofpga_port_number_pipe_write_ack: std_logic_vector(3 downto 0);
  -- aggregate signals for read from pipe tofpga_port_number
  signal tofpga_port_number_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga_port_number_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga_port_number_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module GV_15_initializer_in_click_bc
  -- call arbiter for module GV_15_initializer_in_click_bc
  GV_15_initializer_in_click_bc_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => GV_15_initializer_in_click_bc_call_reqs,
      call_acks => GV_15_initializer_in_click_bc_call_acks,
      return_reqs => GV_15_initializer_in_click_bc_return_reqs,
      return_acks => GV_15_initializer_in_click_bc_return_acks,
      call_tag  => GV_15_initializer_in_click_bc_call_tag,
      return_tag  => GV_15_initializer_in_click_bc_return_tag,
      call_mtag => GV_15_initializer_in_click_bc_tag_in,
      return_mtag => GV_15_initializer_in_click_bc_tag_out,
      call_mreq => GV_15_initializer_in_click_bc_start_req,
      call_mack => GV_15_initializer_in_click_bc_start_ack,
      return_mreq => GV_15_initializer_in_click_bc_fin_req,
      return_mack => GV_15_initializer_in_click_bc_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  GV_15_initializer_in_click_bc_instance:GV_15_initializer_in_click_bc-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => GV_15_initializer_in_click_bc_start_req,
      start_ack => GV_15_initializer_in_click_bc_start_ack,
      fin_req => GV_15_initializer_in_click_bc_fin_req,
      fin_ack => GV_15_initializer_in_click_bc_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(8 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(7 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(7 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(4 downto 0),
      tag_in => GV_15_initializer_in_click_bc_tag_in,
      tag_out => GV_15_initializer_in_click_bc_tag_out-- 
    ); -- 
  -- module GV_16_initializer_in_click_bc
  -- call arbiter for module GV_16_initializer_in_click_bc
  GV_16_initializer_in_click_bc_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => GV_16_initializer_in_click_bc_call_reqs,
      call_acks => GV_16_initializer_in_click_bc_call_acks,
      return_reqs => GV_16_initializer_in_click_bc_return_reqs,
      return_acks => GV_16_initializer_in_click_bc_return_acks,
      call_tag  => GV_16_initializer_in_click_bc_call_tag,
      return_tag  => GV_16_initializer_in_click_bc_return_tag,
      call_mtag => GV_16_initializer_in_click_bc_tag_in,
      return_mtag => GV_16_initializer_in_click_bc_tag_out,
      call_mreq => GV_16_initializer_in_click_bc_start_req,
      call_mack => GV_16_initializer_in_click_bc_start_ack,
      return_mreq => GV_16_initializer_in_click_bc_fin_req,
      return_mack => GV_16_initializer_in_click_bc_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  GV_16_initializer_in_click_bc_instance:GV_16_initializer_in_click_bc-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => GV_16_initializer_in_click_bc_start_req,
      start_ack => GV_16_initializer_in_click_bc_start_ack,
      fin_req => GV_16_initializer_in_click_bc_fin_req,
      fin_ack => GV_16_initializer_in_click_bc_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(4 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(6 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 0),
      tag_in => GV_16_initializer_in_click_bc_tag_in,
      tag_out => GV_16_initializer_in_click_bc_tag_out-- 
    ); -- 
  -- module ahir_glue_bswap_i16
  ahir_glue_bswap_i16_i <= ahir_glue_bswap_i16_in_args(15 downto 0);
  ahir_glue_bswap_i16_out_args <= ahir_glue_bswap_i16_ret_val_x_x ;
  -- call arbiter for module ahir_glue_bswap_i16
  ahir_glue_bswap_i16_arbiter: SplitCallArbiter -- 
    generic map( --
      num_reqs => 6,
      call_data_width => 16,
      return_data_width => 16,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => ahir_glue_bswap_i16_call_reqs,
      call_acks => ahir_glue_bswap_i16_call_acks,
      return_reqs => ahir_glue_bswap_i16_return_reqs,
      return_acks => ahir_glue_bswap_i16_return_acks,
      call_data  => ahir_glue_bswap_i16_call_data,
      call_tag  => ahir_glue_bswap_i16_call_tag,
      return_tag  => ahir_glue_bswap_i16_return_tag,
      call_mtag => ahir_glue_bswap_i16_tag_in,
      return_mtag => ahir_glue_bswap_i16_tag_out,
      return_data =>ahir_glue_bswap_i16_return_data,
      call_mreq => ahir_glue_bswap_i16_start_req,
      call_mack => ahir_glue_bswap_i16_start_ack,
      return_mreq => ahir_glue_bswap_i16_fin_req,
      return_mack => ahir_glue_bswap_i16_fin_ack,
      call_mdata => ahir_glue_bswap_i16_in_args,
      return_mdata => ahir_glue_bswap_i16_out_args,
      clk => clk, 
      reset => reset --
    ); --
  ahir_glue_bswap_i16_instance:ahir_glue_bswap_i16-- 
    generic map(tag_length => 3)
    port map(-- 
      i => ahir_glue_bswap_i16_i,
      ret_val_x_x => ahir_glue_bswap_i16_ret_val_x_x,
      start_req => ahir_glue_bswap_i16_start_req,
      start_ack => ahir_glue_bswap_i16_start_ack,
      fin_req => ahir_glue_bswap_i16_fin_req,
      fin_ack => ahir_glue_bswap_i16_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => ahir_glue_bswap_i16_tag_in,
      tag_out => ahir_glue_bswap_i16_tag_out-- 
    ); -- 
  -- module ahir_glue_chk
  ahir_glue_chk_instance:ahir_glue_chk-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_chk_start_req,
      start_ack => ahir_glue_chk_start_ack,
      fin_req => ahir_glue_chk_fin_req,
      fin_ack => ahir_glue_chk_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(8 downto 8),
      memory_space_5_lr_ack => memory_space_5_lr_ack(8 downto 8),
      memory_space_5_lr_addr => memory_space_5_lr_addr(143 downto 128),
      memory_space_5_lr_tag => memory_space_5_lr_tag(98 downto 88),
      memory_space_5_lc_req => memory_space_5_lc_req(8 downto 8),
      memory_space_5_lc_ack => memory_space_5_lc_ack(8 downto 8),
      memory_space_5_lc_data => memory_space_5_lc_data(71 downto 64),
      memory_space_5_lc_tag => memory_space_5_lc_tag(44 downto 40),
      memory_space_5_sr_req => memory_space_5_sr_req(6 downto 6),
      memory_space_5_sr_ack => memory_space_5_sr_ack(6 downto 6),
      memory_space_5_sr_addr => memory_space_5_sr_addr(111 downto 96),
      memory_space_5_sr_data => memory_space_5_sr_data(55 downto 48),
      memory_space_5_sr_tag => memory_space_5_sr_tag(76 downto 66),
      memory_space_5_sc_req => memory_space_5_sc_req(6 downto 6),
      memory_space_5_sc_ack => memory_space_5_sc_ack(6 downto 6),
      memory_space_5_sc_tag => memory_space_5_sc_tag(34 downto 30),
      chk_in0_pipe_read_req => chk_in0_pipe_read_req(0 downto 0),
      chk_in0_pipe_read_ack => chk_in0_pipe_read_ack(0 downto 0),
      chk_in0_pipe_read_data => chk_in0_pipe_read_data(31 downto 0),
      rtt_in0_pipe_write_req => rtt_in0_pipe_write_req(0 downto 0),
      rtt_in0_pipe_write_ack => rtt_in0_pipe_write_ack(0 downto 0),
      rtt_in0_pipe_write_data => rtt_in0_pipe_write_data(31 downto 0),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(5 downto 5),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(5 downto 5),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(95 downto 80),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(11 downto 10),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(5 downto 5),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(5 downto 5),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(95 downto 80),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(11 downto 10),
      ahir_packet_free_call_reqs => ahir_packet_free_call_reqs(2 downto 2),
      ahir_packet_free_call_acks => ahir_packet_free_call_acks(2 downto 2),
      ahir_packet_free_call_data => ahir_packet_free_call_data(95 downto 64),
      ahir_packet_free_call_tag => ahir_packet_free_call_tag(8 downto 6),
      ahir_packet_free_return_reqs => ahir_packet_free_return_reqs(2 downto 2),
      ahir_packet_free_return_acks => ahir_packet_free_return_acks(2 downto 2),
      ahir_packet_free_return_tag => ahir_packet_free_return_tag(8 downto 6),
      tag_in => ahir_glue_chk_tag_in,
      tag_out => ahir_glue_chk_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_chk_tag_in <= (others => '0');
  ahir_glue_chk_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_chk_start_req, start_ack => ahir_glue_chk_start_ack,  fin_req => ahir_glue_chk_fin_req,  fin_ack => ahir_glue_chk_fin_ack);
  -- module ahir_glue_rtt
  ahir_glue_rtt_instance:ahir_glue_rtt-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_rtt_start_req,
      start_ack => ahir_glue_rtt_start_ack,
      fin_req => ahir_glue_rtt_fin_req,
      fin_ack => ahir_glue_rtt_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(8 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(7 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(7 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(4 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(4 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(6 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(7 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(7 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(4 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(3 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(7 downto 7),
      memory_space_5_lr_ack => memory_space_5_lr_ack(7 downto 7),
      memory_space_5_lr_addr => memory_space_5_lr_addr(127 downto 112),
      memory_space_5_lr_tag => memory_space_5_lr_tag(87 downto 77),
      memory_space_5_lc_req => memory_space_5_lc_req(7 downto 7),
      memory_space_5_lc_ack => memory_space_5_lc_ack(7 downto 7),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 56),
      memory_space_5_lc_tag => memory_space_5_lc_tag(39 downto 35),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(7 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(7 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(31 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(3 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      rtt_in0_pipe_read_req => rtt_in0_pipe_read_req(0 downto 0),
      rtt_in0_pipe_read_ack => rtt_in0_pipe_read_ack(0 downto 0),
      rtt_in0_pipe_read_data => rtt_in0_pipe_read_data(31 downto 0),
      to0_in0_pipe_write_req => to0_in0_pipe_write_req(0 downto 0),
      to0_in0_pipe_write_ack => to0_in0_pipe_write_ack(0 downto 0),
      to0_in0_pipe_write_data => to0_in0_pipe_write_data(31 downto 0),
      to1_in0_pipe_write_req => to1_in0_pipe_write_req(0 downto 0),
      to1_in0_pipe_write_ack => to1_in0_pipe_write_ack(0 downto 0),
      to1_in0_pipe_write_data => to1_in0_pipe_write_data(31 downto 0),
      to2_in0_pipe_write_req => to2_in0_pipe_write_req(0 downto 0),
      to2_in0_pipe_write_ack => to2_in0_pipe_write_ack(0 downto 0),
      to2_in0_pipe_write_data => to2_in0_pipe_write_data(31 downto 0),
      to3_in0_pipe_write_req => to3_in0_pipe_write_req(0 downto 0),
      to3_in0_pipe_write_ack => to3_in0_pipe_write_ack(0 downto 0),
      to3_in0_pipe_write_data => to3_in0_pipe_write_data(31 downto 0),
      ahir_packet_free_call_reqs => ahir_packet_free_call_reqs(1 downto 1),
      ahir_packet_free_call_acks => ahir_packet_free_call_acks(1 downto 1),
      ahir_packet_free_call_data => ahir_packet_free_call_data(63 downto 32),
      ahir_packet_free_call_tag => ahir_packet_free_call_tag(5 downto 3),
      ahir_packet_free_return_reqs => ahir_packet_free_return_reqs(1 downto 1),
      ahir_packet_free_return_acks => ahir_packet_free_return_acks(1 downto 1),
      ahir_packet_free_return_tag => ahir_packet_free_return_tag(5 downto 3),
      tag_in => ahir_glue_rtt_tag_in,
      tag_out => ahir_glue_rtt_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_rtt_tag_in <= (others => '0');
  ahir_glue_rtt_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_rtt_start_req, start_ack => ahir_glue_rtt_start_ack,  fin_req => ahir_glue_rtt_fin_req,  fin_ack => ahir_glue_rtt_fin_ack);
  -- module ahir_glue_src
  ahir_glue_src_instance:ahir_glue_src-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_src_start_req,
      start_ack => ahir_glue_src_start_ack,
      fin_req => ahir_glue_src_fin_req,
      fin_ack => ahir_glue_src_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(6 downto 6),
      memory_space_5_lr_ack => memory_space_5_lr_ack(6 downto 6),
      memory_space_5_lr_addr => memory_space_5_lr_addr(111 downto 96),
      memory_space_5_lr_tag => memory_space_5_lr_tag(76 downto 66),
      memory_space_5_lc_req => memory_space_5_lc_req(6 downto 6),
      memory_space_5_lc_ack => memory_space_5_lc_ack(6 downto 6),
      memory_space_5_lc_data => memory_space_5_lc_data(55 downto 48),
      memory_space_5_lc_tag => memory_space_5_lc_tag(34 downto 30),
      memory_space_5_sr_req => memory_space_5_sr_req(5 downto 5),
      memory_space_5_sr_ack => memory_space_5_sr_ack(5 downto 5),
      memory_space_5_sr_addr => memory_space_5_sr_addr(95 downto 80),
      memory_space_5_sr_data => memory_space_5_sr_data(47 downto 40),
      memory_space_5_sr_tag => memory_space_5_sr_tag(65 downto 55),
      memory_space_5_sc_req => memory_space_5_sc_req(5 downto 5),
      memory_space_5_sc_ack => memory_space_5_sc_ack(5 downto 5),
      memory_space_5_sc_tag => memory_space_5_sc_tag(29 downto 25),
      src_in0_pipe_read_req => src_in0_pipe_read_req(0 downto 0),
      src_in0_pipe_read_ack => src_in0_pipe_read_ack(0 downto 0),
      src_in0_pipe_read_data => src_in0_pipe_read_data(31 downto 0),
      chk_in0_pipe_write_req => chk_in0_pipe_write_req(0 downto 0),
      chk_in0_pipe_write_ack => chk_in0_pipe_write_ack(0 downto 0),
      chk_in0_pipe_write_data => chk_in0_pipe_write_data(31 downto 0),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(4 downto 4),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(4 downto 4),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(79 downto 64),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(9 downto 8),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(4 downto 4),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(4 downto 4),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(79 downto 64),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(9 downto 8),
      tag_in => ahir_glue_src_tag_in,
      tag_out => ahir_glue_src_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_src_tag_in <= (others => '0');
  ahir_glue_src_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_src_start_req, start_ack => ahir_glue_src_start_ack,  fin_req => ahir_glue_src_fin_req,  fin_ack => ahir_glue_src_fin_ack);
  -- module ahir_glue_to0
  ahir_glue_to0_instance:ahir_glue_to0-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to0_start_req,
      start_ack => ahir_glue_to0_start_ack,
      fin_req => ahir_glue_to0_fin_req,
      fin_ack => ahir_glue_to0_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(5 downto 5),
      memory_space_5_lr_ack => memory_space_5_lr_ack(5 downto 5),
      memory_space_5_lr_addr => memory_space_5_lr_addr(95 downto 80),
      memory_space_5_lr_tag => memory_space_5_lr_tag(65 downto 55),
      memory_space_5_lc_req => memory_space_5_lc_req(5 downto 5),
      memory_space_5_lc_ack => memory_space_5_lc_ack(5 downto 5),
      memory_space_5_lc_data => memory_space_5_lc_data(47 downto 40),
      memory_space_5_lc_tag => memory_space_5_lc_tag(29 downto 25),
      memory_space_5_sr_req => memory_space_5_sr_req(4 downto 4),
      memory_space_5_sr_ack => memory_space_5_sr_ack(4 downto 4),
      memory_space_5_sr_addr => memory_space_5_sr_addr(79 downto 64),
      memory_space_5_sr_data => memory_space_5_sr_data(39 downto 32),
      memory_space_5_sr_tag => memory_space_5_sr_tag(54 downto 44),
      memory_space_5_sc_req => memory_space_5_sc_req(4 downto 4),
      memory_space_5_sc_ack => memory_space_5_sc_ack(4 downto 4),
      memory_space_5_sc_tag => memory_space_5_sc_tag(24 downto 20),
      to0_in0_pipe_read_req => to0_in0_pipe_read_req(0 downto 0),
      to0_in0_pipe_read_ack => to0_in0_pipe_read_ack(0 downto 0),
      to0_in0_pipe_read_data => to0_in0_pipe_read_data(31 downto 0),
      tofpga0_out0_pipe_write_req => tofpga0_out0_pipe_write_req(0 downto 0),
      tofpga0_out0_pipe_write_ack => tofpga0_out0_pipe_write_ack(0 downto 0),
      tofpga0_out0_pipe_write_data => tofpga0_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(3 downto 3),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(3 downto 3),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(127 downto 96),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(3 downto 3),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(3 downto 3),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(63 downto 48),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(7 downto 6),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(3 downto 3),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(3 downto 3),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(63 downto 48),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(7 downto 6),
      tag_in => ahir_glue_to0_tag_in,
      tag_out => ahir_glue_to0_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to0_tag_in <= (others => '0');
  ahir_glue_to0_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to0_start_req, start_ack => ahir_glue_to0_start_ack,  fin_req => ahir_glue_to0_fin_req,  fin_ack => ahir_glue_to0_fin_ack);
  -- module ahir_glue_to1
  ahir_glue_to1_instance:ahir_glue_to1-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to1_start_req,
      start_ack => ahir_glue_to1_start_ack,
      fin_req => ahir_glue_to1_fin_req,
      fin_ack => ahir_glue_to1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(4 downto 4),
      memory_space_5_lr_ack => memory_space_5_lr_ack(4 downto 4),
      memory_space_5_lr_addr => memory_space_5_lr_addr(79 downto 64),
      memory_space_5_lr_tag => memory_space_5_lr_tag(54 downto 44),
      memory_space_5_lc_req => memory_space_5_lc_req(4 downto 4),
      memory_space_5_lc_ack => memory_space_5_lc_ack(4 downto 4),
      memory_space_5_lc_data => memory_space_5_lc_data(39 downto 32),
      memory_space_5_lc_tag => memory_space_5_lc_tag(24 downto 20),
      memory_space_5_sr_req => memory_space_5_sr_req(3 downto 3),
      memory_space_5_sr_ack => memory_space_5_sr_ack(3 downto 3),
      memory_space_5_sr_addr => memory_space_5_sr_addr(63 downto 48),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 24),
      memory_space_5_sr_tag => memory_space_5_sr_tag(43 downto 33),
      memory_space_5_sc_req => memory_space_5_sc_req(3 downto 3),
      memory_space_5_sc_ack => memory_space_5_sc_ack(3 downto 3),
      memory_space_5_sc_tag => memory_space_5_sc_tag(19 downto 15),
      to1_in0_pipe_read_req => to1_in0_pipe_read_req(0 downto 0),
      to1_in0_pipe_read_ack => to1_in0_pipe_read_ack(0 downto 0),
      to1_in0_pipe_read_data => to1_in0_pipe_read_data(31 downto 0),
      tofpga1_out0_pipe_write_req => tofpga1_out0_pipe_write_req(0 downto 0),
      tofpga1_out0_pipe_write_ack => tofpga1_out0_pipe_write_ack(0 downto 0),
      tofpga1_out0_pipe_write_data => tofpga1_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(2 downto 2),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(2 downto 2),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(95 downto 64),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(2 downto 2),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(2 downto 2),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(47 downto 32),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(5 downto 4),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(2 downto 2),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(2 downto 2),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(47 downto 32),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(5 downto 4),
      tag_in => ahir_glue_to1_tag_in,
      tag_out => ahir_glue_to1_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to1_tag_in <= (others => '0');
  ahir_glue_to1_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to1_start_req, start_ack => ahir_glue_to1_start_ack,  fin_req => ahir_glue_to1_fin_req,  fin_ack => ahir_glue_to1_fin_ack);
  -- module ahir_glue_to2
  ahir_glue_to2_instance:ahir_glue_to2-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to2_start_req,
      start_ack => ahir_glue_to2_start_ack,
      fin_req => ahir_glue_to2_fin_req,
      fin_ack => ahir_glue_to2_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(3 downto 3),
      memory_space_5_lr_ack => memory_space_5_lr_ack(3 downto 3),
      memory_space_5_lr_addr => memory_space_5_lr_addr(63 downto 48),
      memory_space_5_lr_tag => memory_space_5_lr_tag(43 downto 33),
      memory_space_5_lc_req => memory_space_5_lc_req(3 downto 3),
      memory_space_5_lc_ack => memory_space_5_lc_ack(3 downto 3),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 24),
      memory_space_5_lc_tag => memory_space_5_lc_tag(19 downto 15),
      memory_space_5_sr_req => memory_space_5_sr_req(2 downto 2),
      memory_space_5_sr_ack => memory_space_5_sr_ack(2 downto 2),
      memory_space_5_sr_addr => memory_space_5_sr_addr(47 downto 32),
      memory_space_5_sr_data => memory_space_5_sr_data(23 downto 16),
      memory_space_5_sr_tag => memory_space_5_sr_tag(32 downto 22),
      memory_space_5_sc_req => memory_space_5_sc_req(2 downto 2),
      memory_space_5_sc_ack => memory_space_5_sc_ack(2 downto 2),
      memory_space_5_sc_tag => memory_space_5_sc_tag(14 downto 10),
      to2_in0_pipe_read_req => to2_in0_pipe_read_req(0 downto 0),
      to2_in0_pipe_read_ack => to2_in0_pipe_read_ack(0 downto 0),
      to2_in0_pipe_read_data => to2_in0_pipe_read_data(31 downto 0),
      tofpga2_out0_pipe_write_req => tofpga2_out0_pipe_write_req(0 downto 0),
      tofpga2_out0_pipe_write_ack => tofpga2_out0_pipe_write_ack(0 downto 0),
      tofpga2_out0_pipe_write_data => tofpga2_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(1 downto 1),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(1 downto 1),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(63 downto 32),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(1 downto 1),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(1 downto 1),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(31 downto 16),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(3 downto 2),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(1 downto 1),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(1 downto 1),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(31 downto 16),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(3 downto 2),
      tag_in => ahir_glue_to2_tag_in,
      tag_out => ahir_glue_to2_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to2_tag_in <= (others => '0');
  ahir_glue_to2_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to2_start_req, start_ack => ahir_glue_to2_start_ack,  fin_req => ahir_glue_to2_fin_req,  fin_ack => ahir_glue_to2_fin_ack);
  -- module ahir_glue_to3
  ahir_glue_to3_instance:ahir_glue_to3-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to3_start_req,
      start_ack => ahir_glue_to3_start_ack,
      fin_req => ahir_glue_to3_fin_req,
      fin_ack => ahir_glue_to3_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(2 downto 2),
      memory_space_5_lr_ack => memory_space_5_lr_ack(2 downto 2),
      memory_space_5_lr_addr => memory_space_5_lr_addr(47 downto 32),
      memory_space_5_lr_tag => memory_space_5_lr_tag(32 downto 22),
      memory_space_5_lc_req => memory_space_5_lc_req(2 downto 2),
      memory_space_5_lc_ack => memory_space_5_lc_ack(2 downto 2),
      memory_space_5_lc_data => memory_space_5_lc_data(23 downto 16),
      memory_space_5_lc_tag => memory_space_5_lc_tag(14 downto 10),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(31 downto 16),
      memory_space_5_sr_data => memory_space_5_sr_data(15 downto 8),
      memory_space_5_sr_tag => memory_space_5_sr_tag(21 downto 11),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(9 downto 5),
      to3_in0_pipe_read_req => to3_in0_pipe_read_req(0 downto 0),
      to3_in0_pipe_read_ack => to3_in0_pipe_read_ack(0 downto 0),
      to3_in0_pipe_read_data => to3_in0_pipe_read_data(31 downto 0),
      tofpga3_out0_pipe_write_req => tofpga3_out0_pipe_write_req(0 downto 0),
      tofpga3_out0_pipe_write_ack => tofpga3_out0_pipe_write_ack(0 downto 0),
      tofpga3_out0_pipe_write_data => tofpga3_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(0 downto 0),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(0 downto 0),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(31 downto 0),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(0 downto 0),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(0 downto 0),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(15 downto 0),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(1 downto 0),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(0 downto 0),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(0 downto 0),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(15 downto 0),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(1 downto 0),
      tag_in => ahir_glue_to3_tag_in,
      tag_out => ahir_glue_to3_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to3_tag_in <= (others => '0');
  ahir_glue_to3_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to3_start_req, start_ack => ahir_glue_to3_start_ack,  fin_req => ahir_glue_to3_fin_req,  fin_ack => ahir_glue_to3_fin_ack);
  -- module ahir_packet_free
  ahir_packet_free_pkt <= ahir_packet_free_in_args(31 downto 0);
  -- call arbiter for module ahir_packet_free
  ahir_packet_free_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      num_reqs => 3,
      call_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 3--
    )
    port map(-- 
      call_reqs => ahir_packet_free_call_reqs,
      call_acks => ahir_packet_free_call_acks,
      return_reqs => ahir_packet_free_return_reqs,
      return_acks => ahir_packet_free_return_acks,
      call_data  => ahir_packet_free_call_data,
      call_tag  => ahir_packet_free_call_tag,
      return_tag  => ahir_packet_free_return_tag,
      call_mtag => ahir_packet_free_tag_in,
      return_mtag => ahir_packet_free_tag_out,
      call_mreq => ahir_packet_free_start_req,
      call_mack => ahir_packet_free_start_ack,
      return_mreq => ahir_packet_free_fin_req,
      return_mack => ahir_packet_free_fin_ack,
      call_mdata => ahir_packet_free_in_args,
      clk => clk, 
      reset => reset --
    ); --
  ahir_packet_free_instance:ahir_packet_free-- 
    generic map(tag_length => 2)
    port map(-- 
      pkt => ahir_packet_free_pkt,
      start_req => ahir_packet_free_start_req,
      start_ack => ahir_packet_free_start_ack,
      fin_req => ahir_packet_free_fin_req,
      fin_ack => ahir_packet_free_fin_ack,
      clk => clk,
      reset => reset,
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(1 downto 1),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(1 downto 1),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(63 downto 32),
      tag_in => ahir_packet_free_tag_in,
      tag_out => ahir_packet_free_tag_out-- 
    ); -- 
  -- module ahir_packet_get
  ahir_packet_get_out_args <= ahir_packet_get_buf ;
  -- call arbiter for module ahir_packet_get
  ahir_packet_get_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      num_reqs => 1,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => ahir_packet_get_call_reqs,
      call_acks => ahir_packet_get_call_acks,
      return_reqs => ahir_packet_get_return_reqs,
      return_acks => ahir_packet_get_return_acks,
      call_tag  => ahir_packet_get_call_tag,
      return_tag  => ahir_packet_get_return_tag,
      call_mtag => ahir_packet_get_tag_in,
      return_mtag => ahir_packet_get_tag_out,
      return_data =>ahir_packet_get_return_data,
      call_mreq => ahir_packet_get_start_req,
      call_mack => ahir_packet_get_start_ack,
      return_mreq => ahir_packet_get_fin_req,
      return_mack => ahir_packet_get_fin_ack,
      return_mdata => ahir_packet_get_out_args,
      clk => clk, 
      reset => reset --
    ); --
  ahir_packet_get_instance:ahir_packet_get-- 
    generic map(tag_length => 1)
    port map(-- 
      buf => ahir_packet_get_buf,
      start_req => ahir_packet_get_start_req,
      start_ack => ahir_packet_get_start_ack,
      fin_req => ahir_packet_get_fin_req,
      fin_ack => ahir_packet_get_fin_ack,
      clk => clk,
      reset => reset,
      free_queue_pipe_pipe_read_req => free_queue_pipe_pipe_read_req(0 downto 0),
      free_queue_pipe_pipe_read_ack => free_queue_pipe_pipe_read_ack(0 downto 0),
      free_queue_pipe_pipe_read_data => free_queue_pipe_pipe_read_data(31 downto 0),
      tag_in => ahir_packet_get_tag_in,
      tag_out => ahir_packet_get_tag_out-- 
    ); -- 
  -- module analyze_packet
  analyze_packet_pkt <= analyze_packet_in_args(31 downto 0);
  analyze_packet_out_args <= analyze_packet_buf & analyze_packet_wlen & analyze_packet_blen ;
  -- call arbiter for module analyze_packet
  analyze_packet_arbiter: SplitCallArbiter -- 
    generic map( --
      num_reqs => 1,
      call_data_width => 32,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => analyze_packet_call_reqs,
      call_acks => analyze_packet_call_acks,
      return_reqs => analyze_packet_return_reqs,
      return_acks => analyze_packet_return_acks,
      call_data  => analyze_packet_call_data,
      call_tag  => analyze_packet_call_tag,
      return_tag  => analyze_packet_return_tag,
      call_mtag => analyze_packet_tag_in,
      return_mtag => analyze_packet_tag_out,
      return_data =>analyze_packet_return_data,
      call_mreq => analyze_packet_start_req,
      call_mack => analyze_packet_start_ack,
      return_mreq => analyze_packet_fin_req,
      return_mack => analyze_packet_fin_ack,
      call_mdata => analyze_packet_in_args,
      return_mdata => analyze_packet_out_args,
      clk => clk, 
      reset => reset --
    ); --
  analyze_packet_instance:analyze_packet-- 
    generic map(tag_length => 1)
    port map(-- 
      pkt => analyze_packet_pkt,
      buf => analyze_packet_buf,
      wlen => analyze_packet_wlen,
      blen => analyze_packet_blen,
      start_req => analyze_packet_start_req,
      start_ack => analyze_packet_start_ack,
      fin_req => analyze_packet_fin_req,
      fin_ack => analyze_packet_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(31 downto 16),
      memory_space_5_lr_tag => memory_space_5_lr_tag(21 downto 11),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(15 downto 8),
      memory_space_5_lc_tag => memory_space_5_lc_tag(9 downto 5),
      tag_in => analyze_packet_tag_in,
      tag_out => analyze_packet_tag_out-- 
    ); -- 
  -- module click_bc_storage_initializer_x
  -- call arbiter for module click_bc_storage_initializer_x
  click_bc_storage_initializer_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => click_bc_storage_initializer_x_call_reqs,
      call_acks => click_bc_storage_initializer_x_call_acks,
      return_reqs => click_bc_storage_initializer_x_return_reqs,
      return_acks => click_bc_storage_initializer_x_return_acks,
      call_tag  => click_bc_storage_initializer_x_call_tag,
      return_tag  => click_bc_storage_initializer_x_return_tag,
      call_mtag => click_bc_storage_initializer_x_tag_in,
      return_mtag => click_bc_storage_initializer_x_tag_out,
      call_mreq => click_bc_storage_initializer_x_start_req,
      call_mack => click_bc_storage_initializer_x_start_ack,
      return_mreq => click_bc_storage_initializer_x_fin_req,
      return_mack => click_bc_storage_initializer_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  click_bc_storage_initializer_x_instance:click_bc_storage_initializer_x-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => click_bc_storage_initializer_x_start_req,
      start_ack => click_bc_storage_initializer_x_start_ack,
      fin_req => click_bc_storage_initializer_x_fin_req,
      fin_ack => click_bc_storage_initializer_x_fin_ack,
      clk => clk,
      reset => reset,
      GV_15_initializer_in_click_bc_call_reqs => GV_15_initializer_in_click_bc_call_reqs(0 downto 0),
      GV_15_initializer_in_click_bc_call_acks => GV_15_initializer_in_click_bc_call_acks(0 downto 0),
      GV_15_initializer_in_click_bc_call_tag => GV_15_initializer_in_click_bc_call_tag(0 downto 0),
      GV_15_initializer_in_click_bc_return_reqs => GV_15_initializer_in_click_bc_return_reqs(0 downto 0),
      GV_15_initializer_in_click_bc_return_acks => GV_15_initializer_in_click_bc_return_acks(0 downto 0),
      GV_15_initializer_in_click_bc_return_tag => GV_15_initializer_in_click_bc_return_tag(0 downto 0),
      GV_16_initializer_in_click_bc_call_reqs => GV_16_initializer_in_click_bc_call_reqs(0 downto 0),
      GV_16_initializer_in_click_bc_call_acks => GV_16_initializer_in_click_bc_call_acks(0 downto 0),
      GV_16_initializer_in_click_bc_call_tag => GV_16_initializer_in_click_bc_call_tag(0 downto 0),
      GV_16_initializer_in_click_bc_return_reqs => GV_16_initializer_in_click_bc_return_reqs(0 downto 0),
      GV_16_initializer_in_click_bc_return_acks => GV_16_initializer_in_click_bc_return_acks(0 downto 0),
      GV_16_initializer_in_click_bc_return_tag => GV_16_initializer_in_click_bc_return_tag(0 downto 0),
      tag_in => click_bc_storage_initializer_x_tag_in,
      tag_out => click_bc_storage_initializer_x_tag_out-- 
    ); -- 
  -- module free_queue_init
  -- call arbiter for module free_queue_init
  free_queue_init_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => free_queue_init_call_reqs,
      call_acks => free_queue_init_call_acks,
      return_reqs => free_queue_init_return_reqs,
      return_acks => free_queue_init_return_acks,
      call_tag  => free_queue_init_call_tag,
      return_tag  => free_queue_init_return_tag,
      call_mtag => free_queue_init_tag_in,
      return_mtag => free_queue_init_tag_out,
      call_mreq => free_queue_init_start_req,
      call_mack => free_queue_init_start_ack,
      return_mreq => free_queue_init_fin_req,
      return_mack => free_queue_init_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  free_queue_init_instance:free_queue_init-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => free_queue_init_start_req,
      start_ack => free_queue_init_start_ack,
      fin_req => free_queue_init_fin_req,
      fin_ack => free_queue_init_fin_ack,
      clk => clk,
      reset => reset,
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(0 downto 0),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(0 downto 0),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(31 downto 0),
      tag_in => free_queue_init_tag_in,
      tag_out => free_queue_init_tag_out-- 
    ); -- 
  -- module global_storage_initializer_x
  -- call arbiter for module global_storage_initializer_x
  global_storage_initializer_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => global_storage_initializer_x_call_reqs,
      call_acks => global_storage_initializer_x_call_acks,
      return_reqs => global_storage_initializer_x_return_reqs,
      return_acks => global_storage_initializer_x_return_acks,
      call_tag  => global_storage_initializer_x_call_tag,
      return_tag  => global_storage_initializer_x_return_tag,
      call_mtag => global_storage_initializer_x_tag_in,
      return_mtag => global_storage_initializer_x_tag_out,
      call_mreq => global_storage_initializer_x_start_req,
      call_mack => global_storage_initializer_x_start_ack,
      return_mreq => global_storage_initializer_x_fin_req,
      return_mack => global_storage_initializer_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  global_storage_initializer_x_instance:global_storage_initializer_x-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => global_storage_initializer_x_start_req,
      start_ack => global_storage_initializer_x_start_ack,
      fin_req => global_storage_initializer_x_fin_req,
      fin_ack => global_storage_initializer_x_fin_ack,
      clk => clk,
      reset => reset,
      click_bc_storage_initializer_x_call_reqs => click_bc_storage_initializer_x_call_reqs(0 downto 0),
      click_bc_storage_initializer_x_call_acks => click_bc_storage_initializer_x_call_acks(0 downto 0),
      click_bc_storage_initializer_x_call_tag => click_bc_storage_initializer_x_call_tag(0 downto 0),
      click_bc_storage_initializer_x_return_reqs => click_bc_storage_initializer_x_return_reqs(0 downto 0),
      click_bc_storage_initializer_x_return_acks => click_bc_storage_initializer_x_return_acks(0 downto 0),
      click_bc_storage_initializer_x_return_tag => click_bc_storage_initializer_x_return_tag(0 downto 0),
      tag_in => global_storage_initializer_x_tag_in,
      tag_out => global_storage_initializer_x_tag_out-- 
    ); -- 
  -- module receive_packet_pipeline
  receive_packet_pipeline_instance:receive_packet_pipeline-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => receive_packet_pipeline_start_req,
      start_ack => receive_packet_pipeline_start_ack,
      fin_req => receive_packet_pipeline_fin_req,
      fin_ack => receive_packet_pipeline_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(15 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(7 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(10 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(4 downto 0),
      in_ctrl_pipe_read_req => in_ctrl_pipe_read_req(0 downto 0),
      in_ctrl_pipe_read_ack => in_ctrl_pipe_read_ack(0 downto 0),
      in_ctrl_pipe_read_data => in_ctrl_pipe_read_data(7 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      receive_packet_buf_queue_pipe_read_req => receive_packet_buf_queue_pipe_read_req(0 downto 0),
      receive_packet_buf_queue_pipe_read_ack => receive_packet_buf_queue_pipe_read_ack(0 downto 0),
      receive_packet_buf_queue_pipe_read_data => receive_packet_buf_queue_pipe_read_data(31 downto 0),
      swapped_in_data_pipe_read_req => swapped_in_data_pipe_read_req(0 downto 0),
      swapped_in_data_pipe_read_ack => swapped_in_data_pipe_read_ack(0 downto 0),
      swapped_in_data_pipe_read_data => swapped_in_data_pipe_read_data(63 downto 0),
      receive_packet_buf_queue_pipe_write_req => receive_packet_buf_queue_pipe_write_req(0 downto 0),
      receive_packet_buf_queue_pipe_write_ack => receive_packet_buf_queue_pipe_write_ack(0 downto 0),
      receive_packet_buf_queue_pipe_write_data => receive_packet_buf_queue_pipe_write_data(31 downto 0),
      swapped_in_data_pipe_write_req => swapped_in_data_pipe_write_req(0 downto 0),
      swapped_in_data_pipe_write_ack => swapped_in_data_pipe_write_ack(0 downto 0),
      swapped_in_data_pipe_write_data => swapped_in_data_pipe_write_data(63 downto 0),
      receive_packet_pipe_pipe_write_req => receive_packet_pipe_pipe_write_req(0 downto 0),
      receive_packet_pipe_pipe_write_ack => receive_packet_pipe_pipe_write_ack(0 downto 0),
      receive_packet_pipe_pipe_write_data => receive_packet_pipe_pipe_write_data(31 downto 0),
      ahir_packet_get_call_reqs => ahir_packet_get_call_reqs(0 downto 0),
      ahir_packet_get_call_acks => ahir_packet_get_call_acks(0 downto 0),
      ahir_packet_get_call_tag => ahir_packet_get_call_tag(0 downto 0),
      ahir_packet_get_return_reqs => ahir_packet_get_return_reqs(0 downto 0),
      ahir_packet_get_return_acks => ahir_packet_get_return_acks(0 downto 0),
      ahir_packet_get_return_data => ahir_packet_get_return_data(31 downto 0),
      ahir_packet_get_return_tag => ahir_packet_get_return_tag(0 downto 0),
      tag_in => receive_packet_pipeline_tag_in,
      tag_out => receive_packet_pipeline_tag_out-- 
    ); -- 
  -- module will be run forever 
  receive_packet_pipeline_tag_in <= (others => '0');
  receive_packet_pipeline_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => receive_packet_pipeline_start_req, start_ack => receive_packet_pipeline_start_ack,  fin_req => receive_packet_pipeline_fin_req,  fin_ack => receive_packet_pipeline_fin_ack);
  -- module send_packet_pipeline
  send_packet_pipeline_instance:send_packet_pipeline-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => send_packet_pipeline_start_req,
      start_ack => send_packet_pipeline_start_ack,
      fin_req => send_packet_pipeline_fin_req,
      fin_ack => send_packet_pipeline_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(15 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(10 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(7 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(4 downto 0),
      send_packet_buf_queue_pipe_read_req => send_packet_buf_queue_pipe_read_req(0 downto 0),
      send_packet_buf_queue_pipe_read_ack => send_packet_buf_queue_pipe_read_ack(0 downto 0),
      send_packet_buf_queue_pipe_read_data => send_packet_buf_queue_pipe_read_data(31 downto 0),
      send_packet_pipe_pipe_read_req => send_packet_pipe_pipe_read_req(0 downto 0),
      send_packet_pipe_pipe_read_ack => send_packet_pipe_pipe_read_ack(0 downto 0),
      send_packet_pipe_pipe_read_data => send_packet_pipe_pipe_read_data(31 downto 0),
      out_ctrl_pipe_write_req => out_ctrl_pipe_write_req(0 downto 0),
      out_ctrl_pipe_write_ack => out_ctrl_pipe_write_ack(0 downto 0),
      out_ctrl_pipe_write_data => out_ctrl_pipe_write_data(7 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      send_packet_buf_queue_pipe_write_req => send_packet_buf_queue_pipe_write_req(0 downto 0),
      send_packet_buf_queue_pipe_write_ack => send_packet_buf_queue_pipe_write_ack(0 downto 0),
      send_packet_buf_queue_pipe_write_data => send_packet_buf_queue_pipe_write_data(31 downto 0),
      ahir_packet_free_call_reqs => ahir_packet_free_call_reqs(0 downto 0),
      ahir_packet_free_call_acks => ahir_packet_free_call_acks(0 downto 0),
      ahir_packet_free_call_data => ahir_packet_free_call_data(31 downto 0),
      ahir_packet_free_call_tag => ahir_packet_free_call_tag(2 downto 0),
      ahir_packet_free_return_reqs => ahir_packet_free_return_reqs(0 downto 0),
      ahir_packet_free_return_acks => ahir_packet_free_return_acks(0 downto 0),
      ahir_packet_free_return_tag => ahir_packet_free_return_tag(2 downto 0),
      analyze_packet_call_reqs => analyze_packet_call_reqs(0 downto 0),
      analyze_packet_call_acks => analyze_packet_call_acks(0 downto 0),
      analyze_packet_call_data => analyze_packet_call_data(31 downto 0),
      analyze_packet_call_tag => analyze_packet_call_tag(0 downto 0),
      analyze_packet_return_reqs => analyze_packet_return_reqs(0 downto 0),
      analyze_packet_return_acks => analyze_packet_return_acks(0 downto 0),
      analyze_packet_return_data => analyze_packet_return_data(63 downto 0),
      analyze_packet_return_tag => analyze_packet_return_tag(0 downto 0),
      tag_in => send_packet_pipeline_tag_in,
      tag_out => send_packet_pipeline_tag_out-- 
    ); -- 
  -- module will be run forever 
  send_packet_pipeline_tag_in <= (others => '0');
  send_packet_pipeline_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => send_packet_pipeline_start_req, start_ack => send_packet_pipeline_start_ack,  fin_req => send_packet_pipeline_fin_req,  fin_ack => send_packet_pipeline_fin_ack);
  -- module wrapper_input
  wrapper_input_instance:wrapper_input-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_input_start_req,
      start_ack => wrapper_input_start_ack,
      fin_req => wrapper_input_fin_req,
      fin_ack => wrapper_input_fin_ack,
      clk => clk,
      reset => reset,
      receive_packet_pipe_pipe_read_req => receive_packet_pipe_pipe_read_req(0 downto 0),
      receive_packet_pipe_pipe_read_ack => receive_packet_pipe_pipe_read_ack(0 downto 0),
      receive_packet_pipe_pipe_read_data => receive_packet_pipe_pipe_read_data(31 downto 0),
      src_in0_pipe_write_req => src_in0_pipe_write_req(0 downto 0),
      src_in0_pipe_write_ack => src_in0_pipe_write_ack(0 downto 0),
      src_in0_pipe_write_data => src_in0_pipe_write_data(31 downto 0),
      free_queue_init_call_reqs => free_queue_init_call_reqs(0 downto 0),
      free_queue_init_call_acks => free_queue_init_call_acks(0 downto 0),
      free_queue_init_call_tag => free_queue_init_call_tag(0 downto 0),
      free_queue_init_return_reqs => free_queue_init_return_reqs(0 downto 0),
      free_queue_init_return_acks => free_queue_init_return_acks(0 downto 0),
      free_queue_init_return_tag => free_queue_init_return_tag(0 downto 0),
      global_storage_initializer_x_call_reqs => global_storage_initializer_x_call_reqs(0 downto 0),
      global_storage_initializer_x_call_acks => global_storage_initializer_x_call_acks(0 downto 0),
      global_storage_initializer_x_call_tag => global_storage_initializer_x_call_tag(0 downto 0),
      global_storage_initializer_x_return_reqs => global_storage_initializer_x_return_reqs(0 downto 0),
      global_storage_initializer_x_return_acks => global_storage_initializer_x_return_acks(0 downto 0),
      global_storage_initializer_x_return_tag => global_storage_initializer_x_return_tag(0 downto 0),
      tag_in => wrapper_input_tag_in,
      tag_out => wrapper_input_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_input_tag_in <= (others => '0');
  wrapper_input_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_input_start_req, start_ack => wrapper_input_start_ack,  fin_req => wrapper_input_fin_req,  fin_ack => wrapper_input_fin_ack);
  -- module wrapper_output
  wrapper_output_instance:wrapper_output-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_output_start_req,
      start_ack => wrapper_output_start_ack,
      fin_req => wrapper_output_fin_req,
      fin_ack => wrapper_output_fin_ack,
      clk => clk,
      reset => reset,
      tofpga0_out0_pipe_read_req => tofpga0_out0_pipe_read_req(0 downto 0),
      tofpga0_out0_pipe_read_ack => tofpga0_out0_pipe_read_ack(0 downto 0),
      tofpga0_out0_pipe_read_data => tofpga0_out0_pipe_read_data(31 downto 0),
      tofpga1_out0_pipe_read_req => tofpga1_out0_pipe_read_req(0 downto 0),
      tofpga1_out0_pipe_read_ack => tofpga1_out0_pipe_read_ack(0 downto 0),
      tofpga1_out0_pipe_read_data => tofpga1_out0_pipe_read_data(31 downto 0),
      tofpga2_out0_pipe_read_req => tofpga2_out0_pipe_read_req(0 downto 0),
      tofpga2_out0_pipe_read_ack => tofpga2_out0_pipe_read_ack(0 downto 0),
      tofpga2_out0_pipe_read_data => tofpga2_out0_pipe_read_data(31 downto 0),
      tofpga3_out0_pipe_read_req => tofpga3_out0_pipe_read_req(0 downto 0),
      tofpga3_out0_pipe_read_ack => tofpga3_out0_pipe_read_ack(0 downto 0),
      tofpga3_out0_pipe_read_data => tofpga3_out0_pipe_read_data(31 downto 0),
      tofpga_port_number_pipe_read_req => tofpga_port_number_pipe_read_req(0 downto 0),
      tofpga_port_number_pipe_read_ack => tofpga_port_number_pipe_read_ack(0 downto 0),
      tofpga_port_number_pipe_read_data => tofpga_port_number_pipe_read_data(31 downto 0),
      send_packet_pipe_pipe_write_req => send_packet_pipe_pipe_write_req(0 downto 0),
      send_packet_pipe_pipe_write_ack => send_packet_pipe_pipe_write_ack(0 downto 0),
      send_packet_pipe_pipe_write_data => send_packet_pipe_pipe_write_data(31 downto 0),
      tag_in => wrapper_output_tag_in,
      tag_out => wrapper_output_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_output_tag_in <= (others => '0');
  wrapper_output_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_output_start_req, start_ack => wrapper_output_start_ack,  fin_req => wrapper_output_fin_req,  fin_ack => wrapper_output_fin_ack);
  chk_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => chk_in0_pipe_read_req,
      read_ack => chk_in0_pipe_read_ack,
      read_data => chk_in0_pipe_read_data,
      write_req => chk_in0_pipe_write_req,
      write_ack => chk_in0_pipe_write_ack,
      write_data => chk_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 32,
      depth => 16 --
    )
    port map( -- 
      read_req => free_queue_pipe_pipe_read_req,
      read_ack => free_queue_pipe_pipe_read_ack,
      read_data => free_queue_pipe_pipe_read_data,
      write_req => free_queue_pipe_pipe_write_req,
      write_ack => free_queue_pipe_pipe_write_ack,
      write_data => free_queue_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => in_ctrl_pipe_read_req,
      read_ack => in_ctrl_pipe_read_ack,
      read_data => in_ctrl_pipe_read_data,
      write_req => in_ctrl_pipe_write_req,
      write_ack => in_ctrl_pipe_write_ack,
      write_data => in_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => out_ctrl_pipe_read_req,
      read_ack => out_ctrl_pipe_read_ack,
      read_data => out_ctrl_pipe_read_data,
      write_req => out_ctrl_pipe_write_req,
      write_ack => out_ctrl_pipe_write_ack,
      write_data => out_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  receive_packet_buf_queue_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 4 --
    )
    port map( -- 
      read_req => receive_packet_buf_queue_pipe_read_req,
      read_ack => receive_packet_buf_queue_pipe_read_ack,
      read_data => receive_packet_buf_queue_pipe_read_data,
      write_req => receive_packet_buf_queue_pipe_write_req,
      write_ack => receive_packet_buf_queue_pipe_write_ack,
      write_data => receive_packet_buf_queue_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  receive_packet_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => receive_packet_pipe_pipe_read_req,
      read_ack => receive_packet_pipe_pipe_read_ack,
      read_data => receive_packet_pipe_pipe_read_data,
      write_req => receive_packet_pipe_pipe_write_req,
      write_ack => receive_packet_pipe_pipe_write_ack,
      write_data => receive_packet_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  rtt_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => rtt_in0_pipe_read_req,
      read_ack => rtt_in0_pipe_read_ack,
      read_data => rtt_in0_pipe_read_data,
      write_req => rtt_in0_pipe_write_req,
      write_ack => rtt_in0_pipe_write_ack,
      write_data => rtt_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  send_packet_buf_queue_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 4 --
    )
    port map( -- 
      read_req => send_packet_buf_queue_pipe_read_req,
      read_ack => send_packet_buf_queue_pipe_read_ack,
      read_data => send_packet_buf_queue_pipe_read_data,
      write_req => send_packet_buf_queue_pipe_write_req,
      write_ack => send_packet_buf_queue_pipe_write_ack,
      write_data => send_packet_buf_queue_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  send_packet_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => send_packet_pipe_pipe_read_req,
      read_ack => send_packet_pipe_pipe_read_ack,
      read_data => send_packet_pipe_pipe_read_data,
      write_req => send_packet_pipe_pipe_write_req,
      write_ack => send_packet_pipe_pipe_write_ack,
      write_data => send_packet_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  src_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => src_in0_pipe_read_req,
      read_ack => src_in0_pipe_read_ack,
      read_data => src_in0_pipe_read_data,
      write_req => src_in0_pipe_write_req,
      write_ack => src_in0_pipe_write_ack,
      write_data => src_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  swapped_in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => swapped_in_data_pipe_read_req,
      read_ack => swapped_in_data_pipe_read_ack,
      read_data => swapped_in_data_pipe_read_data,
      write_req => swapped_in_data_pipe_write_req,
      write_ack => swapped_in_data_pipe_write_ack,
      write_data => swapped_in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to0_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to0_in0_pipe_read_req,
      read_ack => to0_in0_pipe_read_ack,
      read_data => to0_in0_pipe_read_data,
      write_req => to0_in0_pipe_write_req,
      write_ack => to0_in0_pipe_write_ack,
      write_data => to0_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to1_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to1_in0_pipe_read_req,
      read_ack => to1_in0_pipe_read_ack,
      read_data => to1_in0_pipe_read_data,
      write_req => to1_in0_pipe_write_req,
      write_ack => to1_in0_pipe_write_ack,
      write_data => to1_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to2_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to2_in0_pipe_read_req,
      read_ack => to2_in0_pipe_read_ack,
      read_data => to2_in0_pipe_read_data,
      write_req => to2_in0_pipe_write_req,
      write_ack => to2_in0_pipe_write_ack,
      write_data => to2_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to3_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to3_in0_pipe_read_req,
      read_ack => to3_in0_pipe_read_ack,
      read_data => to3_in0_pipe_read_data,
      write_req => to3_in0_pipe_write_req,
      write_ack => to3_in0_pipe_write_ack,
      write_data => to3_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga0_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga0_out0_pipe_read_req,
      read_ack => tofpga0_out0_pipe_read_ack,
      read_data => tofpga0_out0_pipe_read_data,
      write_req => tofpga0_out0_pipe_write_req,
      write_ack => tofpga0_out0_pipe_write_ack,
      write_data => tofpga0_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga1_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga1_out0_pipe_read_req,
      read_ack => tofpga1_out0_pipe_read_ack,
      read_data => tofpga1_out0_pipe_read_data,
      write_req => tofpga1_out0_pipe_write_req,
      write_ack => tofpga1_out0_pipe_write_ack,
      write_data => tofpga1_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga2_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga2_out0_pipe_read_req,
      read_ack => tofpga2_out0_pipe_read_ack,
      read_data => tofpga2_out0_pipe_read_data,
      write_req => tofpga2_out0_pipe_write_req,
      write_ack => tofpga2_out0_pipe_write_ack,
      write_data => tofpga2_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga3_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga3_out0_pipe_read_req,
      read_ack => tofpga3_out0_pipe_read_ack,
      read_data => tofpga3_out0_pipe_read_data,
      write_req => tofpga3_out0_pipe_write_req,
      write_ack => tofpga3_out0_pipe_write_ack,
      write_data => tofpga3_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga_port_number_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 4,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga_port_number_pipe_read_req,
      read_ack => tofpga_port_number_pipe_read_ack,
      read_data => tofpga_port_number_pipe_read_data,
      write_req => tofpga_port_number_pipe_write_req,
      write_ack => tofpga_port_number_pipe_write_ack,
      write_data => tofpga_port_number_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 9,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 5,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 5,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 9,
      num_stores => 7,
      addr_width => 16,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 6,
      number_of_banks => 4,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system_Test_Bench is -- 
  -- 
end entity;
architecture Default of ahir_system_Test_Bench is -- 
  component ahir_system is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
      in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
      in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
      in_data_pipe_write_data: in std_logic_vector(63 downto 0);
      in_data_pipe_write_req : in std_logic_vector(0 downto 0);
      in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
      out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
      out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
      out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
      out_data_pipe_read_data: out std_logic_vector(63 downto 0);
      out_data_pipe_read_req : in std_logic_vector(0 downto 0);
      out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  signal clk: std_logic := '0';
  signal reset: std_logic := '1';
  signal ahir_glue_chk_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_chk_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_chk_start_req : std_logic := '0';
  signal ahir_glue_chk_start_ack : std_logic := '0';
  signal ahir_glue_chk_fin_req   : std_logic := '0';
  signal ahir_glue_chk_fin_ack   : std_logic := '0';
  signal ahir_glue_rtt_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_rtt_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_rtt_start_req : std_logic := '0';
  signal ahir_glue_rtt_start_ack : std_logic := '0';
  signal ahir_glue_rtt_fin_req   : std_logic := '0';
  signal ahir_glue_rtt_fin_ack   : std_logic := '0';
  signal ahir_glue_src_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_src_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_src_start_req : std_logic := '0';
  signal ahir_glue_src_start_ack : std_logic := '0';
  signal ahir_glue_src_fin_req   : std_logic := '0';
  signal ahir_glue_src_fin_ack   : std_logic := '0';
  signal ahir_glue_to0_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to0_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to0_start_req : std_logic := '0';
  signal ahir_glue_to0_start_ack : std_logic := '0';
  signal ahir_glue_to0_fin_req   : std_logic := '0';
  signal ahir_glue_to0_fin_ack   : std_logic := '0';
  signal ahir_glue_to1_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to1_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to1_start_req : std_logic := '0';
  signal ahir_glue_to1_start_ack : std_logic := '0';
  signal ahir_glue_to1_fin_req   : std_logic := '0';
  signal ahir_glue_to1_fin_ack   : std_logic := '0';
  signal ahir_glue_to2_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to2_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to2_start_req : std_logic := '0';
  signal ahir_glue_to2_start_ack : std_logic := '0';
  signal ahir_glue_to2_fin_req   : std_logic := '0';
  signal ahir_glue_to2_fin_ack   : std_logic := '0';
  signal ahir_glue_to3_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to3_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to3_start_req : std_logic := '0';
  signal ahir_glue_to3_start_ack : std_logic := '0';
  signal ahir_glue_to3_fin_req   : std_logic := '0';
  signal ahir_glue_to3_fin_ack   : std_logic := '0';
  signal receive_packet_pipeline_tag_in: std_logic_vector(0 downto 0);
  signal receive_packet_pipeline_tag_out: std_logic_vector(0 downto 0);
  signal receive_packet_pipeline_start_req : std_logic := '0';
  signal receive_packet_pipeline_start_ack : std_logic := '0';
  signal receive_packet_pipeline_fin_req   : std_logic := '0';
  signal receive_packet_pipeline_fin_ack   : std_logic := '0';
  signal send_packet_pipeline_tag_in: std_logic_vector(0 downto 0);
  signal send_packet_pipeline_tag_out: std_logic_vector(0 downto 0);
  signal send_packet_pipeline_start_req : std_logic := '0';
  signal send_packet_pipeline_start_ack : std_logic := '0';
  signal send_packet_pipeline_fin_req   : std_logic := '0';
  signal send_packet_pipeline_fin_ack   : std_logic := '0';
  signal wrapper_input_tag_in: std_logic_vector(0 downto 0);
  signal wrapper_input_tag_out: std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic := '0';
  signal wrapper_input_start_ack : std_logic := '0';
  signal wrapper_input_fin_req   : std_logic := '0';
  signal wrapper_input_fin_ack   : std_logic := '0';
  signal wrapper_output_tag_in: std_logic_vector(0 downto 0);
  signal wrapper_output_tag_out: std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic := '0';
  signal wrapper_output_start_ack : std_logic := '0';
  signal wrapper_output_fin_req   : std_logic := '0';
  signal wrapper_output_fin_ack   : std_logic := '0';
  -- write to pipe in_ctrl
  signal in_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_write_req : std_logic_vector(0 downto 0) := (others => '0');
  signal in_ctrl_pipe_write_ack : std_logic_vector(0 downto 0);
  -- write to pipe in_data
  signal in_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_write_req : std_logic_vector(0 downto 0) := (others => '0');
  signal in_data_pipe_write_ack : std_logic_vector(0 downto 0);
  -- read from pipe out_ctrl
  signal out_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_read_req : std_logic_vector(0 downto 0) := (others => '0');
  signal out_ctrl_pipe_read_ack : std_logic_vector(0 downto 0);
  -- read from pipe out_data
  signal out_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_read_req : std_logic_vector(0 downto 0) := (others => '0');
  signal out_data_pipe_read_ack : std_logic_vector(0 downto 0);
  -- 
begin --
  -- clock/reset generation 
  clk <= not clk after 5 ns;
  process
  begin --
    wait until clk = '1';
    reset <= '0';
    wait;
    --
  end process;
  -- a rudimentary tb.. will start all the top-level modules ..
  ahir_system_instance: ahir_system -- 
    port map ( -- 
      clk => clk,
      reset => reset,
      in_ctrl_pipe_write_data  => in_ctrl_pipe_write_data, 
      in_ctrl_pipe_write_req  => in_ctrl_pipe_write_req, 
      in_ctrl_pipe_write_ack  => in_ctrl_pipe_write_ack,
      in_data_pipe_write_data  => in_data_pipe_write_data, 
      in_data_pipe_write_req  => in_data_pipe_write_req, 
      in_data_pipe_write_ack  => in_data_pipe_write_ack,
      out_ctrl_pipe_read_data  => out_ctrl_pipe_read_data, 
      out_ctrl_pipe_read_req  => out_ctrl_pipe_read_req, 
      out_ctrl_pipe_read_ack  => out_ctrl_pipe_read_ack ,
      out_data_pipe_read_data  => out_data_pipe_read_data, 
      out_data_pipe_read_req  => out_data_pipe_read_req, 
      out_data_pipe_read_ack  => out_data_pipe_read_ack ); -- 
  -- 
end Default;
