-------------------------------------------------------
--  Copyright (c) 2011 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version : 11.1
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : X_BUFG_LB.vhd
-- \   \  /  \      
--  \__ \/\__ \                   
--                                 
--  Generated by    : /home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
--  Revision: 1.0
--    11/15/11 - 634082 - connected ouput.
--  End Revision
-------------------------------------------------------

----- CELL X_BUFG_LB -----

library IEEE;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

library simprim;
use simprim.VCOMPONENTS.all;
use simprim.VPACKAGE.all;

  entity X_BUFG_LB is
    generic (
      TimingChecksOn : boolean := TRUE;
      InstancePath   : string  := "*";
      Xon            : boolean := TRUE;
      MsgOn          : boolean := FALSE;
      LOC            : string  := "UNPLACED";
      tipd_CLKIN : VitalDelayType01 :=  (0 ps, 0 ps);
      tpd_CLKIN_CLKOUT : VitalDelayType01 := (0 ps, 0 ps);
      ticd_CLKIN : VitalDelayType := 0 ps
    );

    port (
      CLKOUT               : out std_ulogic;
      CLKIN                : in std_ulogic      
    );
    attribute VITAL_LEVEL0 of X_BUFG_LB :     entity is true;
  end X_BUFG_LB;

  architecture X_BUFG_LB_V of X_BUFG_LB is
    TYPE VitalTimingDataArrayType IS ARRAY (NATURAL RANGE <>) OF VitalTimingDataType;
    
    signal CLKOUT_out : std_ulogic;
    signal CLKIN_ipd : std_ulogic;
    signal CLKIN_dly : std_ulogic;
    
    
    begin
    
    WireDelay : block
    begin
      VitalWireDelay (CLKIN_ipd,CLKIN,tipd_CLKIN);
    end block;
    
    SignalDelay : block
    begin
      VitalSignalDelay (CLKIN_dly,CLKIN_ipd,ticd_CLKIN);
    end block;

    CLKOUT_out <= CLKIN_dly;
    
    TIMING : process
      variable CLKOUT_GlitchData : VitalGlitchDataType;

      begin

        VitalPathDelay01
        (
          OutSignal     => CLKOUT,
          GlitchData    => CLKOUT_GlitchData,
          OutSignalName => "CLKOUT",
          OutTemp       => CLKOUT_out,
          Paths       => (0 => (CLKIN_dly'last_event, tpd_CLKIN_CLKOUT,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
      wait on
        CLKOUT_out;
    end process TIMING;
  end X_BUFG_LB_V;
